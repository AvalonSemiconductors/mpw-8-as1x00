// This is the unpowered netlist.
module wrapped_tms1x00 (oram_csb,
    ram_csb,
    ram_web,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_dat_i,
    wbs_stb_i,
    wbs_we_i,
    io_in,
    io_oeb,
    io_out,
    oram_addr,
    oram_value,
    ram_adrb,
    ram_wmask,
    wbs_adr_i);
 output oram_csb;
 output ram_csb;
 output ram_web;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_dat_i;
 input wbs_stb_i;
 input wbs_we_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 output [8:0] oram_addr;
 input [31:0] oram_value;
 output [8:0] ram_adrb;
 output [3:0] ram_wmask;
 input [31:0] wbs_adr_i;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire net126;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net127;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net128;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net129;
 wire net130;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net112;
 wire net113;
 wire net114;
 wire net122;
 wire net123;
 wire net124;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net125;
 wire net131;
 wire net132;
 wire net133;
 wire clknet_leaf_0_wb_clk_i;
 wire \tms1x00.A[0] ;
 wire \tms1x00.A[1] ;
 wire \tms1x00.A[2] ;
 wire \tms1x00.A[3] ;
 wire \tms1x00.CL ;
 wire \tms1x00.K_latch[0] ;
 wire \tms1x00.K_latch[1] ;
 wire \tms1x00.K_latch[2] ;
 wire \tms1x00.K_latch[3] ;
 wire \tms1x00.N[0] ;
 wire \tms1x00.N[1] ;
 wire \tms1x00.N[2] ;
 wire \tms1x00.N[3] ;
 wire \tms1x00.PA[0] ;
 wire \tms1x00.PA[1] ;
 wire \tms1x00.PA[2] ;
 wire \tms1x00.PA[3] ;
 wire \tms1x00.PB[0] ;
 wire \tms1x00.PB[1] ;
 wire \tms1x00.PB[2] ;
 wire \tms1x00.PB[3] ;
 wire \tms1x00.PC[0] ;
 wire \tms1x00.PC[1] ;
 wire \tms1x00.PC[2] ;
 wire \tms1x00.PC[3] ;
 wire \tms1x00.PC[4] ;
 wire \tms1x00.PC[5] ;
 wire \tms1x00.P[0] ;
 wire \tms1x00.P[1] ;
 wire \tms1x00.P[2] ;
 wire \tms1x00.P[3] ;
 wire \tms1x00.RAM[0][0] ;
 wire \tms1x00.RAM[0][1] ;
 wire \tms1x00.RAM[0][2] ;
 wire \tms1x00.RAM[0][3] ;
 wire \tms1x00.RAM[100][0] ;
 wire \tms1x00.RAM[100][1] ;
 wire \tms1x00.RAM[100][2] ;
 wire \tms1x00.RAM[100][3] ;
 wire \tms1x00.RAM[101][0] ;
 wire \tms1x00.RAM[101][1] ;
 wire \tms1x00.RAM[101][2] ;
 wire \tms1x00.RAM[101][3] ;
 wire \tms1x00.RAM[102][0] ;
 wire \tms1x00.RAM[102][1] ;
 wire \tms1x00.RAM[102][2] ;
 wire \tms1x00.RAM[102][3] ;
 wire \tms1x00.RAM[103][0] ;
 wire \tms1x00.RAM[103][1] ;
 wire \tms1x00.RAM[103][2] ;
 wire \tms1x00.RAM[103][3] ;
 wire \tms1x00.RAM[104][0] ;
 wire \tms1x00.RAM[104][1] ;
 wire \tms1x00.RAM[104][2] ;
 wire \tms1x00.RAM[104][3] ;
 wire \tms1x00.RAM[105][0] ;
 wire \tms1x00.RAM[105][1] ;
 wire \tms1x00.RAM[105][2] ;
 wire \tms1x00.RAM[105][3] ;
 wire \tms1x00.RAM[106][0] ;
 wire \tms1x00.RAM[106][1] ;
 wire \tms1x00.RAM[106][2] ;
 wire \tms1x00.RAM[106][3] ;
 wire \tms1x00.RAM[107][0] ;
 wire \tms1x00.RAM[107][1] ;
 wire \tms1x00.RAM[107][2] ;
 wire \tms1x00.RAM[107][3] ;
 wire \tms1x00.RAM[108][0] ;
 wire \tms1x00.RAM[108][1] ;
 wire \tms1x00.RAM[108][2] ;
 wire \tms1x00.RAM[108][3] ;
 wire \tms1x00.RAM[109][0] ;
 wire \tms1x00.RAM[109][1] ;
 wire \tms1x00.RAM[109][2] ;
 wire \tms1x00.RAM[109][3] ;
 wire \tms1x00.RAM[10][0] ;
 wire \tms1x00.RAM[10][1] ;
 wire \tms1x00.RAM[10][2] ;
 wire \tms1x00.RAM[10][3] ;
 wire \tms1x00.RAM[110][0] ;
 wire \tms1x00.RAM[110][1] ;
 wire \tms1x00.RAM[110][2] ;
 wire \tms1x00.RAM[110][3] ;
 wire \tms1x00.RAM[111][0] ;
 wire \tms1x00.RAM[111][1] ;
 wire \tms1x00.RAM[111][2] ;
 wire \tms1x00.RAM[111][3] ;
 wire \tms1x00.RAM[112][0] ;
 wire \tms1x00.RAM[112][1] ;
 wire \tms1x00.RAM[112][2] ;
 wire \tms1x00.RAM[112][3] ;
 wire \tms1x00.RAM[113][0] ;
 wire \tms1x00.RAM[113][1] ;
 wire \tms1x00.RAM[113][2] ;
 wire \tms1x00.RAM[113][3] ;
 wire \tms1x00.RAM[114][0] ;
 wire \tms1x00.RAM[114][1] ;
 wire \tms1x00.RAM[114][2] ;
 wire \tms1x00.RAM[114][3] ;
 wire \tms1x00.RAM[115][0] ;
 wire \tms1x00.RAM[115][1] ;
 wire \tms1x00.RAM[115][2] ;
 wire \tms1x00.RAM[115][3] ;
 wire \tms1x00.RAM[116][0] ;
 wire \tms1x00.RAM[116][1] ;
 wire \tms1x00.RAM[116][2] ;
 wire \tms1x00.RAM[116][3] ;
 wire \tms1x00.RAM[117][0] ;
 wire \tms1x00.RAM[117][1] ;
 wire \tms1x00.RAM[117][2] ;
 wire \tms1x00.RAM[117][3] ;
 wire \tms1x00.RAM[118][0] ;
 wire \tms1x00.RAM[118][1] ;
 wire \tms1x00.RAM[118][2] ;
 wire \tms1x00.RAM[118][3] ;
 wire \tms1x00.RAM[119][0] ;
 wire \tms1x00.RAM[119][1] ;
 wire \tms1x00.RAM[119][2] ;
 wire \tms1x00.RAM[119][3] ;
 wire \tms1x00.RAM[11][0] ;
 wire \tms1x00.RAM[11][1] ;
 wire \tms1x00.RAM[11][2] ;
 wire \tms1x00.RAM[11][3] ;
 wire \tms1x00.RAM[120][0] ;
 wire \tms1x00.RAM[120][1] ;
 wire \tms1x00.RAM[120][2] ;
 wire \tms1x00.RAM[120][3] ;
 wire \tms1x00.RAM[121][0] ;
 wire \tms1x00.RAM[121][1] ;
 wire \tms1x00.RAM[121][2] ;
 wire \tms1x00.RAM[121][3] ;
 wire \tms1x00.RAM[122][0] ;
 wire \tms1x00.RAM[122][1] ;
 wire \tms1x00.RAM[122][2] ;
 wire \tms1x00.RAM[122][3] ;
 wire \tms1x00.RAM[123][0] ;
 wire \tms1x00.RAM[123][1] ;
 wire \tms1x00.RAM[123][2] ;
 wire \tms1x00.RAM[123][3] ;
 wire \tms1x00.RAM[124][0] ;
 wire \tms1x00.RAM[124][1] ;
 wire \tms1x00.RAM[124][2] ;
 wire \tms1x00.RAM[124][3] ;
 wire \tms1x00.RAM[125][0] ;
 wire \tms1x00.RAM[125][1] ;
 wire \tms1x00.RAM[125][2] ;
 wire \tms1x00.RAM[125][3] ;
 wire \tms1x00.RAM[126][0] ;
 wire \tms1x00.RAM[126][1] ;
 wire \tms1x00.RAM[126][2] ;
 wire \tms1x00.RAM[126][3] ;
 wire \tms1x00.RAM[127][0] ;
 wire \tms1x00.RAM[127][1] ;
 wire \tms1x00.RAM[127][2] ;
 wire \tms1x00.RAM[127][3] ;
 wire \tms1x00.RAM[12][0] ;
 wire \tms1x00.RAM[12][1] ;
 wire \tms1x00.RAM[12][2] ;
 wire \tms1x00.RAM[12][3] ;
 wire \tms1x00.RAM[13][0] ;
 wire \tms1x00.RAM[13][1] ;
 wire \tms1x00.RAM[13][2] ;
 wire \tms1x00.RAM[13][3] ;
 wire \tms1x00.RAM[14][0] ;
 wire \tms1x00.RAM[14][1] ;
 wire \tms1x00.RAM[14][2] ;
 wire \tms1x00.RAM[14][3] ;
 wire \tms1x00.RAM[15][0] ;
 wire \tms1x00.RAM[15][1] ;
 wire \tms1x00.RAM[15][2] ;
 wire \tms1x00.RAM[15][3] ;
 wire \tms1x00.RAM[16][0] ;
 wire \tms1x00.RAM[16][1] ;
 wire \tms1x00.RAM[16][2] ;
 wire \tms1x00.RAM[16][3] ;
 wire \tms1x00.RAM[17][0] ;
 wire \tms1x00.RAM[17][1] ;
 wire \tms1x00.RAM[17][2] ;
 wire \tms1x00.RAM[17][3] ;
 wire \tms1x00.RAM[18][0] ;
 wire \tms1x00.RAM[18][1] ;
 wire \tms1x00.RAM[18][2] ;
 wire \tms1x00.RAM[18][3] ;
 wire \tms1x00.RAM[19][0] ;
 wire \tms1x00.RAM[19][1] ;
 wire \tms1x00.RAM[19][2] ;
 wire \tms1x00.RAM[19][3] ;
 wire \tms1x00.RAM[1][0] ;
 wire \tms1x00.RAM[1][1] ;
 wire \tms1x00.RAM[1][2] ;
 wire \tms1x00.RAM[1][3] ;
 wire \tms1x00.RAM[20][0] ;
 wire \tms1x00.RAM[20][1] ;
 wire \tms1x00.RAM[20][2] ;
 wire \tms1x00.RAM[20][3] ;
 wire \tms1x00.RAM[21][0] ;
 wire \tms1x00.RAM[21][1] ;
 wire \tms1x00.RAM[21][2] ;
 wire \tms1x00.RAM[21][3] ;
 wire \tms1x00.RAM[22][0] ;
 wire \tms1x00.RAM[22][1] ;
 wire \tms1x00.RAM[22][2] ;
 wire \tms1x00.RAM[22][3] ;
 wire \tms1x00.RAM[23][0] ;
 wire \tms1x00.RAM[23][1] ;
 wire \tms1x00.RAM[23][2] ;
 wire \tms1x00.RAM[23][3] ;
 wire \tms1x00.RAM[24][0] ;
 wire \tms1x00.RAM[24][1] ;
 wire \tms1x00.RAM[24][2] ;
 wire \tms1x00.RAM[24][3] ;
 wire \tms1x00.RAM[25][0] ;
 wire \tms1x00.RAM[25][1] ;
 wire \tms1x00.RAM[25][2] ;
 wire \tms1x00.RAM[25][3] ;
 wire \tms1x00.RAM[26][0] ;
 wire \tms1x00.RAM[26][1] ;
 wire \tms1x00.RAM[26][2] ;
 wire \tms1x00.RAM[26][3] ;
 wire \tms1x00.RAM[27][0] ;
 wire \tms1x00.RAM[27][1] ;
 wire \tms1x00.RAM[27][2] ;
 wire \tms1x00.RAM[27][3] ;
 wire \tms1x00.RAM[28][0] ;
 wire \tms1x00.RAM[28][1] ;
 wire \tms1x00.RAM[28][2] ;
 wire \tms1x00.RAM[28][3] ;
 wire \tms1x00.RAM[29][0] ;
 wire \tms1x00.RAM[29][1] ;
 wire \tms1x00.RAM[29][2] ;
 wire \tms1x00.RAM[29][3] ;
 wire \tms1x00.RAM[2][0] ;
 wire \tms1x00.RAM[2][1] ;
 wire \tms1x00.RAM[2][2] ;
 wire \tms1x00.RAM[2][3] ;
 wire \tms1x00.RAM[30][0] ;
 wire \tms1x00.RAM[30][1] ;
 wire \tms1x00.RAM[30][2] ;
 wire \tms1x00.RAM[30][3] ;
 wire \tms1x00.RAM[31][0] ;
 wire \tms1x00.RAM[31][1] ;
 wire \tms1x00.RAM[31][2] ;
 wire \tms1x00.RAM[31][3] ;
 wire \tms1x00.RAM[32][0] ;
 wire \tms1x00.RAM[32][1] ;
 wire \tms1x00.RAM[32][2] ;
 wire \tms1x00.RAM[32][3] ;
 wire \tms1x00.RAM[33][0] ;
 wire \tms1x00.RAM[33][1] ;
 wire \tms1x00.RAM[33][2] ;
 wire \tms1x00.RAM[33][3] ;
 wire \tms1x00.RAM[34][0] ;
 wire \tms1x00.RAM[34][1] ;
 wire \tms1x00.RAM[34][2] ;
 wire \tms1x00.RAM[34][3] ;
 wire \tms1x00.RAM[35][0] ;
 wire \tms1x00.RAM[35][1] ;
 wire \tms1x00.RAM[35][2] ;
 wire \tms1x00.RAM[35][3] ;
 wire \tms1x00.RAM[36][0] ;
 wire \tms1x00.RAM[36][1] ;
 wire \tms1x00.RAM[36][2] ;
 wire \tms1x00.RAM[36][3] ;
 wire \tms1x00.RAM[37][0] ;
 wire \tms1x00.RAM[37][1] ;
 wire \tms1x00.RAM[37][2] ;
 wire \tms1x00.RAM[37][3] ;
 wire \tms1x00.RAM[38][0] ;
 wire \tms1x00.RAM[38][1] ;
 wire \tms1x00.RAM[38][2] ;
 wire \tms1x00.RAM[38][3] ;
 wire \tms1x00.RAM[39][0] ;
 wire \tms1x00.RAM[39][1] ;
 wire \tms1x00.RAM[39][2] ;
 wire \tms1x00.RAM[39][3] ;
 wire \tms1x00.RAM[3][0] ;
 wire \tms1x00.RAM[3][1] ;
 wire \tms1x00.RAM[3][2] ;
 wire \tms1x00.RAM[3][3] ;
 wire \tms1x00.RAM[40][0] ;
 wire \tms1x00.RAM[40][1] ;
 wire \tms1x00.RAM[40][2] ;
 wire \tms1x00.RAM[40][3] ;
 wire \tms1x00.RAM[41][0] ;
 wire \tms1x00.RAM[41][1] ;
 wire \tms1x00.RAM[41][2] ;
 wire \tms1x00.RAM[41][3] ;
 wire \tms1x00.RAM[42][0] ;
 wire \tms1x00.RAM[42][1] ;
 wire \tms1x00.RAM[42][2] ;
 wire \tms1x00.RAM[42][3] ;
 wire \tms1x00.RAM[43][0] ;
 wire \tms1x00.RAM[43][1] ;
 wire \tms1x00.RAM[43][2] ;
 wire \tms1x00.RAM[43][3] ;
 wire \tms1x00.RAM[44][0] ;
 wire \tms1x00.RAM[44][1] ;
 wire \tms1x00.RAM[44][2] ;
 wire \tms1x00.RAM[44][3] ;
 wire \tms1x00.RAM[45][0] ;
 wire \tms1x00.RAM[45][1] ;
 wire \tms1x00.RAM[45][2] ;
 wire \tms1x00.RAM[45][3] ;
 wire \tms1x00.RAM[46][0] ;
 wire \tms1x00.RAM[46][1] ;
 wire \tms1x00.RAM[46][2] ;
 wire \tms1x00.RAM[46][3] ;
 wire \tms1x00.RAM[47][0] ;
 wire \tms1x00.RAM[47][1] ;
 wire \tms1x00.RAM[47][2] ;
 wire \tms1x00.RAM[47][3] ;
 wire \tms1x00.RAM[48][0] ;
 wire \tms1x00.RAM[48][1] ;
 wire \tms1x00.RAM[48][2] ;
 wire \tms1x00.RAM[48][3] ;
 wire \tms1x00.RAM[49][0] ;
 wire \tms1x00.RAM[49][1] ;
 wire \tms1x00.RAM[49][2] ;
 wire \tms1x00.RAM[49][3] ;
 wire \tms1x00.RAM[4][0] ;
 wire \tms1x00.RAM[4][1] ;
 wire \tms1x00.RAM[4][2] ;
 wire \tms1x00.RAM[4][3] ;
 wire \tms1x00.RAM[50][0] ;
 wire \tms1x00.RAM[50][1] ;
 wire \tms1x00.RAM[50][2] ;
 wire \tms1x00.RAM[50][3] ;
 wire \tms1x00.RAM[51][0] ;
 wire \tms1x00.RAM[51][1] ;
 wire \tms1x00.RAM[51][2] ;
 wire \tms1x00.RAM[51][3] ;
 wire \tms1x00.RAM[52][0] ;
 wire \tms1x00.RAM[52][1] ;
 wire \tms1x00.RAM[52][2] ;
 wire \tms1x00.RAM[52][3] ;
 wire \tms1x00.RAM[53][0] ;
 wire \tms1x00.RAM[53][1] ;
 wire \tms1x00.RAM[53][2] ;
 wire \tms1x00.RAM[53][3] ;
 wire \tms1x00.RAM[54][0] ;
 wire \tms1x00.RAM[54][1] ;
 wire \tms1x00.RAM[54][2] ;
 wire \tms1x00.RAM[54][3] ;
 wire \tms1x00.RAM[55][0] ;
 wire \tms1x00.RAM[55][1] ;
 wire \tms1x00.RAM[55][2] ;
 wire \tms1x00.RAM[55][3] ;
 wire \tms1x00.RAM[56][0] ;
 wire \tms1x00.RAM[56][1] ;
 wire \tms1x00.RAM[56][2] ;
 wire \tms1x00.RAM[56][3] ;
 wire \tms1x00.RAM[57][0] ;
 wire \tms1x00.RAM[57][1] ;
 wire \tms1x00.RAM[57][2] ;
 wire \tms1x00.RAM[57][3] ;
 wire \tms1x00.RAM[58][0] ;
 wire \tms1x00.RAM[58][1] ;
 wire \tms1x00.RAM[58][2] ;
 wire \tms1x00.RAM[58][3] ;
 wire \tms1x00.RAM[59][0] ;
 wire \tms1x00.RAM[59][1] ;
 wire \tms1x00.RAM[59][2] ;
 wire \tms1x00.RAM[59][3] ;
 wire \tms1x00.RAM[5][0] ;
 wire \tms1x00.RAM[5][1] ;
 wire \tms1x00.RAM[5][2] ;
 wire \tms1x00.RAM[5][3] ;
 wire \tms1x00.RAM[60][0] ;
 wire \tms1x00.RAM[60][1] ;
 wire \tms1x00.RAM[60][2] ;
 wire \tms1x00.RAM[60][3] ;
 wire \tms1x00.RAM[61][0] ;
 wire \tms1x00.RAM[61][1] ;
 wire \tms1x00.RAM[61][2] ;
 wire \tms1x00.RAM[61][3] ;
 wire \tms1x00.RAM[62][0] ;
 wire \tms1x00.RAM[62][1] ;
 wire \tms1x00.RAM[62][2] ;
 wire \tms1x00.RAM[62][3] ;
 wire \tms1x00.RAM[63][0] ;
 wire \tms1x00.RAM[63][1] ;
 wire \tms1x00.RAM[63][2] ;
 wire \tms1x00.RAM[63][3] ;
 wire \tms1x00.RAM[64][0] ;
 wire \tms1x00.RAM[64][1] ;
 wire \tms1x00.RAM[64][2] ;
 wire \tms1x00.RAM[64][3] ;
 wire \tms1x00.RAM[65][0] ;
 wire \tms1x00.RAM[65][1] ;
 wire \tms1x00.RAM[65][2] ;
 wire \tms1x00.RAM[65][3] ;
 wire \tms1x00.RAM[66][0] ;
 wire \tms1x00.RAM[66][1] ;
 wire \tms1x00.RAM[66][2] ;
 wire \tms1x00.RAM[66][3] ;
 wire \tms1x00.RAM[67][0] ;
 wire \tms1x00.RAM[67][1] ;
 wire \tms1x00.RAM[67][2] ;
 wire \tms1x00.RAM[67][3] ;
 wire \tms1x00.RAM[68][0] ;
 wire \tms1x00.RAM[68][1] ;
 wire \tms1x00.RAM[68][2] ;
 wire \tms1x00.RAM[68][3] ;
 wire \tms1x00.RAM[69][0] ;
 wire \tms1x00.RAM[69][1] ;
 wire \tms1x00.RAM[69][2] ;
 wire \tms1x00.RAM[69][3] ;
 wire \tms1x00.RAM[6][0] ;
 wire \tms1x00.RAM[6][1] ;
 wire \tms1x00.RAM[6][2] ;
 wire \tms1x00.RAM[6][3] ;
 wire \tms1x00.RAM[70][0] ;
 wire \tms1x00.RAM[70][1] ;
 wire \tms1x00.RAM[70][2] ;
 wire \tms1x00.RAM[70][3] ;
 wire \tms1x00.RAM[71][0] ;
 wire \tms1x00.RAM[71][1] ;
 wire \tms1x00.RAM[71][2] ;
 wire \tms1x00.RAM[71][3] ;
 wire \tms1x00.RAM[72][0] ;
 wire \tms1x00.RAM[72][1] ;
 wire \tms1x00.RAM[72][2] ;
 wire \tms1x00.RAM[72][3] ;
 wire \tms1x00.RAM[73][0] ;
 wire \tms1x00.RAM[73][1] ;
 wire \tms1x00.RAM[73][2] ;
 wire \tms1x00.RAM[73][3] ;
 wire \tms1x00.RAM[74][0] ;
 wire \tms1x00.RAM[74][1] ;
 wire \tms1x00.RAM[74][2] ;
 wire \tms1x00.RAM[74][3] ;
 wire \tms1x00.RAM[75][0] ;
 wire \tms1x00.RAM[75][1] ;
 wire \tms1x00.RAM[75][2] ;
 wire \tms1x00.RAM[75][3] ;
 wire \tms1x00.RAM[76][0] ;
 wire \tms1x00.RAM[76][1] ;
 wire \tms1x00.RAM[76][2] ;
 wire \tms1x00.RAM[76][3] ;
 wire \tms1x00.RAM[77][0] ;
 wire \tms1x00.RAM[77][1] ;
 wire \tms1x00.RAM[77][2] ;
 wire \tms1x00.RAM[77][3] ;
 wire \tms1x00.RAM[78][0] ;
 wire \tms1x00.RAM[78][1] ;
 wire \tms1x00.RAM[78][2] ;
 wire \tms1x00.RAM[78][3] ;
 wire \tms1x00.RAM[79][0] ;
 wire \tms1x00.RAM[79][1] ;
 wire \tms1x00.RAM[79][2] ;
 wire \tms1x00.RAM[79][3] ;
 wire \tms1x00.RAM[7][0] ;
 wire \tms1x00.RAM[7][1] ;
 wire \tms1x00.RAM[7][2] ;
 wire \tms1x00.RAM[7][3] ;
 wire \tms1x00.RAM[80][0] ;
 wire \tms1x00.RAM[80][1] ;
 wire \tms1x00.RAM[80][2] ;
 wire \tms1x00.RAM[80][3] ;
 wire \tms1x00.RAM[81][0] ;
 wire \tms1x00.RAM[81][1] ;
 wire \tms1x00.RAM[81][2] ;
 wire \tms1x00.RAM[81][3] ;
 wire \tms1x00.RAM[82][0] ;
 wire \tms1x00.RAM[82][1] ;
 wire \tms1x00.RAM[82][2] ;
 wire \tms1x00.RAM[82][3] ;
 wire \tms1x00.RAM[83][0] ;
 wire \tms1x00.RAM[83][1] ;
 wire \tms1x00.RAM[83][2] ;
 wire \tms1x00.RAM[83][3] ;
 wire \tms1x00.RAM[84][0] ;
 wire \tms1x00.RAM[84][1] ;
 wire \tms1x00.RAM[84][2] ;
 wire \tms1x00.RAM[84][3] ;
 wire \tms1x00.RAM[85][0] ;
 wire \tms1x00.RAM[85][1] ;
 wire \tms1x00.RAM[85][2] ;
 wire \tms1x00.RAM[85][3] ;
 wire \tms1x00.RAM[86][0] ;
 wire \tms1x00.RAM[86][1] ;
 wire \tms1x00.RAM[86][2] ;
 wire \tms1x00.RAM[86][3] ;
 wire \tms1x00.RAM[87][0] ;
 wire \tms1x00.RAM[87][1] ;
 wire \tms1x00.RAM[87][2] ;
 wire \tms1x00.RAM[87][3] ;
 wire \tms1x00.RAM[88][0] ;
 wire \tms1x00.RAM[88][1] ;
 wire \tms1x00.RAM[88][2] ;
 wire \tms1x00.RAM[88][3] ;
 wire \tms1x00.RAM[89][0] ;
 wire \tms1x00.RAM[89][1] ;
 wire \tms1x00.RAM[89][2] ;
 wire \tms1x00.RAM[89][3] ;
 wire \tms1x00.RAM[8][0] ;
 wire \tms1x00.RAM[8][1] ;
 wire \tms1x00.RAM[8][2] ;
 wire \tms1x00.RAM[8][3] ;
 wire \tms1x00.RAM[90][0] ;
 wire \tms1x00.RAM[90][1] ;
 wire \tms1x00.RAM[90][2] ;
 wire \tms1x00.RAM[90][3] ;
 wire \tms1x00.RAM[91][0] ;
 wire \tms1x00.RAM[91][1] ;
 wire \tms1x00.RAM[91][2] ;
 wire \tms1x00.RAM[91][3] ;
 wire \tms1x00.RAM[92][0] ;
 wire \tms1x00.RAM[92][1] ;
 wire \tms1x00.RAM[92][2] ;
 wire \tms1x00.RAM[92][3] ;
 wire \tms1x00.RAM[93][0] ;
 wire \tms1x00.RAM[93][1] ;
 wire \tms1x00.RAM[93][2] ;
 wire \tms1x00.RAM[93][3] ;
 wire \tms1x00.RAM[94][0] ;
 wire \tms1x00.RAM[94][1] ;
 wire \tms1x00.RAM[94][2] ;
 wire \tms1x00.RAM[94][3] ;
 wire \tms1x00.RAM[95][0] ;
 wire \tms1x00.RAM[95][1] ;
 wire \tms1x00.RAM[95][2] ;
 wire \tms1x00.RAM[95][3] ;
 wire \tms1x00.RAM[96][0] ;
 wire \tms1x00.RAM[96][1] ;
 wire \tms1x00.RAM[96][2] ;
 wire \tms1x00.RAM[96][3] ;
 wire \tms1x00.RAM[97][0] ;
 wire \tms1x00.RAM[97][1] ;
 wire \tms1x00.RAM[97][2] ;
 wire \tms1x00.RAM[97][3] ;
 wire \tms1x00.RAM[98][0] ;
 wire \tms1x00.RAM[98][1] ;
 wire \tms1x00.RAM[98][2] ;
 wire \tms1x00.RAM[98][3] ;
 wire \tms1x00.RAM[99][0] ;
 wire \tms1x00.RAM[99][1] ;
 wire \tms1x00.RAM[99][2] ;
 wire \tms1x00.RAM[99][3] ;
 wire \tms1x00.RAM[9][0] ;
 wire \tms1x00.RAM[9][1] ;
 wire \tms1x00.RAM[9][2] ;
 wire \tms1x00.RAM[9][3] ;
 wire \tms1x00.SR[0] ;
 wire \tms1x00.SR[1] ;
 wire \tms1x00.SR[2] ;
 wire \tms1x00.SR[3] ;
 wire \tms1x00.SR[4] ;
 wire \tms1x00.SR[5] ;
 wire \tms1x00.X[0] ;
 wire \tms1x00.X[1] ;
 wire \tms1x00.X[2] ;
 wire \tms1x00.Y[0] ;
 wire \tms1x00.Y[1] ;
 wire \tms1x00.Y[2] ;
 wire \tms1x00.Y[3] ;
 wire \tms1x00.ins_in[0] ;
 wire \tms1x00.ins_in[1] ;
 wire \tms1x00.ins_in[2] ;
 wire \tms1x00.ins_in[3] ;
 wire \tms1x00.ins_in[4] ;
 wire \tms1x00.ins_in[5] ;
 wire \tms1x00.ins_in[6] ;
 wire \tms1x00.ins_in[7] ;
 wire \tms1x00.ram_addr_buff[0] ;
 wire \tms1x00.ram_addr_buff[1] ;
 wire \tms1x00.ram_addr_buff[2] ;
 wire \tms1x00.ram_addr_buff[3] ;
 wire \tms1x00.ram_addr_buff[4] ;
 wire \tms1x00.ram_addr_buff[5] ;
 wire \tms1x00.ram_addr_buff[6] ;
 wire \tms1x00.rom_addr[0] ;
 wire \tms1x00.rom_addr[1] ;
 wire \tms1x00.status ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire clknet_leaf_1_wb_clk_i;
 wire clknet_leaf_2_wb_clk_i;
 wire clknet_leaf_3_wb_clk_i;
 wire clknet_leaf_4_wb_clk_i;
 wire clknet_leaf_5_wb_clk_i;
 wire clknet_leaf_6_wb_clk_i;
 wire clknet_leaf_7_wb_clk_i;
 wire clknet_leaf_8_wb_clk_i;
 wire clknet_leaf_9_wb_clk_i;
 wire clknet_leaf_10_wb_clk_i;
 wire clknet_leaf_11_wb_clk_i;
 wire clknet_leaf_12_wb_clk_i;
 wire clknet_leaf_13_wb_clk_i;
 wire clknet_leaf_14_wb_clk_i;
 wire clknet_leaf_15_wb_clk_i;
 wire clknet_leaf_16_wb_clk_i;
 wire clknet_leaf_17_wb_clk_i;
 wire clknet_leaf_18_wb_clk_i;
 wire clknet_leaf_19_wb_clk_i;
 wire clknet_leaf_20_wb_clk_i;
 wire clknet_leaf_21_wb_clk_i;
 wire clknet_leaf_22_wb_clk_i;
 wire clknet_leaf_23_wb_clk_i;
 wire clknet_leaf_24_wb_clk_i;
 wire clknet_leaf_25_wb_clk_i;
 wire clknet_leaf_26_wb_clk_i;
 wire clknet_leaf_27_wb_clk_i;
 wire clknet_leaf_28_wb_clk_i;
 wire clknet_leaf_29_wb_clk_i;
 wire clknet_leaf_30_wb_clk_i;
 wire clknet_leaf_31_wb_clk_i;
 wire clknet_leaf_32_wb_clk_i;
 wire clknet_leaf_33_wb_clk_i;
 wire clknet_leaf_34_wb_clk_i;
 wire clknet_leaf_35_wb_clk_i;
 wire clknet_leaf_36_wb_clk_i;
 wire clknet_leaf_37_wb_clk_i;
 wire clknet_leaf_38_wb_clk_i;
 wire clknet_leaf_39_wb_clk_i;
 wire clknet_leaf_40_wb_clk_i;
 wire clknet_leaf_41_wb_clk_i;
 wire clknet_leaf_42_wb_clk_i;
 wire clknet_0_wb_clk_i;
 wire clknet_2_0__leaf_wb_clk_i;
 wire clknet_2_1__leaf_wb_clk_i;
 wire clknet_2_2__leaf_wb_clk_i;
 wire clknet_2_3__leaf_wb_clk_i;

 sky130_fd_sc_hd__and3_1 _2089_ (.A(net30),
    .B(net28),
    .C(net31),
    .X(_0618_));
 sky130_fd_sc_hd__clkbuf_1 _2090_ (.A(_0618_),
    .X(_0000_));
 sky130_fd_sc_hd__clkbuf_4 _2091_ (.A(\tms1x00.Y[0] ),
    .X(_0619_));
 sky130_fd_sc_hd__buf_2 _2092_ (.A(\tms1x00.ram_addr_buff[0] ),
    .X(_0620_));
 sky130_fd_sc_hd__inv_2 _2093_ (.A(net16),
    .Y(_0621_));
 sky130_fd_sc_hd__nand2b_1 _2094_ (.A_N(net37),
    .B(net39),
    .Y(_0622_));
 sky130_fd_sc_hd__nor2_4 _2095_ (.A(net38),
    .B(_0622_),
    .Y(_0623_));
 sky130_fd_sc_hd__nand2_2 _2096_ (.A(_0621_),
    .B(_0623_),
    .Y(_0624_));
 sky130_fd_sc_hd__clkbuf_4 _2097_ (.A(_0624_),
    .X(_0625_));
 sky130_fd_sc_hd__mux2_1 _2098_ (.A0(_0619_),
    .A1(_0620_),
    .S(_0625_),
    .X(_0626_));
 sky130_fd_sc_hd__clkbuf_1 _2099_ (.A(_0626_),
    .X(_0008_));
 sky130_fd_sc_hd__clkbuf_4 _2100_ (.A(\tms1x00.Y[1] ),
    .X(_0627_));
 sky130_fd_sc_hd__buf_2 _2101_ (.A(\tms1x00.ram_addr_buff[1] ),
    .X(_0628_));
 sky130_fd_sc_hd__mux2_1 _2102_ (.A0(_0627_),
    .A1(_0628_),
    .S(_0625_),
    .X(_0629_));
 sky130_fd_sc_hd__clkbuf_1 _2103_ (.A(_0629_),
    .X(_0009_));
 sky130_fd_sc_hd__buf_2 _2104_ (.A(\tms1x00.Y[2] ),
    .X(_0630_));
 sky130_fd_sc_hd__mux2_1 _2105_ (.A0(_0630_),
    .A1(\tms1x00.ram_addr_buff[2] ),
    .S(_0625_),
    .X(_0631_));
 sky130_fd_sc_hd__clkbuf_1 _2106_ (.A(_0631_),
    .X(_0010_));
 sky130_fd_sc_hd__clkbuf_4 _2107_ (.A(\tms1x00.Y[3] ),
    .X(_0632_));
 sky130_fd_sc_hd__clkbuf_4 _2108_ (.A(_0632_),
    .X(_0633_));
 sky130_fd_sc_hd__mux2_1 _2109_ (.A0(_0633_),
    .A1(\tms1x00.ram_addr_buff[3] ),
    .S(_0625_),
    .X(_0634_));
 sky130_fd_sc_hd__clkbuf_1 _2110_ (.A(_0634_),
    .X(_0011_));
 sky130_fd_sc_hd__buf_4 _2111_ (.A(\tms1x00.ram_addr_buff[4] ),
    .X(_0635_));
 sky130_fd_sc_hd__mux2_1 _2112_ (.A0(\tms1x00.X[2] ),
    .A1(_0635_),
    .S(_0625_),
    .X(_0636_));
 sky130_fd_sc_hd__clkbuf_1 _2113_ (.A(_0636_),
    .X(_0012_));
 sky130_fd_sc_hd__clkbuf_8 _2114_ (.A(\tms1x00.ram_addr_buff[5] ),
    .X(_0637_));
 sky130_fd_sc_hd__mux2_1 _2115_ (.A0(\tms1x00.X[0] ),
    .A1(_0637_),
    .S(_0625_),
    .X(_0638_));
 sky130_fd_sc_hd__clkbuf_1 _2116_ (.A(_0638_),
    .X(_0013_));
 sky130_fd_sc_hd__buf_4 _2117_ (.A(\tms1x00.ram_addr_buff[6] ),
    .X(_0639_));
 sky130_fd_sc_hd__mux2_1 _2118_ (.A0(\tms1x00.X[1] ),
    .A1(_0639_),
    .S(_0625_),
    .X(_0640_));
 sky130_fd_sc_hd__clkbuf_1 _2119_ (.A(_0640_),
    .X(_0014_));
 sky130_fd_sc_hd__inv_2 _2120_ (.A(net31),
    .Y(net76));
 sky130_fd_sc_hd__nand3_2 _2121_ (.A(net30),
    .B(net28),
    .C(net18),
    .Y(net75));
 sky130_fd_sc_hd__or3_1 _2122_ (.A(_0630_),
    .B(_0627_),
    .C(_0619_),
    .X(_0641_));
 sky130_fd_sc_hd__clkbuf_4 _2123_ (.A(\tms1x00.ins_in[7] ),
    .X(_0642_));
 sky130_fd_sc_hd__clkbuf_4 _2124_ (.A(\tms1x00.ins_in[6] ),
    .X(_0643_));
 sky130_fd_sc_hd__or4_1 _2125_ (.A(\tms1x00.ins_in[3] ),
    .B(\tms1x00.ins_in[2] ),
    .C(\tms1x00.ins_in[1] ),
    .D(\tms1x00.ins_in[0] ),
    .X(_0644_));
 sky130_fd_sc_hd__nand2_1 _2126_ (.A(\tms1x00.ins_in[5] ),
    .B(\tms1x00.ins_in[4] ),
    .Y(_0645_));
 sky130_fd_sc_hd__or2_2 _2127_ (.A(_0644_),
    .B(_0645_),
    .X(_0646_));
 sky130_fd_sc_hd__nand3b_2 _2128_ (.A_N(net39),
    .B(net37),
    .C(net38),
    .Y(_0647_));
 sky130_fd_sc_hd__or4_4 _2129_ (.A(_0642_),
    .B(_0643_),
    .C(_0646_),
    .D(_0647_),
    .X(_0648_));
 sky130_fd_sc_hd__clkbuf_4 _2130_ (.A(_0648_),
    .X(_0649_));
 sky130_fd_sc_hd__inv_2 _2131_ (.A(\tms1x00.Y[3] ),
    .Y(_0650_));
 sky130_fd_sc_hd__buf_2 _2132_ (.A(_0650_),
    .X(_0651_));
 sky130_fd_sc_hd__nor3_1 _2133_ (.A(_0630_),
    .B(_0627_),
    .C(_0619_),
    .Y(_0652_));
 sky130_fd_sc_hd__or2b_1 _2134_ (.A(\tms1x00.ins_in[6] ),
    .B_N(\tms1x00.ins_in[7] ),
    .X(_0653_));
 sky130_fd_sc_hd__or2_2 _2135_ (.A(_0647_),
    .B(_0653_),
    .X(_0654_));
 sky130_fd_sc_hd__nor2_4 _2136_ (.A(_0646_),
    .B(_0654_),
    .Y(_0655_));
 sky130_fd_sc_hd__clkbuf_4 _2137_ (.A(_0655_),
    .X(_0656_));
 sky130_fd_sc_hd__a31o_1 _2138_ (.A1(_0651_),
    .A2(_0652_),
    .A3(_0656_),
    .B1(net40),
    .X(_0657_));
 sky130_fd_sc_hd__buf_2 _2139_ (.A(_0621_),
    .X(_0658_));
 sky130_fd_sc_hd__o311a_1 _2140_ (.A1(_0633_),
    .A2(_0641_),
    .A3(_0649_),
    .B1(_0657_),
    .C1(_0658_),
    .X(_0015_));
 sky130_fd_sc_hd__and4b_1 _2141_ (.A_N(\tms1x00.ins_in[5] ),
    .B(\tms1x00.ins_in[4] ),
    .C(\tms1x00.ins_in[7] ),
    .D(\tms1x00.ins_in[6] ),
    .X(_0659_));
 sky130_fd_sc_hd__nand3b_1 _2142_ (.A_N(\tms1x00.ins_in[3] ),
    .B(\tms1x00.ins_in[2] ),
    .C(_0659_),
    .Y(_0660_));
 sky130_fd_sc_hd__or3b_1 _2143_ (.A(\tms1x00.ins_in[1] ),
    .B(net37),
    .C_N(net38),
    .X(_0661_));
 sky130_fd_sc_hd__or4_2 _2144_ (.A(net39),
    .B(net16),
    .C(_0660_),
    .D(_0661_),
    .X(_0662_));
 sky130_fd_sc_hd__buf_2 _2145_ (.A(_0006_),
    .X(_0663_));
 sky130_fd_sc_hd__buf_6 _2146_ (.A(_0002_),
    .X(_0664_));
 sky130_fd_sc_hd__buf_4 _2147_ (.A(_0664_),
    .X(_0665_));
 sky130_fd_sc_hd__clkbuf_4 _2148_ (.A(_0665_),
    .X(_0666_));
 sky130_fd_sc_hd__buf_6 _2149_ (.A(_0001_),
    .X(_0667_));
 sky130_fd_sc_hd__mux2_1 _2150_ (.A0(\tms1x00.RAM[92][0] ),
    .A1(\tms1x00.RAM[93][0] ),
    .S(_0667_),
    .X(_0668_));
 sky130_fd_sc_hd__inv_2 _2151_ (.A(_0668_),
    .Y(_0669_));
 sky130_fd_sc_hd__buf_2 _2152_ (.A(_0665_),
    .X(_0670_));
 sky130_fd_sc_hd__buf_6 _2153_ (.A(_0001_),
    .X(_0671_));
 sky130_fd_sc_hd__buf_4 _2154_ (.A(_0671_),
    .X(_0672_));
 sky130_fd_sc_hd__mux2_1 _2155_ (.A0(\tms1x00.RAM[94][0] ),
    .A1(\tms1x00.RAM[95][0] ),
    .S(_0672_),
    .X(_0673_));
 sky130_fd_sc_hd__nand2_1 _2156_ (.A(_0670_),
    .B(_0673_),
    .Y(_0674_));
 sky130_fd_sc_hd__buf_2 _2157_ (.A(_0003_),
    .X(_0675_));
 sky130_fd_sc_hd__o211a_1 _2158_ (.A1(_0666_),
    .A2(_0669_),
    .B1(_0674_),
    .C1(_0675_),
    .X(_0676_));
 sky130_fd_sc_hd__clkbuf_4 _2159_ (.A(_0003_),
    .X(_0677_));
 sky130_fd_sc_hd__clkbuf_4 _2160_ (.A(_0677_),
    .X(_0678_));
 sky130_fd_sc_hd__buf_6 _2161_ (.A(_0671_),
    .X(_0679_));
 sky130_fd_sc_hd__clkbuf_8 _2162_ (.A(_0664_),
    .X(_0680_));
 sky130_fd_sc_hd__mux4_2 _2163_ (.A0(\tms1x00.RAM[88][0] ),
    .A1(\tms1x00.RAM[89][0] ),
    .A2(\tms1x00.RAM[90][0] ),
    .A3(\tms1x00.RAM[91][0] ),
    .S0(_0679_),
    .S1(_0680_),
    .X(_0681_));
 sky130_fd_sc_hd__buf_2 _2164_ (.A(_0004_),
    .X(_0682_));
 sky130_fd_sc_hd__o21ai_1 _2165_ (.A1(_0678_),
    .A2(_0681_),
    .B1(_0682_),
    .Y(_0683_));
 sky130_fd_sc_hd__buf_2 _2166_ (.A(_0677_),
    .X(_0684_));
 sky130_fd_sc_hd__buf_6 _2167_ (.A(_0001_),
    .X(_0685_));
 sky130_fd_sc_hd__buf_6 _2168_ (.A(_0685_),
    .X(_0686_));
 sky130_fd_sc_hd__clkbuf_8 _2169_ (.A(_0002_),
    .X(_0687_));
 sky130_fd_sc_hd__buf_6 _2170_ (.A(_0687_),
    .X(_0688_));
 sky130_fd_sc_hd__mux4_1 _2171_ (.A0(\tms1x00.RAM[80][0] ),
    .A1(\tms1x00.RAM[81][0] ),
    .A2(\tms1x00.RAM[82][0] ),
    .A3(\tms1x00.RAM[83][0] ),
    .S0(_0686_),
    .S1(_0688_),
    .X(_0689_));
 sky130_fd_sc_hd__nor2_1 _2172_ (.A(_0684_),
    .B(_0689_),
    .Y(_0690_));
 sky130_fd_sc_hd__inv_2 _2173_ (.A(_0003_),
    .Y(_0691_));
 sky130_fd_sc_hd__clkbuf_4 _2174_ (.A(_0691_),
    .X(_0692_));
 sky130_fd_sc_hd__buf_6 _2175_ (.A(_0667_),
    .X(_0693_));
 sky130_fd_sc_hd__buf_4 _2176_ (.A(_0664_),
    .X(_0694_));
 sky130_fd_sc_hd__mux4_1 _2177_ (.A0(\tms1x00.RAM[84][0] ),
    .A1(\tms1x00.RAM[85][0] ),
    .A2(\tms1x00.RAM[86][0] ),
    .A3(\tms1x00.RAM[87][0] ),
    .S0(_0693_),
    .S1(_0694_),
    .X(_0695_));
 sky130_fd_sc_hd__inv_2 _2178_ (.A(_0004_),
    .Y(_0696_));
 sky130_fd_sc_hd__clkbuf_4 _2179_ (.A(_0696_),
    .X(_0697_));
 sky130_fd_sc_hd__o21ai_1 _2180_ (.A1(_0692_),
    .A2(_0695_),
    .B1(_0697_),
    .Y(_0698_));
 sky130_fd_sc_hd__buf_2 _2181_ (.A(_0005_),
    .X(_0699_));
 sky130_fd_sc_hd__o221a_1 _2182_ (.A1(_0676_),
    .A2(_0683_),
    .B1(_0690_),
    .B2(_0698_),
    .C1(_0699_),
    .X(_0700_));
 sky130_fd_sc_hd__buf_2 _2183_ (.A(_0005_),
    .X(_0701_));
 sky130_fd_sc_hd__buf_6 _2184_ (.A(_0002_),
    .X(_0702_));
 sky130_fd_sc_hd__buf_4 _2185_ (.A(_0702_),
    .X(_0703_));
 sky130_fd_sc_hd__buf_6 _2186_ (.A(_0671_),
    .X(_0704_));
 sky130_fd_sc_hd__mux2_1 _2187_ (.A0(\tms1x00.RAM[76][0] ),
    .A1(\tms1x00.RAM[77][0] ),
    .S(_0704_),
    .X(_0705_));
 sky130_fd_sc_hd__and2b_1 _2188_ (.A_N(_0703_),
    .B(_0705_),
    .X(_0706_));
 sky130_fd_sc_hd__buf_6 _2189_ (.A(_0002_),
    .X(_0707_));
 sky130_fd_sc_hd__clkbuf_4 _2190_ (.A(_0707_),
    .X(_0708_));
 sky130_fd_sc_hd__buf_6 _2191_ (.A(_0671_),
    .X(_0709_));
 sky130_fd_sc_hd__mux2_1 _2192_ (.A0(\tms1x00.RAM[78][0] ),
    .A1(\tms1x00.RAM[79][0] ),
    .S(_0709_),
    .X(_0710_));
 sky130_fd_sc_hd__clkbuf_4 _2193_ (.A(_0691_),
    .X(_0711_));
 sky130_fd_sc_hd__a21o_1 _2194_ (.A1(_0708_),
    .A2(_0710_),
    .B1(_0711_),
    .X(_0712_));
 sky130_fd_sc_hd__mux4_2 _2195_ (.A0(\tms1x00.RAM[72][0] ),
    .A1(\tms1x00.RAM[73][0] ),
    .A2(\tms1x00.RAM[74][0] ),
    .A3(\tms1x00.RAM[75][0] ),
    .S0(_0693_),
    .S1(_0694_),
    .X(_0713_));
 sky130_fd_sc_hd__buf_2 _2196_ (.A(_0677_),
    .X(_0714_));
 sky130_fd_sc_hd__buf_2 _2197_ (.A(_0004_),
    .X(_0715_));
 sky130_fd_sc_hd__o221a_1 _2198_ (.A1(_0706_),
    .A2(_0712_),
    .B1(_0713_),
    .B2(_0714_),
    .C1(_0715_),
    .X(_0716_));
 sky130_fd_sc_hd__mux2_1 _2199_ (.A0(\tms1x00.RAM[68][0] ),
    .A1(\tms1x00.RAM[69][0] ),
    .S(_0672_),
    .X(_0717_));
 sky130_fd_sc_hd__and2b_1 _2200_ (.A_N(_0708_),
    .B(_0717_),
    .X(_0718_));
 sky130_fd_sc_hd__buf_4 _2201_ (.A(_0671_),
    .X(_0719_));
 sky130_fd_sc_hd__mux2_1 _2202_ (.A0(\tms1x00.RAM[70][0] ),
    .A1(\tms1x00.RAM[71][0] ),
    .S(_0719_),
    .X(_0720_));
 sky130_fd_sc_hd__clkbuf_4 _2203_ (.A(_0691_),
    .X(_0721_));
 sky130_fd_sc_hd__a21o_1 _2204_ (.A1(_0670_),
    .A2(_0720_),
    .B1(_0721_),
    .X(_0722_));
 sky130_fd_sc_hd__buf_6 _2205_ (.A(_0001_),
    .X(_0723_));
 sky130_fd_sc_hd__buf_6 _2206_ (.A(_0723_),
    .X(_0724_));
 sky130_fd_sc_hd__mux4_2 _2207_ (.A0(\tms1x00.RAM[64][0] ),
    .A1(\tms1x00.RAM[65][0] ),
    .A2(\tms1x00.RAM[66][0] ),
    .A3(\tms1x00.RAM[67][0] ),
    .S0(_0724_),
    .S1(_0688_),
    .X(_0725_));
 sky130_fd_sc_hd__clkbuf_4 _2208_ (.A(_0003_),
    .X(_0726_));
 sky130_fd_sc_hd__buf_2 _2209_ (.A(_0726_),
    .X(_0727_));
 sky130_fd_sc_hd__clkbuf_4 _2210_ (.A(_0696_),
    .X(_0728_));
 sky130_fd_sc_hd__buf_2 _2211_ (.A(_0728_),
    .X(_0729_));
 sky130_fd_sc_hd__o221a_1 _2212_ (.A1(_0718_),
    .A2(_0722_),
    .B1(_0725_),
    .B2(_0727_),
    .C1(_0729_),
    .X(_0730_));
 sky130_fd_sc_hd__nor3_1 _2213_ (.A(_0701_),
    .B(_0716_),
    .C(_0730_),
    .Y(_0731_));
 sky130_fd_sc_hd__mux2_1 _2214_ (.A0(\tms1x00.RAM[118][0] ),
    .A1(\tms1x00.RAM[119][0] ),
    .S(_0719_),
    .X(_0732_));
 sky130_fd_sc_hd__nand2_1 _2215_ (.A(_0666_),
    .B(_0732_),
    .Y(_0733_));
 sky130_fd_sc_hd__mux2_1 _2216_ (.A0(\tms1x00.RAM[116][0] ),
    .A1(\tms1x00.RAM[117][0] ),
    .S(_0723_),
    .X(_0734_));
 sky130_fd_sc_hd__or2b_1 _2217_ (.A(_0680_),
    .B_N(_0734_),
    .X(_0735_));
 sky130_fd_sc_hd__buf_6 _2218_ (.A(_0002_),
    .X(_0736_));
 sky130_fd_sc_hd__mux4_1 _2219_ (.A0(\tms1x00.RAM[112][0] ),
    .A1(\tms1x00.RAM[113][0] ),
    .A2(\tms1x00.RAM[114][0] ),
    .A3(\tms1x00.RAM[115][0] ),
    .S0(_0723_),
    .S1(_0736_),
    .X(_0737_));
 sky130_fd_sc_hd__o21ai_1 _2220_ (.A1(_0726_),
    .A2(_0737_),
    .B1(_0728_),
    .Y(_0738_));
 sky130_fd_sc_hd__a31o_1 _2221_ (.A1(_0678_),
    .A2(_0733_),
    .A3(_0735_),
    .B1(_0738_),
    .X(_0739_));
 sky130_fd_sc_hd__clkbuf_4 _2222_ (.A(_0711_),
    .X(_0740_));
 sky130_fd_sc_hd__mux4_1 _2223_ (.A0(\tms1x00.RAM[124][0] ),
    .A1(\tms1x00.RAM[125][0] ),
    .A2(\tms1x00.RAM[126][0] ),
    .A3(\tms1x00.RAM[127][0] ),
    .S0(_0724_),
    .S1(_0688_),
    .X(_0741_));
 sky130_fd_sc_hd__clkbuf_4 _2224_ (.A(_0003_),
    .X(_0742_));
 sky130_fd_sc_hd__buf_6 _2225_ (.A(_0001_),
    .X(_0743_));
 sky130_fd_sc_hd__buf_8 _2226_ (.A(_0002_),
    .X(_0744_));
 sky130_fd_sc_hd__mux4_1 _2227_ (.A0(\tms1x00.RAM[120][0] ),
    .A1(\tms1x00.RAM[121][0] ),
    .A2(\tms1x00.RAM[122][0] ),
    .A3(\tms1x00.RAM[123][0] ),
    .S0(_0743_),
    .S1(_0744_),
    .X(_0745_));
 sky130_fd_sc_hd__clkbuf_4 _2228_ (.A(_0004_),
    .X(_0746_));
 sky130_fd_sc_hd__o21a_1 _2229_ (.A1(_0742_),
    .A2(_0745_),
    .B1(_0746_),
    .X(_0747_));
 sky130_fd_sc_hd__o21ai_1 _2230_ (.A1(_0740_),
    .A2(_0741_),
    .B1(_0747_),
    .Y(_0748_));
 sky130_fd_sc_hd__clkinv_2 _2231_ (.A(_0006_),
    .Y(_0749_));
 sky130_fd_sc_hd__buf_6 _2232_ (.A(_0001_),
    .X(_0750_));
 sky130_fd_sc_hd__mux4_2 _2233_ (.A0(\tms1x00.RAM[108][0] ),
    .A1(\tms1x00.RAM[109][0] ),
    .A2(\tms1x00.RAM[110][0] ),
    .A3(\tms1x00.RAM[111][0] ),
    .S0(_0750_),
    .S1(_0702_),
    .X(_0751_));
 sky130_fd_sc_hd__nor2_1 _2234_ (.A(_0721_),
    .B(_0751_),
    .Y(_0752_));
 sky130_fd_sc_hd__mux4_1 _2235_ (.A0(\tms1x00.RAM[104][0] ),
    .A1(\tms1x00.RAM[105][0] ),
    .A2(\tms1x00.RAM[106][0] ),
    .A3(\tms1x00.RAM[107][0] ),
    .S0(_0685_),
    .S1(_0664_),
    .X(_0753_));
 sky130_fd_sc_hd__o21ai_1 _2236_ (.A1(_0677_),
    .A2(_0753_),
    .B1(_0746_),
    .Y(_0754_));
 sky130_fd_sc_hd__buf_6 _2237_ (.A(_0001_),
    .X(_0755_));
 sky130_fd_sc_hd__mux4_1 _2238_ (.A0(\tms1x00.RAM[96][0] ),
    .A1(\tms1x00.RAM[97][0] ),
    .A2(\tms1x00.RAM[98][0] ),
    .A3(\tms1x00.RAM[99][0] ),
    .S0(_0755_),
    .S1(_0744_),
    .X(_0756_));
 sky130_fd_sc_hd__nor2_1 _2239_ (.A(_0742_),
    .B(_0756_),
    .Y(_0757_));
 sky130_fd_sc_hd__clkbuf_4 _2240_ (.A(_0691_),
    .X(_0758_));
 sky130_fd_sc_hd__mux4_2 _2241_ (.A0(\tms1x00.RAM[100][0] ),
    .A1(\tms1x00.RAM[101][0] ),
    .A2(\tms1x00.RAM[102][0] ),
    .A3(\tms1x00.RAM[103][0] ),
    .S0(_0685_),
    .S1(_0736_),
    .X(_0759_));
 sky130_fd_sc_hd__o21ai_1 _2242_ (.A1(_0758_),
    .A2(_0759_),
    .B1(_0728_),
    .Y(_0760_));
 sky130_fd_sc_hd__inv_2 _2243_ (.A(_0005_),
    .Y(_0761_));
 sky130_fd_sc_hd__o221a_1 _2244_ (.A1(_0752_),
    .A2(_0754_),
    .B1(_0757_),
    .B2(_0760_),
    .C1(_0761_),
    .X(_0762_));
 sky130_fd_sc_hd__a311o_1 _2245_ (.A1(_0699_),
    .A2(_0739_),
    .A3(_0748_),
    .B1(_0749_),
    .C1(_0762_),
    .X(_0763_));
 sky130_fd_sc_hd__o311a_2 _2246_ (.A1(_0663_),
    .A2(_0700_),
    .A3(_0731_),
    .B1(_0763_),
    .C1(_0007_),
    .X(_0764_));
 sky130_fd_sc_hd__clkbuf_4 _2247_ (.A(_0665_),
    .X(_0765_));
 sky130_fd_sc_hd__buf_6 _2248_ (.A(_0743_),
    .X(_0766_));
 sky130_fd_sc_hd__mux2_1 _2249_ (.A0(\tms1x00.RAM[6][0] ),
    .A1(\tms1x00.RAM[7][0] ),
    .S(_0766_),
    .X(_0767_));
 sky130_fd_sc_hd__mux2_1 _2250_ (.A0(\tms1x00.RAM[4][0] ),
    .A1(\tms1x00.RAM[5][0] ),
    .S(_0704_),
    .X(_0768_));
 sky130_fd_sc_hd__and2b_1 _2251_ (.A_N(_0703_),
    .B(_0768_),
    .X(_0769_));
 sky130_fd_sc_hd__a211o_1 _2252_ (.A1(_0765_),
    .A2(_0767_),
    .B1(_0769_),
    .C1(_0740_),
    .X(_0770_));
 sky130_fd_sc_hd__mux4_1 _2253_ (.A0(\tms1x00.RAM[0][0] ),
    .A1(\tms1x00.RAM[1][0] ),
    .A2(\tms1x00.RAM[2][0] ),
    .A3(\tms1x00.RAM[3][0] ),
    .S0(_0693_),
    .S1(_0694_),
    .X(_0771_));
 sky130_fd_sc_hd__or2_1 _2254_ (.A(_0714_),
    .B(_0771_),
    .X(_0772_));
 sky130_fd_sc_hd__clkbuf_4 _2255_ (.A(_0744_),
    .X(_0773_));
 sky130_fd_sc_hd__mux2_1 _2256_ (.A0(\tms1x00.RAM[12][0] ),
    .A1(\tms1x00.RAM[13][0] ),
    .S(_0709_),
    .X(_0774_));
 sky130_fd_sc_hd__and2b_1 _2257_ (.A_N(_0773_),
    .B(_0774_),
    .X(_0775_));
 sky130_fd_sc_hd__mux2_1 _2258_ (.A0(\tms1x00.RAM[14][0] ),
    .A1(\tms1x00.RAM[15][0] ),
    .S(_0719_),
    .X(_0776_));
 sky130_fd_sc_hd__a21o_1 _2259_ (.A1(_0670_),
    .A2(_0776_),
    .B1(_0758_),
    .X(_0777_));
 sky130_fd_sc_hd__mux4_1 _2260_ (.A0(\tms1x00.RAM[8][0] ),
    .A1(\tms1x00.RAM[9][0] ),
    .A2(\tms1x00.RAM[10][0] ),
    .A3(\tms1x00.RAM[11][0] ),
    .S0(_0686_),
    .S1(_0688_),
    .X(_0778_));
 sky130_fd_sc_hd__o221a_1 _2261_ (.A1(_0775_),
    .A2(_0777_),
    .B1(_0778_),
    .B2(_0727_),
    .C1(_0715_),
    .X(_0779_));
 sky130_fd_sc_hd__a311oi_1 _2262_ (.A1(_0729_),
    .A2(_0770_),
    .A3(_0772_),
    .B1(_0701_),
    .C1(_0779_),
    .Y(_0780_));
 sky130_fd_sc_hd__buf_4 _2263_ (.A(_0736_),
    .X(_0781_));
 sky130_fd_sc_hd__buf_6 _2264_ (.A(_0671_),
    .X(_0782_));
 sky130_fd_sc_hd__mux2_1 _2265_ (.A0(\tms1x00.RAM[28][0] ),
    .A1(\tms1x00.RAM[29][0] ),
    .S(_0782_),
    .X(_0783_));
 sky130_fd_sc_hd__or2b_1 _2266_ (.A(_0781_),
    .B_N(_0783_),
    .X(_0784_));
 sky130_fd_sc_hd__mux2_1 _2267_ (.A0(\tms1x00.RAM[30][0] ),
    .A1(\tms1x00.RAM[31][0] ),
    .S(_0679_),
    .X(_0785_));
 sky130_fd_sc_hd__nand2_1 _2268_ (.A(_0765_),
    .B(_0785_),
    .Y(_0786_));
 sky130_fd_sc_hd__mux4_1 _2269_ (.A0(\tms1x00.RAM[24][0] ),
    .A1(\tms1x00.RAM[25][0] ),
    .A2(\tms1x00.RAM[26][0] ),
    .A3(\tms1x00.RAM[27][0] ),
    .S0(_0743_),
    .S1(_0744_),
    .X(_0787_));
 sky130_fd_sc_hd__o21ai_1 _2270_ (.A1(_0742_),
    .A2(_0787_),
    .B1(_0682_),
    .Y(_0788_));
 sky130_fd_sc_hd__a31o_1 _2271_ (.A1(_0714_),
    .A2(_0784_),
    .A3(_0786_),
    .B1(_0788_),
    .X(_0789_));
 sky130_fd_sc_hd__mux4_1 _2272_ (.A0(\tms1x00.RAM[16][0] ),
    .A1(\tms1x00.RAM[17][0] ),
    .A2(\tms1x00.RAM[18][0] ),
    .A3(\tms1x00.RAM[19][0] ),
    .S0(_0766_),
    .S1(_0708_),
    .X(_0790_));
 sky130_fd_sc_hd__mux4_1 _2273_ (.A0(\tms1x00.RAM[20][0] ),
    .A1(\tms1x00.RAM[21][0] ),
    .A2(\tms1x00.RAM[22][0] ),
    .A3(\tms1x00.RAM[23][0] ),
    .S0(_0709_),
    .S1(_0665_),
    .X(_0791_));
 sky130_fd_sc_hd__o21a_1 _2274_ (.A1(_0692_),
    .A2(_0791_),
    .B1(_0697_),
    .X(_0792_));
 sky130_fd_sc_hd__o21ai_1 _2275_ (.A1(_0727_),
    .A2(_0790_),
    .B1(_0792_),
    .Y(_0793_));
 sky130_fd_sc_hd__a31o_1 _2276_ (.A1(_0701_),
    .A2(_0789_),
    .A3(_0793_),
    .B1(_0663_),
    .X(_0794_));
 sky130_fd_sc_hd__mux2_1 _2277_ (.A0(\tms1x00.RAM[54][0] ),
    .A1(\tms1x00.RAM[55][0] ),
    .S(_0679_),
    .X(_0795_));
 sky130_fd_sc_hd__nand2_1 _2278_ (.A(_0765_),
    .B(_0795_),
    .Y(_0796_));
 sky130_fd_sc_hd__mux2_1 _2279_ (.A0(\tms1x00.RAM[52][0] ),
    .A1(\tms1x00.RAM[53][0] ),
    .S(_0755_),
    .X(_0797_));
 sky130_fd_sc_hd__or2b_1 _2280_ (.A(_0694_),
    .B_N(_0797_),
    .X(_0798_));
 sky130_fd_sc_hd__mux4_1 _2281_ (.A0(\tms1x00.RAM[48][0] ),
    .A1(\tms1x00.RAM[49][0] ),
    .A2(\tms1x00.RAM[50][0] ),
    .A3(\tms1x00.RAM[51][0] ),
    .S0(_0750_),
    .S1(_0702_),
    .X(_0799_));
 sky130_fd_sc_hd__o21ai_1 _2282_ (.A1(_0726_),
    .A2(_0799_),
    .B1(_0697_),
    .Y(_0800_));
 sky130_fd_sc_hd__a31o_1 _2283_ (.A1(_0678_),
    .A2(_0796_),
    .A3(_0798_),
    .B1(_0800_),
    .X(_0801_));
 sky130_fd_sc_hd__mux4_1 _2284_ (.A0(\tms1x00.RAM[60][0] ),
    .A1(\tms1x00.RAM[61][0] ),
    .A2(\tms1x00.RAM[62][0] ),
    .A3(\tms1x00.RAM[63][0] ),
    .S0(_0724_),
    .S1(_0703_),
    .X(_0802_));
 sky130_fd_sc_hd__mux4_1 _2285_ (.A0(\tms1x00.RAM[56][0] ),
    .A1(\tms1x00.RAM[57][0] ),
    .A2(\tms1x00.RAM[58][0] ),
    .A3(\tms1x00.RAM[59][0] ),
    .S0(_0704_),
    .S1(_0707_),
    .X(_0803_));
 sky130_fd_sc_hd__o21a_1 _2286_ (.A1(_0675_),
    .A2(_0803_),
    .B1(_0682_),
    .X(_0804_));
 sky130_fd_sc_hd__o21ai_1 _2287_ (.A1(_0740_),
    .A2(_0802_),
    .B1(_0804_),
    .Y(_0805_));
 sky130_fd_sc_hd__mux4_1 _2288_ (.A0(\tms1x00.RAM[44][0] ),
    .A1(\tms1x00.RAM[45][0] ),
    .A2(\tms1x00.RAM[46][0] ),
    .A3(\tms1x00.RAM[47][0] ),
    .S0(_0755_),
    .S1(_0702_),
    .X(_0806_));
 sky130_fd_sc_hd__nor2_1 _2289_ (.A(_0721_),
    .B(_0806_),
    .Y(_0807_));
 sky130_fd_sc_hd__mux4_1 _2290_ (.A0(\tms1x00.RAM[40][0] ),
    .A1(\tms1x00.RAM[41][0] ),
    .A2(\tms1x00.RAM[42][0] ),
    .A3(\tms1x00.RAM[43][0] ),
    .S0(_0685_),
    .S1(_0736_),
    .X(_0808_));
 sky130_fd_sc_hd__o21ai_1 _2291_ (.A1(_0677_),
    .A2(_0808_),
    .B1(_0746_),
    .Y(_0809_));
 sky130_fd_sc_hd__mux4_1 _2292_ (.A0(\tms1x00.RAM[32][0] ),
    .A1(\tms1x00.RAM[33][0] ),
    .A2(\tms1x00.RAM[34][0] ),
    .A3(\tms1x00.RAM[35][0] ),
    .S0(_0755_),
    .S1(_0744_),
    .X(_0810_));
 sky130_fd_sc_hd__nor2_1 _2293_ (.A(_0742_),
    .B(_0810_),
    .Y(_0811_));
 sky130_fd_sc_hd__mux4_1 _2294_ (.A0(\tms1x00.RAM[36][0] ),
    .A1(\tms1x00.RAM[37][0] ),
    .A2(\tms1x00.RAM[38][0] ),
    .A3(\tms1x00.RAM[39][0] ),
    .S0(_0685_),
    .S1(_0736_),
    .X(_0812_));
 sky130_fd_sc_hd__o21ai_1 _2295_ (.A1(_0758_),
    .A2(_0812_),
    .B1(_0728_),
    .Y(_0813_));
 sky130_fd_sc_hd__o221a_1 _2296_ (.A1(_0807_),
    .A2(_0809_),
    .B1(_0811_),
    .B2(_0813_),
    .C1(_0761_),
    .X(_0814_));
 sky130_fd_sc_hd__a311o_1 _2297_ (.A1(_0699_),
    .A2(_0801_),
    .A3(_0805_),
    .B1(_0814_),
    .C1(_0749_),
    .X(_0815_));
 sky130_fd_sc_hd__inv_2 _2298_ (.A(_0007_),
    .Y(_0816_));
 sky130_fd_sc_hd__o211a_1 _2299_ (.A1(_0780_),
    .A2(_0794_),
    .B1(_0815_),
    .C1(_0816_),
    .X(_0817_));
 sky130_fd_sc_hd__o22ai_1 _2300_ (.A1(\tms1x00.ins_in[7] ),
    .A2(_0643_),
    .B1(_0764_),
    .B2(_0817_),
    .Y(_0818_));
 sky130_fd_sc_hd__nor2_1 _2301_ (.A(\tms1x00.ins_in[1] ),
    .B(\tms1x00.ins_in[0] ),
    .Y(_0819_));
 sky130_fd_sc_hd__and3_1 _2302_ (.A(\tms1x00.ins_in[3] ),
    .B(\tms1x00.ins_in[2] ),
    .C(_0819_),
    .X(_0820_));
 sky130_fd_sc_hd__or4b_1 _2303_ (.A(\tms1x00.ins_in[4] ),
    .B(net16),
    .C(_0647_),
    .D_N(_0820_),
    .X(_0821_));
 sky130_fd_sc_hd__nor2_1 _2304_ (.A(\tms1x00.ins_in[5] ),
    .B(_0821_),
    .Y(_0822_));
 sky130_fd_sc_hd__or3_1 _2305_ (.A(\tms1x00.ins_in[7] ),
    .B(\tms1x00.ins_in[6] ),
    .C(_0822_),
    .X(_0823_));
 sky130_fd_sc_hd__nor3_2 _2306_ (.A(\tms1x00.ins_in[1] ),
    .B(\tms1x00.ins_in[0] ),
    .C(_0662_),
    .Y(_0824_));
 sky130_fd_sc_hd__a32o_1 _2307_ (.A1(_0662_),
    .A2(_0818_),
    .A3(_0823_),
    .B1(_0824_),
    .B2(\tms1x00.A[0] ),
    .X(_0825_));
 sky130_fd_sc_hd__buf_4 _2308_ (.A(_0825_),
    .X(_0826_));
 sky130_fd_sc_hd__clkbuf_4 _2309_ (.A(_0826_),
    .X(_0827_));
 sky130_fd_sc_hd__nand3b_1 _2310_ (.A_N(\tms1x00.ram_addr_buff[4] ),
    .B(\tms1x00.ram_addr_buff[5] ),
    .C(\tms1x00.ram_addr_buff[6] ),
    .Y(_0828_));
 sky130_fd_sc_hd__buf_4 _2311_ (.A(_0828_),
    .X(_0829_));
 sky130_fd_sc_hd__and2_1 _2312_ (.A(_0821_),
    .B(_0662_),
    .X(_0830_));
 sky130_fd_sc_hd__or3_1 _2313_ (.A(\tms1x00.ram_addr_buff[2] ),
    .B(\tms1x00.ram_addr_buff[3] ),
    .C(_0830_),
    .X(_0831_));
 sky130_fd_sc_hd__nand2_1 _2314_ (.A(\tms1x00.ram_addr_buff[0] ),
    .B(\tms1x00.ram_addr_buff[1] ),
    .Y(_0832_));
 sky130_fd_sc_hd__or2_4 _2315_ (.A(_0831_),
    .B(_0832_),
    .X(_0833_));
 sky130_fd_sc_hd__or2_2 _2316_ (.A(_0829_),
    .B(_0833_),
    .X(_0834_));
 sky130_fd_sc_hd__mux2_1 _2317_ (.A0(_0827_),
    .A1(\tms1x00.RAM[99][0] ),
    .S(_0834_),
    .X(_0835_));
 sky130_fd_sc_hd__clkbuf_1 _2318_ (.A(_0835_),
    .X(_0016_));
 sky130_fd_sc_hd__mux2_1 _2319_ (.A0(\tms1x00.RAM[92][1] ),
    .A1(\tms1x00.RAM[93][1] ),
    .S(_0671_),
    .X(_0836_));
 sky130_fd_sc_hd__inv_2 _2320_ (.A(_0836_),
    .Y(_0837_));
 sky130_fd_sc_hd__mux2_1 _2321_ (.A0(\tms1x00.RAM[94][1] ),
    .A1(\tms1x00.RAM[95][1] ),
    .S(_0709_),
    .X(_0838_));
 sky130_fd_sc_hd__nand2_1 _2322_ (.A(_0670_),
    .B(_0838_),
    .Y(_0839_));
 sky130_fd_sc_hd__o211a_1 _2323_ (.A1(_0666_),
    .A2(_0837_),
    .B1(_0839_),
    .C1(_0675_),
    .X(_0840_));
 sky130_fd_sc_hd__mux4_1 _2324_ (.A0(\tms1x00.RAM[88][1] ),
    .A1(\tms1x00.RAM[89][1] ),
    .A2(\tms1x00.RAM[90][1] ),
    .A3(\tms1x00.RAM[91][1] ),
    .S0(_0679_),
    .S1(_0665_),
    .X(_0841_));
 sky130_fd_sc_hd__o21ai_1 _2325_ (.A1(_0678_),
    .A2(_0841_),
    .B1(_0682_),
    .Y(_0842_));
 sky130_fd_sc_hd__mux4_1 _2326_ (.A0(\tms1x00.RAM[80][1] ),
    .A1(\tms1x00.RAM[81][1] ),
    .A2(\tms1x00.RAM[82][1] ),
    .A3(\tms1x00.RAM[83][1] ),
    .S0(_0686_),
    .S1(_0781_),
    .X(_0843_));
 sky130_fd_sc_hd__nor2_1 _2327_ (.A(_0684_),
    .B(_0843_),
    .Y(_0844_));
 sky130_fd_sc_hd__mux4_1 _2328_ (.A0(\tms1x00.RAM[84][1] ),
    .A1(\tms1x00.RAM[85][1] ),
    .A2(\tms1x00.RAM[86][1] ),
    .A3(\tms1x00.RAM[87][1] ),
    .S0(_0693_),
    .S1(_0680_),
    .X(_0845_));
 sky130_fd_sc_hd__o21ai_1 _2329_ (.A1(_0692_),
    .A2(_0845_),
    .B1(_0697_),
    .Y(_0846_));
 sky130_fd_sc_hd__o221a_1 _2330_ (.A1(_0840_),
    .A2(_0842_),
    .B1(_0844_),
    .B2(_0846_),
    .C1(_0005_),
    .X(_0847_));
 sky130_fd_sc_hd__mux2_1 _2331_ (.A0(\tms1x00.RAM[76][1] ),
    .A1(\tms1x00.RAM[77][1] ),
    .S(_0782_),
    .X(_0848_));
 sky130_fd_sc_hd__and2b_1 _2332_ (.A_N(_0703_),
    .B(_0848_),
    .X(_0849_));
 sky130_fd_sc_hd__mux2_1 _2333_ (.A0(\tms1x00.RAM[78][1] ),
    .A1(\tms1x00.RAM[79][1] ),
    .S(_0709_),
    .X(_0850_));
 sky130_fd_sc_hd__a21o_1 _2334_ (.A1(_0708_),
    .A2(_0850_),
    .B1(_0711_),
    .X(_0851_));
 sky130_fd_sc_hd__mux4_2 _2335_ (.A0(\tms1x00.RAM[72][1] ),
    .A1(\tms1x00.RAM[73][1] ),
    .A2(\tms1x00.RAM[74][1] ),
    .A3(\tms1x00.RAM[75][1] ),
    .S0(_0693_),
    .S1(_0694_),
    .X(_0852_));
 sky130_fd_sc_hd__o221a_1 _2336_ (.A1(_0849_),
    .A2(_0851_),
    .B1(_0852_),
    .B2(_0714_),
    .C1(_0715_),
    .X(_0853_));
 sky130_fd_sc_hd__mux2_1 _2337_ (.A0(\tms1x00.RAM[68][1] ),
    .A1(\tms1x00.RAM[69][1] ),
    .S(_0709_),
    .X(_0854_));
 sky130_fd_sc_hd__and2b_1 _2338_ (.A_N(_0773_),
    .B(_0854_),
    .X(_0855_));
 sky130_fd_sc_hd__mux2_1 _2339_ (.A0(\tms1x00.RAM[70][1] ),
    .A1(\tms1x00.RAM[71][1] ),
    .S(_0719_),
    .X(_0856_));
 sky130_fd_sc_hd__a21o_1 _2340_ (.A1(_0670_),
    .A2(_0856_),
    .B1(_0758_),
    .X(_0857_));
 sky130_fd_sc_hd__mux4_2 _2341_ (.A0(\tms1x00.RAM[64][1] ),
    .A1(\tms1x00.RAM[65][1] ),
    .A2(\tms1x00.RAM[66][1] ),
    .A3(\tms1x00.RAM[67][1] ),
    .S0(_0686_),
    .S1(_0781_),
    .X(_0858_));
 sky130_fd_sc_hd__o221a_1 _2342_ (.A1(_0855_),
    .A2(_0857_),
    .B1(_0858_),
    .B2(_0684_),
    .C1(_0729_),
    .X(_0859_));
 sky130_fd_sc_hd__nor3_1 _2343_ (.A(_0701_),
    .B(_0853_),
    .C(_0859_),
    .Y(_0860_));
 sky130_fd_sc_hd__mux2_1 _2344_ (.A0(\tms1x00.RAM[118][1] ),
    .A1(\tms1x00.RAM[119][1] ),
    .S(_0679_),
    .X(_0861_));
 sky130_fd_sc_hd__nand2_1 _2345_ (.A(_0666_),
    .B(_0861_),
    .Y(_0862_));
 sky130_fd_sc_hd__mux2_1 _2346_ (.A0(\tms1x00.RAM[116][1] ),
    .A1(\tms1x00.RAM[117][1] ),
    .S(_0750_),
    .X(_0863_));
 sky130_fd_sc_hd__or2b_1 _2347_ (.A(_0680_),
    .B_N(_0863_),
    .X(_0864_));
 sky130_fd_sc_hd__mux4_1 _2348_ (.A0(\tms1x00.RAM[112][1] ),
    .A1(\tms1x00.RAM[113][1] ),
    .A2(\tms1x00.RAM[114][1] ),
    .A3(\tms1x00.RAM[115][1] ),
    .S0(_0723_),
    .S1(_0687_),
    .X(_0865_));
 sky130_fd_sc_hd__o21ai_1 _2349_ (.A1(_0726_),
    .A2(_0865_),
    .B1(_0728_),
    .Y(_0866_));
 sky130_fd_sc_hd__a31o_1 _2350_ (.A1(_0678_),
    .A2(_0862_),
    .A3(_0864_),
    .B1(_0866_),
    .X(_0867_));
 sky130_fd_sc_hd__mux4_1 _2351_ (.A0(\tms1x00.RAM[124][1] ),
    .A1(\tms1x00.RAM[125][1] ),
    .A2(\tms1x00.RAM[126][1] ),
    .A3(\tms1x00.RAM[127][1] ),
    .S0(_0724_),
    .S1(_0703_),
    .X(_0868_));
 sky130_fd_sc_hd__mux4_1 _2352_ (.A0(\tms1x00.RAM[120][1] ),
    .A1(\tms1x00.RAM[121][1] ),
    .A2(\tms1x00.RAM[122][1] ),
    .A3(\tms1x00.RAM[123][1] ),
    .S0(_0782_),
    .S1(_0707_),
    .X(_0869_));
 sky130_fd_sc_hd__o21a_1 _2353_ (.A1(_0675_),
    .A2(_0869_),
    .B1(_0746_),
    .X(_0870_));
 sky130_fd_sc_hd__o21ai_1 _2354_ (.A1(_0740_),
    .A2(_0868_),
    .B1(_0870_),
    .Y(_0871_));
 sky130_fd_sc_hd__mux4_1 _2355_ (.A0(\tms1x00.RAM[108][1] ),
    .A1(\tms1x00.RAM[109][1] ),
    .A2(\tms1x00.RAM[110][1] ),
    .A3(\tms1x00.RAM[111][1] ),
    .S0(_0750_),
    .S1(_0687_),
    .X(_0872_));
 sky130_fd_sc_hd__nor2_1 _2356_ (.A(_0721_),
    .B(_0872_),
    .Y(_0873_));
 sky130_fd_sc_hd__mux4_1 _2357_ (.A0(\tms1x00.RAM[104][1] ),
    .A1(\tms1x00.RAM[105][1] ),
    .A2(\tms1x00.RAM[106][1] ),
    .A3(\tms1x00.RAM[107][1] ),
    .S0(_0667_),
    .S1(_0664_),
    .X(_0874_));
 sky130_fd_sc_hd__o21ai_1 _2358_ (.A1(_0677_),
    .A2(_0874_),
    .B1(_0746_),
    .Y(_0875_));
 sky130_fd_sc_hd__mux4_1 _2359_ (.A0(\tms1x00.RAM[96][1] ),
    .A1(\tms1x00.RAM[97][1] ),
    .A2(\tms1x00.RAM[98][1] ),
    .A3(\tms1x00.RAM[99][1] ),
    .S0(_0755_),
    .S1(_0702_),
    .X(_0876_));
 sky130_fd_sc_hd__nor2_1 _2360_ (.A(_0726_),
    .B(_0876_),
    .Y(_0877_));
 sky130_fd_sc_hd__mux4_2 _2361_ (.A0(\tms1x00.RAM[100][1] ),
    .A1(\tms1x00.RAM[101][1] ),
    .A2(\tms1x00.RAM[102][1] ),
    .A3(\tms1x00.RAM[103][1] ),
    .S0(_0685_),
    .S1(_0736_),
    .X(_0878_));
 sky130_fd_sc_hd__o21ai_2 _2362_ (.A1(_0711_),
    .A2(_0878_),
    .B1(_0696_),
    .Y(_0879_));
 sky130_fd_sc_hd__o221a_1 _2363_ (.A1(_0873_),
    .A2(_0875_),
    .B1(_0877_),
    .B2(_0879_),
    .C1(_0761_),
    .X(_0880_));
 sky130_fd_sc_hd__a311o_1 _2364_ (.A1(_0699_),
    .A2(_0867_),
    .A3(_0871_),
    .B1(_0880_),
    .C1(_0749_),
    .X(_0881_));
 sky130_fd_sc_hd__o311a_2 _2365_ (.A1(_0663_),
    .A2(_0847_),
    .A3(_0860_),
    .B1(_0007_),
    .C1(_0881_),
    .X(_0882_));
 sky130_fd_sc_hd__mux2_1 _2366_ (.A0(\tms1x00.RAM[6][1] ),
    .A1(\tms1x00.RAM[7][1] ),
    .S(_0766_),
    .X(_0883_));
 sky130_fd_sc_hd__mux2_1 _2367_ (.A0(\tms1x00.RAM[4][1] ),
    .A1(\tms1x00.RAM[5][1] ),
    .S(_0782_),
    .X(_0884_));
 sky130_fd_sc_hd__and2b_1 _2368_ (.A_N(_0703_),
    .B(_0884_),
    .X(_0885_));
 sky130_fd_sc_hd__a211o_1 _2369_ (.A1(_0765_),
    .A2(_0883_),
    .B1(_0885_),
    .C1(_0740_),
    .X(_0886_));
 sky130_fd_sc_hd__mux4_1 _2370_ (.A0(\tms1x00.RAM[0][1] ),
    .A1(\tms1x00.RAM[1][1] ),
    .A2(\tms1x00.RAM[2][1] ),
    .A3(\tms1x00.RAM[3][1] ),
    .S0(_0693_),
    .S1(_0680_),
    .X(_0887_));
 sky130_fd_sc_hd__or2_1 _2371_ (.A(_0714_),
    .B(_0887_),
    .X(_0888_));
 sky130_fd_sc_hd__mux2_1 _2372_ (.A0(\tms1x00.RAM[12][1] ),
    .A1(\tms1x00.RAM[13][1] ),
    .S(_0704_),
    .X(_0889_));
 sky130_fd_sc_hd__and2b_1 _2373_ (.A_N(_0773_),
    .B(_0889_),
    .X(_0890_));
 sky130_fd_sc_hd__mux2_1 _2374_ (.A0(\tms1x00.RAM[14][1] ),
    .A1(\tms1x00.RAM[15][1] ),
    .S(_0719_),
    .X(_0891_));
 sky130_fd_sc_hd__a21o_1 _2375_ (.A1(_0670_),
    .A2(_0891_),
    .B1(_0758_),
    .X(_0892_));
 sky130_fd_sc_hd__mux4_1 _2376_ (.A0(\tms1x00.RAM[8][1] ),
    .A1(\tms1x00.RAM[9][1] ),
    .A2(\tms1x00.RAM[10][1] ),
    .A3(\tms1x00.RAM[11][1] ),
    .S0(_0686_),
    .S1(_0781_),
    .X(_0893_));
 sky130_fd_sc_hd__o221a_1 _2377_ (.A1(_0890_),
    .A2(_0892_),
    .B1(_0893_),
    .B2(_0684_),
    .C1(_0715_),
    .X(_0894_));
 sky130_fd_sc_hd__a311oi_1 _2378_ (.A1(_0729_),
    .A2(_0886_),
    .A3(_0888_),
    .B1(_0701_),
    .C1(_0894_),
    .Y(_0895_));
 sky130_fd_sc_hd__mux2_1 _2379_ (.A0(\tms1x00.RAM[28][1] ),
    .A1(\tms1x00.RAM[29][1] ),
    .S(_0743_),
    .X(_0896_));
 sky130_fd_sc_hd__or2b_1 _2380_ (.A(_0781_),
    .B_N(_0896_),
    .X(_0897_));
 sky130_fd_sc_hd__mux2_1 _2381_ (.A0(\tms1x00.RAM[30][1] ),
    .A1(\tms1x00.RAM[31][1] ),
    .S(_0679_),
    .X(_0898_));
 sky130_fd_sc_hd__nand2_1 _2382_ (.A(_0765_),
    .B(_0898_),
    .Y(_0899_));
 sky130_fd_sc_hd__mux4_1 _2383_ (.A0(\tms1x00.RAM[24][1] ),
    .A1(\tms1x00.RAM[25][1] ),
    .A2(\tms1x00.RAM[26][1] ),
    .A3(\tms1x00.RAM[27][1] ),
    .S0(_0743_),
    .S1(_0744_),
    .X(_0900_));
 sky130_fd_sc_hd__o21ai_1 _2384_ (.A1(_0742_),
    .A2(_0900_),
    .B1(_0682_),
    .Y(_0901_));
 sky130_fd_sc_hd__a31o_1 _2385_ (.A1(_0714_),
    .A2(_0897_),
    .A3(_0899_),
    .B1(_0901_),
    .X(_0902_));
 sky130_fd_sc_hd__mux4_1 _2386_ (.A0(\tms1x00.RAM[16][1] ),
    .A1(\tms1x00.RAM[17][1] ),
    .A2(\tms1x00.RAM[18][1] ),
    .A3(\tms1x00.RAM[19][1] ),
    .S0(_0766_),
    .S1(_0773_),
    .X(_0903_));
 sky130_fd_sc_hd__mux4_1 _2387_ (.A0(\tms1x00.RAM[20][1] ),
    .A1(\tms1x00.RAM[21][1] ),
    .A2(\tms1x00.RAM[22][1] ),
    .A3(\tms1x00.RAM[23][1] ),
    .S0(_0709_),
    .S1(_0707_),
    .X(_0904_));
 sky130_fd_sc_hd__o21a_1 _2388_ (.A1(_0692_),
    .A2(_0904_),
    .B1(_0697_),
    .X(_0905_));
 sky130_fd_sc_hd__o21ai_1 _2389_ (.A1(_0727_),
    .A2(_0903_),
    .B1(_0905_),
    .Y(_0906_));
 sky130_fd_sc_hd__a31o_1 _2390_ (.A1(_0699_),
    .A2(_0902_),
    .A3(_0906_),
    .B1(_0663_),
    .X(_0907_));
 sky130_fd_sc_hd__mux2_1 _2391_ (.A0(\tms1x00.RAM[54][1] ),
    .A1(\tms1x00.RAM[55][1] ),
    .S(_0679_),
    .X(_0908_));
 sky130_fd_sc_hd__nand2_1 _2392_ (.A(_0666_),
    .B(_0908_),
    .Y(_0909_));
 sky130_fd_sc_hd__mux2_1 _2393_ (.A0(\tms1x00.RAM[52][1] ),
    .A1(\tms1x00.RAM[53][1] ),
    .S(_0750_),
    .X(_0910_));
 sky130_fd_sc_hd__or2b_1 _2394_ (.A(_0694_),
    .B_N(_0910_),
    .X(_0911_));
 sky130_fd_sc_hd__mux4_1 _2395_ (.A0(\tms1x00.RAM[48][1] ),
    .A1(\tms1x00.RAM[49][1] ),
    .A2(\tms1x00.RAM[50][1] ),
    .A3(\tms1x00.RAM[51][1] ),
    .S0(_0723_),
    .S1(_0687_),
    .X(_0912_));
 sky130_fd_sc_hd__o21ai_1 _2396_ (.A1(_0726_),
    .A2(_0912_),
    .B1(_0697_),
    .Y(_0913_));
 sky130_fd_sc_hd__a31o_1 _2397_ (.A1(_0678_),
    .A2(_0909_),
    .A3(_0911_),
    .B1(_0913_),
    .X(_0914_));
 sky130_fd_sc_hd__mux4_1 _2398_ (.A0(\tms1x00.RAM[60][1] ),
    .A1(\tms1x00.RAM[61][1] ),
    .A2(\tms1x00.RAM[62][1] ),
    .A3(\tms1x00.RAM[63][1] ),
    .S0(_0724_),
    .S1(_0703_),
    .X(_0915_));
 sky130_fd_sc_hd__mux4_1 _2399_ (.A0(\tms1x00.RAM[56][1] ),
    .A1(\tms1x00.RAM[57][1] ),
    .A2(\tms1x00.RAM[58][1] ),
    .A3(\tms1x00.RAM[59][1] ),
    .S0(_0782_),
    .S1(_0707_),
    .X(_0916_));
 sky130_fd_sc_hd__o21a_1 _2400_ (.A1(_0675_),
    .A2(_0916_),
    .B1(_0682_),
    .X(_0917_));
 sky130_fd_sc_hd__o21ai_1 _2401_ (.A1(_0740_),
    .A2(_0915_),
    .B1(_0917_),
    .Y(_0918_));
 sky130_fd_sc_hd__mux4_1 _2402_ (.A0(\tms1x00.RAM[44][1] ),
    .A1(\tms1x00.RAM[45][1] ),
    .A2(\tms1x00.RAM[46][1] ),
    .A3(\tms1x00.RAM[47][1] ),
    .S0(_0750_),
    .S1(_0702_),
    .X(_0919_));
 sky130_fd_sc_hd__nor2_1 _2403_ (.A(_0721_),
    .B(_0919_),
    .Y(_0920_));
 sky130_fd_sc_hd__mux4_1 _2404_ (.A0(\tms1x00.RAM[40][1] ),
    .A1(\tms1x00.RAM[41][1] ),
    .A2(\tms1x00.RAM[42][1] ),
    .A3(\tms1x00.RAM[43][1] ),
    .S0(_0667_),
    .S1(_0664_),
    .X(_0921_));
 sky130_fd_sc_hd__o21ai_1 _2405_ (.A1(_0677_),
    .A2(_0921_),
    .B1(_0746_),
    .Y(_0922_));
 sky130_fd_sc_hd__mux4_1 _2406_ (.A0(\tms1x00.RAM[32][1] ),
    .A1(\tms1x00.RAM[33][1] ),
    .A2(\tms1x00.RAM[34][1] ),
    .A3(\tms1x00.RAM[35][1] ),
    .S0(_0755_),
    .S1(_0702_),
    .X(_0923_));
 sky130_fd_sc_hd__nor2_1 _2407_ (.A(_0742_),
    .B(_0923_),
    .Y(_0924_));
 sky130_fd_sc_hd__mux4_1 _2408_ (.A0(\tms1x00.RAM[36][1] ),
    .A1(\tms1x00.RAM[37][1] ),
    .A2(\tms1x00.RAM[38][1] ),
    .A3(\tms1x00.RAM[39][1] ),
    .S0(_0685_),
    .S1(_0736_),
    .X(_0925_));
 sky130_fd_sc_hd__o21ai_1 _2409_ (.A1(_0711_),
    .A2(_0925_),
    .B1(_0696_),
    .Y(_0926_));
 sky130_fd_sc_hd__o221a_1 _2410_ (.A1(_0920_),
    .A2(_0922_),
    .B1(_0924_),
    .B2(_0926_),
    .C1(_0761_),
    .X(_0927_));
 sky130_fd_sc_hd__a311o_1 _2411_ (.A1(_0699_),
    .A2(_0914_),
    .A3(_0918_),
    .B1(_0927_),
    .C1(_0749_),
    .X(_0928_));
 sky130_fd_sc_hd__o211a_1 _2412_ (.A1(_0895_),
    .A2(_0907_),
    .B1(_0928_),
    .C1(_0816_),
    .X(_0929_));
 sky130_fd_sc_hd__and2b_1 _2413_ (.A_N(\tms1x00.ins_in[7] ),
    .B(\tms1x00.ins_in[6] ),
    .X(_0930_));
 sky130_fd_sc_hd__o21bai_1 _2414_ (.A1(_0882_),
    .A2(_0929_),
    .B1_N(_0930_),
    .Y(_0931_));
 sky130_fd_sc_hd__o21ai_1 _2415_ (.A1(\tms1x00.ins_in[5] ),
    .A2(_0821_),
    .B1(_0930_),
    .Y(_0932_));
 sky130_fd_sc_hd__a32o_1 _2416_ (.A1(_0662_),
    .A2(_0931_),
    .A3(_0932_),
    .B1(_0824_),
    .B2(\tms1x00.A[1] ),
    .X(_0933_));
 sky130_fd_sc_hd__buf_4 _2417_ (.A(_0933_),
    .X(_0934_));
 sky130_fd_sc_hd__clkbuf_4 _2418_ (.A(_0934_),
    .X(_0935_));
 sky130_fd_sc_hd__mux2_1 _2419_ (.A0(_0935_),
    .A1(\tms1x00.RAM[99][1] ),
    .S(_0834_),
    .X(_0936_));
 sky130_fd_sc_hd__clkbuf_1 _2420_ (.A(_0936_),
    .X(_0017_));
 sky130_fd_sc_hd__mux2_1 _2421_ (.A0(\tms1x00.RAM[92][2] ),
    .A1(\tms1x00.RAM[93][2] ),
    .S(_0667_),
    .X(_0937_));
 sky130_fd_sc_hd__inv_2 _2422_ (.A(_0937_),
    .Y(_0938_));
 sky130_fd_sc_hd__mux2_1 _2423_ (.A0(\tms1x00.RAM[94][2] ),
    .A1(\tms1x00.RAM[95][2] ),
    .S(_0672_),
    .X(_0939_));
 sky130_fd_sc_hd__nand2_1 _2424_ (.A(_0670_),
    .B(_0939_),
    .Y(_0940_));
 sky130_fd_sc_hd__o211a_1 _2425_ (.A1(_0666_),
    .A2(_0938_),
    .B1(_0940_),
    .C1(_0675_),
    .X(_0941_));
 sky130_fd_sc_hd__mux4_2 _2426_ (.A0(\tms1x00.RAM[88][2] ),
    .A1(\tms1x00.RAM[89][2] ),
    .A2(\tms1x00.RAM[90][2] ),
    .A3(\tms1x00.RAM[91][2] ),
    .S0(_0679_),
    .S1(_0680_),
    .X(_0942_));
 sky130_fd_sc_hd__o21ai_1 _2427_ (.A1(_0678_),
    .A2(_0942_),
    .B1(_0682_),
    .Y(_0943_));
 sky130_fd_sc_hd__mux4_1 _2428_ (.A0(\tms1x00.RAM[80][2] ),
    .A1(\tms1x00.RAM[81][2] ),
    .A2(\tms1x00.RAM[82][2] ),
    .A3(\tms1x00.RAM[83][2] ),
    .S0(_0686_),
    .S1(_0781_),
    .X(_0944_));
 sky130_fd_sc_hd__nor2_1 _2429_ (.A(_0684_),
    .B(_0944_),
    .Y(_0945_));
 sky130_fd_sc_hd__mux4_1 _2430_ (.A0(\tms1x00.RAM[84][2] ),
    .A1(\tms1x00.RAM[85][2] ),
    .A2(\tms1x00.RAM[86][2] ),
    .A3(\tms1x00.RAM[87][2] ),
    .S0(_0693_),
    .S1(_0694_),
    .X(_0946_));
 sky130_fd_sc_hd__o21ai_1 _2431_ (.A1(_0692_),
    .A2(_0946_),
    .B1(_0697_),
    .Y(_0947_));
 sky130_fd_sc_hd__o221a_1 _2432_ (.A1(_0941_),
    .A2(_0943_),
    .B1(_0945_),
    .B2(_0947_),
    .C1(_0699_),
    .X(_0948_));
 sky130_fd_sc_hd__mux2_1 _2433_ (.A0(\tms1x00.RAM[76][2] ),
    .A1(\tms1x00.RAM[77][2] ),
    .S(_0782_),
    .X(_0949_));
 sky130_fd_sc_hd__and2b_1 _2434_ (.A_N(_0703_),
    .B(_0949_),
    .X(_0950_));
 sky130_fd_sc_hd__mux2_1 _2435_ (.A0(\tms1x00.RAM[78][2] ),
    .A1(\tms1x00.RAM[79][2] ),
    .S(_0709_),
    .X(_0951_));
 sky130_fd_sc_hd__a21o_1 _2436_ (.A1(_0708_),
    .A2(_0951_),
    .B1(_0711_),
    .X(_0952_));
 sky130_fd_sc_hd__mux4_1 _2437_ (.A0(\tms1x00.RAM[72][2] ),
    .A1(\tms1x00.RAM[73][2] ),
    .A2(\tms1x00.RAM[74][2] ),
    .A3(\tms1x00.RAM[75][2] ),
    .S0(_0693_),
    .S1(_0694_),
    .X(_0953_));
 sky130_fd_sc_hd__o221a_1 _2438_ (.A1(_0950_),
    .A2(_0952_),
    .B1(_0953_),
    .B2(_0714_),
    .C1(_0715_),
    .X(_0954_));
 sky130_fd_sc_hd__mux2_1 _2439_ (.A0(\tms1x00.RAM[68][2] ),
    .A1(\tms1x00.RAM[69][2] ),
    .S(_0672_),
    .X(_0955_));
 sky130_fd_sc_hd__and2b_1 _2440_ (.A_N(_0708_),
    .B(_0955_),
    .X(_0956_));
 sky130_fd_sc_hd__mux2_1 _2441_ (.A0(\tms1x00.RAM[70][2] ),
    .A1(\tms1x00.RAM[71][2] ),
    .S(_0719_),
    .X(_0957_));
 sky130_fd_sc_hd__a21o_1 _2442_ (.A1(_0670_),
    .A2(_0957_),
    .B1(_0721_),
    .X(_0958_));
 sky130_fd_sc_hd__mux4_2 _2443_ (.A0(\tms1x00.RAM[64][2] ),
    .A1(\tms1x00.RAM[65][2] ),
    .A2(\tms1x00.RAM[66][2] ),
    .A3(\tms1x00.RAM[67][2] ),
    .S0(_0724_),
    .S1(_0688_),
    .X(_0959_));
 sky130_fd_sc_hd__o221a_1 _2444_ (.A1(_0956_),
    .A2(_0958_),
    .B1(_0959_),
    .B2(_0727_),
    .C1(_0729_),
    .X(_0960_));
 sky130_fd_sc_hd__nor3_1 _2445_ (.A(_0701_),
    .B(_0954_),
    .C(_0960_),
    .Y(_0961_));
 sky130_fd_sc_hd__mux2_1 _2446_ (.A0(\tms1x00.RAM[118][2] ),
    .A1(\tms1x00.RAM[119][2] ),
    .S(_0719_),
    .X(_0962_));
 sky130_fd_sc_hd__nand2_1 _2447_ (.A(_0666_),
    .B(_0962_),
    .Y(_0963_));
 sky130_fd_sc_hd__mux2_1 _2448_ (.A0(\tms1x00.RAM[116][2] ),
    .A1(\tms1x00.RAM[117][2] ),
    .S(_0723_),
    .X(_0964_));
 sky130_fd_sc_hd__or2b_1 _2449_ (.A(_0680_),
    .B_N(_0964_),
    .X(_0965_));
 sky130_fd_sc_hd__mux4_1 _2450_ (.A0(\tms1x00.RAM[112][2] ),
    .A1(\tms1x00.RAM[113][2] ),
    .A2(\tms1x00.RAM[114][2] ),
    .A3(\tms1x00.RAM[115][2] ),
    .S0(_0685_),
    .S1(_0736_),
    .X(_0966_));
 sky130_fd_sc_hd__o21ai_1 _2451_ (.A1(_0726_),
    .A2(_0966_),
    .B1(_0728_),
    .Y(_0967_));
 sky130_fd_sc_hd__a31o_1 _2452_ (.A1(_0678_),
    .A2(_0963_),
    .A3(_0965_),
    .B1(_0967_),
    .X(_0968_));
 sky130_fd_sc_hd__mux4_1 _2453_ (.A0(\tms1x00.RAM[124][2] ),
    .A1(\tms1x00.RAM[125][2] ),
    .A2(\tms1x00.RAM[126][2] ),
    .A3(\tms1x00.RAM[127][2] ),
    .S0(_0724_),
    .S1(_0688_),
    .X(_0969_));
 sky130_fd_sc_hd__mux4_1 _2454_ (.A0(\tms1x00.RAM[120][2] ),
    .A1(\tms1x00.RAM[121][2] ),
    .A2(\tms1x00.RAM[122][2] ),
    .A3(\tms1x00.RAM[123][2] ),
    .S0(_0743_),
    .S1(_0744_),
    .X(_0970_));
 sky130_fd_sc_hd__o21a_1 _2455_ (.A1(_0742_),
    .A2(_0970_),
    .B1(_0746_),
    .X(_0971_));
 sky130_fd_sc_hd__o21ai_1 _2456_ (.A1(_0740_),
    .A2(_0969_),
    .B1(_0971_),
    .Y(_0972_));
 sky130_fd_sc_hd__mux4_2 _2457_ (.A0(\tms1x00.RAM[108][2] ),
    .A1(\tms1x00.RAM[109][2] ),
    .A2(\tms1x00.RAM[110][2] ),
    .A3(\tms1x00.RAM[111][2] ),
    .S0(_0750_),
    .S1(_0702_),
    .X(_0973_));
 sky130_fd_sc_hd__nor2_1 _2458_ (.A(_0721_),
    .B(_0973_),
    .Y(_0974_));
 sky130_fd_sc_hd__mux4_1 _2459_ (.A0(\tms1x00.RAM[104][2] ),
    .A1(\tms1x00.RAM[105][2] ),
    .A2(\tms1x00.RAM[106][2] ),
    .A3(\tms1x00.RAM[107][2] ),
    .S0(_0667_),
    .S1(_0664_),
    .X(_0975_));
 sky130_fd_sc_hd__o21ai_1 _2460_ (.A1(_0677_),
    .A2(_0975_),
    .B1(_0746_),
    .Y(_0976_));
 sky130_fd_sc_hd__mux4_1 _2461_ (.A0(\tms1x00.RAM[96][2] ),
    .A1(\tms1x00.RAM[97][2] ),
    .A2(\tms1x00.RAM[98][2] ),
    .A3(\tms1x00.RAM[99][2] ),
    .S0(_0755_),
    .S1(_0744_),
    .X(_0977_));
 sky130_fd_sc_hd__nor2_1 _2462_ (.A(_0742_),
    .B(_0977_),
    .Y(_0978_));
 sky130_fd_sc_hd__mux4_2 _2463_ (.A0(\tms1x00.RAM[100][2] ),
    .A1(\tms1x00.RAM[101][2] ),
    .A2(\tms1x00.RAM[102][2] ),
    .A3(\tms1x00.RAM[103][2] ),
    .S0(_0685_),
    .S1(_0736_),
    .X(_0979_));
 sky130_fd_sc_hd__o21ai_1 _2464_ (.A1(_0758_),
    .A2(_0979_),
    .B1(_0728_),
    .Y(_0980_));
 sky130_fd_sc_hd__o221a_1 _2465_ (.A1(_0974_),
    .A2(_0976_),
    .B1(_0978_),
    .B2(_0980_),
    .C1(_0761_),
    .X(_0981_));
 sky130_fd_sc_hd__a311o_1 _2466_ (.A1(_0699_),
    .A2(_0968_),
    .A3(_0972_),
    .B1(_0749_),
    .C1(_0981_),
    .X(_0982_));
 sky130_fd_sc_hd__o311a_2 _2467_ (.A1(_0663_),
    .A2(_0948_),
    .A3(_0961_),
    .B1(_0982_),
    .C1(_0007_),
    .X(_0983_));
 sky130_fd_sc_hd__mux2_1 _2468_ (.A0(\tms1x00.RAM[6][2] ),
    .A1(\tms1x00.RAM[7][2] ),
    .S(_0766_),
    .X(_0984_));
 sky130_fd_sc_hd__mux2_1 _2469_ (.A0(\tms1x00.RAM[4][2] ),
    .A1(\tms1x00.RAM[5][2] ),
    .S(_0782_),
    .X(_0985_));
 sky130_fd_sc_hd__and2b_1 _2470_ (.A_N(_0703_),
    .B(_0985_),
    .X(_0986_));
 sky130_fd_sc_hd__a211o_1 _2471_ (.A1(_0765_),
    .A2(_0984_),
    .B1(_0986_),
    .C1(_0692_),
    .X(_0987_));
 sky130_fd_sc_hd__mux4_1 _2472_ (.A0(\tms1x00.RAM[0][2] ),
    .A1(\tms1x00.RAM[1][2] ),
    .A2(\tms1x00.RAM[2][2] ),
    .A3(\tms1x00.RAM[3][2] ),
    .S0(_0693_),
    .S1(_0680_),
    .X(_0988_));
 sky130_fd_sc_hd__or2_1 _2473_ (.A(_0714_),
    .B(_0988_),
    .X(_0989_));
 sky130_fd_sc_hd__mux2_1 _2474_ (.A0(\tms1x00.RAM[12][2] ),
    .A1(\tms1x00.RAM[13][2] ),
    .S(_0704_),
    .X(_0990_));
 sky130_fd_sc_hd__and2b_1 _2475_ (.A_N(_0773_),
    .B(_0990_),
    .X(_0991_));
 sky130_fd_sc_hd__mux2_1 _2476_ (.A0(\tms1x00.RAM[14][2] ),
    .A1(\tms1x00.RAM[15][2] ),
    .S(_0672_),
    .X(_0992_));
 sky130_fd_sc_hd__a21o_1 _2477_ (.A1(_0670_),
    .A2(_0992_),
    .B1(_0758_),
    .X(_0993_));
 sky130_fd_sc_hd__mux4_1 _2478_ (.A0(\tms1x00.RAM[8][2] ),
    .A1(\tms1x00.RAM[9][2] ),
    .A2(\tms1x00.RAM[10][2] ),
    .A3(\tms1x00.RAM[11][2] ),
    .S0(_0686_),
    .S1(_0781_),
    .X(_0994_));
 sky130_fd_sc_hd__o221a_1 _2479_ (.A1(_0991_),
    .A2(_0993_),
    .B1(_0994_),
    .B2(_0684_),
    .C1(_0715_),
    .X(_0995_));
 sky130_fd_sc_hd__a311oi_1 _2480_ (.A1(_0729_),
    .A2(_0987_),
    .A3(_0989_),
    .B1(_0701_),
    .C1(_0995_),
    .Y(_0996_));
 sky130_fd_sc_hd__mux2_1 _2481_ (.A0(\tms1x00.RAM[28][2] ),
    .A1(\tms1x00.RAM[29][2] ),
    .S(_0743_),
    .X(_0997_));
 sky130_fd_sc_hd__or2b_1 _2482_ (.A(_0781_),
    .B_N(_0997_),
    .X(_0998_));
 sky130_fd_sc_hd__mux2_1 _2483_ (.A0(\tms1x00.RAM[30][2] ),
    .A1(\tms1x00.RAM[31][2] ),
    .S(_0679_),
    .X(_0999_));
 sky130_fd_sc_hd__nand2_1 _2484_ (.A(_0765_),
    .B(_0999_),
    .Y(_1000_));
 sky130_fd_sc_hd__mux4_1 _2485_ (.A0(\tms1x00.RAM[24][2] ),
    .A1(\tms1x00.RAM[25][2] ),
    .A2(\tms1x00.RAM[26][2] ),
    .A3(\tms1x00.RAM[27][2] ),
    .S0(_0743_),
    .S1(_0744_),
    .X(_1001_));
 sky130_fd_sc_hd__o21ai_1 _2486_ (.A1(_0742_),
    .A2(_1001_),
    .B1(_0682_),
    .Y(_1002_));
 sky130_fd_sc_hd__a31o_1 _2487_ (.A1(_0714_),
    .A2(_0998_),
    .A3(_1000_),
    .B1(_1002_),
    .X(_1003_));
 sky130_fd_sc_hd__mux4_1 _2488_ (.A0(\tms1x00.RAM[16][2] ),
    .A1(\tms1x00.RAM[17][2] ),
    .A2(\tms1x00.RAM[18][2] ),
    .A3(\tms1x00.RAM[19][2] ),
    .S0(_0766_),
    .S1(_0773_),
    .X(_1004_));
 sky130_fd_sc_hd__mux4_1 _2489_ (.A0(\tms1x00.RAM[20][2] ),
    .A1(\tms1x00.RAM[21][2] ),
    .A2(\tms1x00.RAM[22][2] ),
    .A3(\tms1x00.RAM[23][2] ),
    .S0(_0704_),
    .S1(_0707_),
    .X(_1005_));
 sky130_fd_sc_hd__o21a_1 _2490_ (.A1(_0692_),
    .A2(_1005_),
    .B1(_0697_),
    .X(_1006_));
 sky130_fd_sc_hd__o21ai_1 _2491_ (.A1(_0727_),
    .A2(_1004_),
    .B1(_1006_),
    .Y(_1007_));
 sky130_fd_sc_hd__a31o_1 _2492_ (.A1(_0699_),
    .A2(_1003_),
    .A3(_1007_),
    .B1(_0663_),
    .X(_1008_));
 sky130_fd_sc_hd__mux2_1 _2493_ (.A0(\tms1x00.RAM[54][2] ),
    .A1(\tms1x00.RAM[55][2] ),
    .S(_0719_),
    .X(_1009_));
 sky130_fd_sc_hd__nand2_1 _2494_ (.A(_0666_),
    .B(_1009_),
    .Y(_1010_));
 sky130_fd_sc_hd__mux2_1 _2495_ (.A0(\tms1x00.RAM[52][2] ),
    .A1(\tms1x00.RAM[53][2] ),
    .S(_0750_),
    .X(_1011_));
 sky130_fd_sc_hd__or2b_1 _2496_ (.A(_0680_),
    .B_N(_1011_),
    .X(_1012_));
 sky130_fd_sc_hd__mux4_1 _2497_ (.A0(\tms1x00.RAM[48][2] ),
    .A1(\tms1x00.RAM[49][2] ),
    .A2(\tms1x00.RAM[50][2] ),
    .A3(\tms1x00.RAM[51][2] ),
    .S0(_0723_),
    .S1(_0687_),
    .X(_1013_));
 sky130_fd_sc_hd__o21ai_1 _2498_ (.A1(_0726_),
    .A2(_1013_),
    .B1(_0728_),
    .Y(_1014_));
 sky130_fd_sc_hd__a31o_1 _2499_ (.A1(_0678_),
    .A2(_1010_),
    .A3(_1012_),
    .B1(_1014_),
    .X(_1015_));
 sky130_fd_sc_hd__mux4_1 _2500_ (.A0(\tms1x00.RAM[60][2] ),
    .A1(\tms1x00.RAM[61][2] ),
    .A2(\tms1x00.RAM[62][2] ),
    .A3(\tms1x00.RAM[63][2] ),
    .S0(_0724_),
    .S1(_0688_),
    .X(_1016_));
 sky130_fd_sc_hd__mux4_1 _2501_ (.A0(\tms1x00.RAM[56][2] ),
    .A1(\tms1x00.RAM[57][2] ),
    .A2(\tms1x00.RAM[58][2] ),
    .A3(\tms1x00.RAM[59][2] ),
    .S0(_0743_),
    .S1(_0707_),
    .X(_1017_));
 sky130_fd_sc_hd__o21a_1 _2502_ (.A1(_0675_),
    .A2(_1017_),
    .B1(_0746_),
    .X(_1018_));
 sky130_fd_sc_hd__o21ai_1 _2503_ (.A1(_0740_),
    .A2(_1016_),
    .B1(_1018_),
    .Y(_1019_));
 sky130_fd_sc_hd__mux4_1 _2504_ (.A0(\tms1x00.RAM[44][2] ),
    .A1(\tms1x00.RAM[45][2] ),
    .A2(\tms1x00.RAM[46][2] ),
    .A3(\tms1x00.RAM[47][2] ),
    .S0(_0750_),
    .S1(_0687_),
    .X(_1020_));
 sky130_fd_sc_hd__nor2_1 _2505_ (.A(_0721_),
    .B(_1020_),
    .Y(_1021_));
 sky130_fd_sc_hd__mux4_1 _2506_ (.A0(\tms1x00.RAM[40][2] ),
    .A1(\tms1x00.RAM[41][2] ),
    .A2(\tms1x00.RAM[42][2] ),
    .A3(\tms1x00.RAM[43][2] ),
    .S0(_0667_),
    .S1(_0664_),
    .X(_1022_));
 sky130_fd_sc_hd__o21ai_1 _2507_ (.A1(_0677_),
    .A2(_1022_),
    .B1(_0004_),
    .Y(_1023_));
 sky130_fd_sc_hd__mux4_2 _2508_ (.A0(\tms1x00.RAM[32][2] ),
    .A1(\tms1x00.RAM[33][2] ),
    .A2(\tms1x00.RAM[34][2] ),
    .A3(\tms1x00.RAM[35][2] ),
    .S0(_0755_),
    .S1(_0702_),
    .X(_1024_));
 sky130_fd_sc_hd__nor2_1 _2509_ (.A(_0726_),
    .B(_1024_),
    .Y(_1025_));
 sky130_fd_sc_hd__mux4_1 _2510_ (.A0(\tms1x00.RAM[36][2] ),
    .A1(\tms1x00.RAM[37][2] ),
    .A2(\tms1x00.RAM[38][2] ),
    .A3(\tms1x00.RAM[39][2] ),
    .S0(_0685_),
    .S1(_0736_),
    .X(_1026_));
 sky130_fd_sc_hd__o21ai_1 _2511_ (.A1(_0711_),
    .A2(_1026_),
    .B1(_0696_),
    .Y(_1027_));
 sky130_fd_sc_hd__o221a_1 _2512_ (.A1(_1021_),
    .A2(_1023_),
    .B1(_1025_),
    .B2(_1027_),
    .C1(_0761_),
    .X(_1028_));
 sky130_fd_sc_hd__a311o_1 _2513_ (.A1(_0699_),
    .A2(_1015_),
    .A3(_1019_),
    .B1(_1028_),
    .C1(_0749_),
    .X(_1029_));
 sky130_fd_sc_hd__o211a_1 _2514_ (.A1(_0996_),
    .A2(_1008_),
    .B1(_1029_),
    .C1(_0816_),
    .X(_1030_));
 sky130_fd_sc_hd__o21ai_1 _2515_ (.A1(_0983_),
    .A2(_1030_),
    .B1(_0653_),
    .Y(_1031_));
 sky130_fd_sc_hd__or3b_1 _2516_ (.A(_0643_),
    .B(_0822_),
    .C_N(\tms1x00.ins_in[7] ),
    .X(_1032_));
 sky130_fd_sc_hd__a32o_1 _2517_ (.A1(_0662_),
    .A2(_1031_),
    .A3(_1032_),
    .B1(_0824_),
    .B2(\tms1x00.A[2] ),
    .X(_1033_));
 sky130_fd_sc_hd__buf_4 _2518_ (.A(_1033_),
    .X(_1034_));
 sky130_fd_sc_hd__clkbuf_4 _2519_ (.A(_1034_),
    .X(_1035_));
 sky130_fd_sc_hd__mux2_1 _2520_ (.A0(_1035_),
    .A1(\tms1x00.RAM[99][2] ),
    .S(_0834_),
    .X(_1036_));
 sky130_fd_sc_hd__clkbuf_1 _2521_ (.A(_1036_),
    .X(_0018_));
 sky130_fd_sc_hd__mux2_1 _2522_ (.A0(\tms1x00.RAM[116][3] ),
    .A1(\tms1x00.RAM[117][3] ),
    .S(_0671_),
    .X(_1037_));
 sky130_fd_sc_hd__and2b_1 _2523_ (.A_N(_0665_),
    .B(_1037_),
    .X(_1038_));
 sky130_fd_sc_hd__mux2_1 _2524_ (.A0(\tms1x00.RAM[118][3] ),
    .A1(\tms1x00.RAM[119][3] ),
    .S(_0667_),
    .X(_1039_));
 sky130_fd_sc_hd__a21o_1 _2525_ (.A1(_0665_),
    .A2(_1039_),
    .B1(_0691_),
    .X(_1040_));
 sky130_fd_sc_hd__mux4_1 _2526_ (.A0(\tms1x00.RAM[112][3] ),
    .A1(\tms1x00.RAM[113][3] ),
    .A2(\tms1x00.RAM[114][3] ),
    .A3(\tms1x00.RAM[115][3] ),
    .S0(_0782_),
    .S1(_0707_),
    .X(_1041_));
 sky130_fd_sc_hd__o221a_1 _2527_ (.A1(_1038_),
    .A2(_1040_),
    .B1(_1041_),
    .B2(_0675_),
    .C1(_0697_),
    .X(_1042_));
 sky130_fd_sc_hd__mux4_1 _2528_ (.A0(\tms1x00.RAM[120][3] ),
    .A1(\tms1x00.RAM[121][3] ),
    .A2(\tms1x00.RAM[122][3] ),
    .A3(\tms1x00.RAM[123][3] ),
    .S0(_0709_),
    .S1(_0665_),
    .X(_1043_));
 sky130_fd_sc_hd__mux4_1 _2529_ (.A0(\tms1x00.RAM[124][3] ),
    .A1(\tms1x00.RAM[125][3] ),
    .A2(\tms1x00.RAM[126][3] ),
    .A3(\tms1x00.RAM[127][3] ),
    .S0(_0671_),
    .S1(_0002_),
    .X(_1044_));
 sky130_fd_sc_hd__or2_1 _2530_ (.A(_0691_),
    .B(_1044_),
    .X(_1045_));
 sky130_fd_sc_hd__o211a_1 _2531_ (.A1(_0675_),
    .A2(_1043_),
    .B1(_1045_),
    .C1(_0682_),
    .X(_1046_));
 sky130_fd_sc_hd__o31a_1 _2532_ (.A1(_0761_),
    .A2(_1042_),
    .A3(_1046_),
    .B1(_0663_),
    .X(_1047_));
 sky130_fd_sc_hd__mux4_2 _2533_ (.A0(\tms1x00.RAM[100][3] ),
    .A1(\tms1x00.RAM[101][3] ),
    .A2(\tms1x00.RAM[102][3] ),
    .A3(\tms1x00.RAM[103][3] ),
    .S0(_0782_),
    .S1(_0707_),
    .X(_1048_));
 sky130_fd_sc_hd__or2_1 _2534_ (.A(_0692_),
    .B(_1048_),
    .X(_1049_));
 sky130_fd_sc_hd__mux4_1 _2535_ (.A0(\tms1x00.RAM[96][3] ),
    .A1(\tms1x00.RAM[97][3] ),
    .A2(\tms1x00.RAM[98][3] ),
    .A3(\tms1x00.RAM[99][3] ),
    .S0(_0782_),
    .S1(_0707_),
    .X(_1050_));
 sky130_fd_sc_hd__or2_1 _2536_ (.A(_0675_),
    .B(_1050_),
    .X(_1051_));
 sky130_fd_sc_hd__mux4_2 _2537_ (.A0(\tms1x00.RAM[108][3] ),
    .A1(\tms1x00.RAM[109][3] ),
    .A2(\tms1x00.RAM[110][3] ),
    .A3(\tms1x00.RAM[111][3] ),
    .S0(_0672_),
    .S1(_0665_),
    .X(_1052_));
 sky130_fd_sc_hd__mux4_1 _2538_ (.A0(\tms1x00.RAM[104][3] ),
    .A1(\tms1x00.RAM[105][3] ),
    .A2(\tms1x00.RAM[106][3] ),
    .A3(\tms1x00.RAM[107][3] ),
    .S0(_0671_),
    .S1(_0664_),
    .X(_1053_));
 sky130_fd_sc_hd__or2_1 _2539_ (.A(_0003_),
    .B(_1053_),
    .X(_1054_));
 sky130_fd_sc_hd__o211a_1 _2540_ (.A1(_0692_),
    .A2(_1052_),
    .B1(_1054_),
    .C1(_0682_),
    .X(_1055_));
 sky130_fd_sc_hd__a311o_1 _2541_ (.A1(_0729_),
    .A2(_1049_),
    .A3(_1051_),
    .B1(_0005_),
    .C1(_1055_),
    .X(_1056_));
 sky130_fd_sc_hd__mux2_1 _2542_ (.A0(\tms1x00.RAM[92][3] ),
    .A1(\tms1x00.RAM[93][3] ),
    .S(_0667_),
    .X(_1057_));
 sky130_fd_sc_hd__or2b_1 _2543_ (.A(_0665_),
    .B_N(_1057_),
    .X(_1058_));
 sky130_fd_sc_hd__mux2_1 _2544_ (.A0(\tms1x00.RAM[94][3] ),
    .A1(\tms1x00.RAM[95][3] ),
    .S(_0719_),
    .X(_1059_));
 sky130_fd_sc_hd__nand2_1 _2545_ (.A(_0666_),
    .B(_1059_),
    .Y(_1060_));
 sky130_fd_sc_hd__mux4_2 _2546_ (.A0(\tms1x00.RAM[88][3] ),
    .A1(\tms1x00.RAM[89][3] ),
    .A2(\tms1x00.RAM[90][3] ),
    .A3(\tms1x00.RAM[91][3] ),
    .S0(_0667_),
    .S1(_0664_),
    .X(_1061_));
 sky130_fd_sc_hd__o21ai_1 _2547_ (.A1(_0677_),
    .A2(_1061_),
    .B1(_0004_),
    .Y(_1062_));
 sky130_fd_sc_hd__a31o_1 _2548_ (.A1(_0678_),
    .A2(_1058_),
    .A3(_1060_),
    .B1(_1062_),
    .X(_1063_));
 sky130_fd_sc_hd__mux4_1 _2549_ (.A0(\tms1x00.RAM[80][3] ),
    .A1(\tms1x00.RAM[81][3] ),
    .A2(\tms1x00.RAM[82][3] ),
    .A3(\tms1x00.RAM[83][3] ),
    .S0(_0686_),
    .S1(_0694_),
    .X(_1064_));
 sky130_fd_sc_hd__mux4_1 _2550_ (.A0(\tms1x00.RAM[84][3] ),
    .A1(\tms1x00.RAM[85][3] ),
    .A2(\tms1x00.RAM[86][3] ),
    .A3(\tms1x00.RAM[87][3] ),
    .S0(_0723_),
    .S1(_0687_),
    .X(_1065_));
 sky130_fd_sc_hd__o21a_1 _2551_ (.A1(_0721_),
    .A2(_1065_),
    .B1(_0728_),
    .X(_1066_));
 sky130_fd_sc_hd__o21ai_1 _2552_ (.A1(_0684_),
    .A2(_1064_),
    .B1(_1066_),
    .Y(_1067_));
 sky130_fd_sc_hd__a31o_1 _2553_ (.A1(_0005_),
    .A2(_1063_),
    .A3(_1067_),
    .B1(_0663_),
    .X(_1068_));
 sky130_fd_sc_hd__mux2_1 _2554_ (.A0(\tms1x00.RAM[76][3] ),
    .A1(\tms1x00.RAM[77][3] ),
    .S(_0743_),
    .X(_1069_));
 sky130_fd_sc_hd__and2b_1 _2555_ (.A_N(_0688_),
    .B(_1069_),
    .X(_1070_));
 sky130_fd_sc_hd__mux2_1 _2556_ (.A0(\tms1x00.RAM[78][3] ),
    .A1(\tms1x00.RAM[79][3] ),
    .S(_0704_),
    .X(_1071_));
 sky130_fd_sc_hd__a21o_1 _2557_ (.A1(_0773_),
    .A2(_1071_),
    .B1(_0711_),
    .X(_1072_));
 sky130_fd_sc_hd__mux4_2 _2558_ (.A0(\tms1x00.RAM[72][3] ),
    .A1(\tms1x00.RAM[73][3] ),
    .A2(\tms1x00.RAM[74][3] ),
    .A3(\tms1x00.RAM[75][3] ),
    .S0(_0679_),
    .S1(_0680_),
    .X(_1073_));
 sky130_fd_sc_hd__o221a_1 _2559_ (.A1(_1070_),
    .A2(_1072_),
    .B1(_1073_),
    .B2(_0714_),
    .C1(_0715_),
    .X(_1074_));
 sky130_fd_sc_hd__mux2_1 _2560_ (.A0(\tms1x00.RAM[68][3] ),
    .A1(\tms1x00.RAM[69][3] ),
    .S(_0704_),
    .X(_1075_));
 sky130_fd_sc_hd__and2b_1 _2561_ (.A_N(_0773_),
    .B(_1075_),
    .X(_1076_));
 sky130_fd_sc_hd__mux2_1 _2562_ (.A0(\tms1x00.RAM[70][3] ),
    .A1(\tms1x00.RAM[71][3] ),
    .S(_0672_),
    .X(_1077_));
 sky130_fd_sc_hd__a21o_1 _2563_ (.A1(_0708_),
    .A2(_1077_),
    .B1(_0711_),
    .X(_1078_));
 sky130_fd_sc_hd__mux4_2 _2564_ (.A0(\tms1x00.RAM[64][3] ),
    .A1(\tms1x00.RAM[65][3] ),
    .A2(\tms1x00.RAM[66][3] ),
    .A3(\tms1x00.RAM[67][3] ),
    .S0(_0686_),
    .S1(_0781_),
    .X(_1079_));
 sky130_fd_sc_hd__o221a_1 _2565_ (.A1(_1076_),
    .A2(_1078_),
    .B1(_1079_),
    .B2(_0684_),
    .C1(_0729_),
    .X(_1080_));
 sky130_fd_sc_hd__nor3_1 _2566_ (.A(_0701_),
    .B(_1074_),
    .C(_1080_),
    .Y(_1081_));
 sky130_fd_sc_hd__o2bb2a_1 _2567_ (.A1_N(_1047_),
    .A2_N(_1056_),
    .B1(_1068_),
    .B2(_1081_),
    .X(_1082_));
 sky130_fd_sc_hd__mux4_1 _2568_ (.A0(\tms1x00.RAM[24][3] ),
    .A1(\tms1x00.RAM[25][3] ),
    .A2(\tms1x00.RAM[26][3] ),
    .A3(\tms1x00.RAM[27][3] ),
    .S0(_0766_),
    .S1(_0765_),
    .X(_1083_));
 sky130_fd_sc_hd__mux2_1 _2569_ (.A0(\tms1x00.RAM[30][3] ),
    .A1(\tms1x00.RAM[31][3] ),
    .S(_0766_),
    .X(_1084_));
 sky130_fd_sc_hd__mux2_1 _2570_ (.A0(\tms1x00.RAM[28][3] ),
    .A1(\tms1x00.RAM[29][3] ),
    .S(_0709_),
    .X(_1085_));
 sky130_fd_sc_hd__and2b_1 _2571_ (.A_N(_0773_),
    .B(_1085_),
    .X(_1086_));
 sky130_fd_sc_hd__a211o_1 _2572_ (.A1(_0765_),
    .A2(_1084_),
    .B1(_1086_),
    .C1(_0740_),
    .X(_1087_));
 sky130_fd_sc_hd__o211ai_1 _2573_ (.A1(_0727_),
    .A2(_1083_),
    .B1(_1087_),
    .C1(_0715_),
    .Y(_1088_));
 sky130_fd_sc_hd__mux4_1 _2574_ (.A0(\tms1x00.RAM[16][3] ),
    .A1(\tms1x00.RAM[17][3] ),
    .A2(\tms1x00.RAM[18][3] ),
    .A3(\tms1x00.RAM[19][3] ),
    .S0(_0766_),
    .S1(_0765_),
    .X(_1089_));
 sky130_fd_sc_hd__mux4_1 _2575_ (.A0(\tms1x00.RAM[20][3] ),
    .A1(\tms1x00.RAM[21][3] ),
    .A2(\tms1x00.RAM[22][3] ),
    .A3(\tms1x00.RAM[23][3] ),
    .S0(_0766_),
    .S1(_0708_),
    .X(_1090_));
 sky130_fd_sc_hd__o21a_1 _2576_ (.A1(_0740_),
    .A2(_1090_),
    .B1(_0729_),
    .X(_1091_));
 sky130_fd_sc_hd__o21ai_1 _2577_ (.A1(_0727_),
    .A2(_1089_),
    .B1(_1091_),
    .Y(_1092_));
 sky130_fd_sc_hd__mux2_1 _2578_ (.A0(\tms1x00.RAM[12][3] ),
    .A1(\tms1x00.RAM[13][3] ),
    .S(_0704_),
    .X(_1093_));
 sky130_fd_sc_hd__and2b_1 _2579_ (.A_N(_0773_),
    .B(_1093_),
    .X(_1094_));
 sky130_fd_sc_hd__mux2_1 _2580_ (.A0(\tms1x00.RAM[14][3] ),
    .A1(\tms1x00.RAM[15][3] ),
    .S(_0672_),
    .X(_1095_));
 sky130_fd_sc_hd__a21o_1 _2581_ (.A1(_0670_),
    .A2(_1095_),
    .B1(_0758_),
    .X(_1096_));
 sky130_fd_sc_hd__mux4_1 _2582_ (.A0(\tms1x00.RAM[8][3] ),
    .A1(\tms1x00.RAM[9][3] ),
    .A2(\tms1x00.RAM[10][3] ),
    .A3(\tms1x00.RAM[11][3] ),
    .S0(_0686_),
    .S1(_0781_),
    .X(_1097_));
 sky130_fd_sc_hd__o221a_1 _2583_ (.A1(_1094_),
    .A2(_1096_),
    .B1(_1097_),
    .B2(_0684_),
    .C1(_0715_),
    .X(_1098_));
 sky130_fd_sc_hd__mux2_1 _2584_ (.A0(\tms1x00.RAM[4][3] ),
    .A1(\tms1x00.RAM[5][3] ),
    .S(_0672_),
    .X(_1099_));
 sky130_fd_sc_hd__and2b_1 _2585_ (.A_N(_0708_),
    .B(_1099_),
    .X(_1100_));
 sky130_fd_sc_hd__mux2_1 _2586_ (.A0(\tms1x00.RAM[6][3] ),
    .A1(\tms1x00.RAM[7][3] ),
    .S(_0719_),
    .X(_1101_));
 sky130_fd_sc_hd__a21o_1 _2587_ (.A1(_0666_),
    .A2(_1101_),
    .B1(_0721_),
    .X(_1102_));
 sky130_fd_sc_hd__mux4_1 _2588_ (.A0(\tms1x00.RAM[0][3] ),
    .A1(\tms1x00.RAM[1][3] ),
    .A2(\tms1x00.RAM[2][3] ),
    .A3(\tms1x00.RAM[3][3] ),
    .S0(_0724_),
    .S1(_0688_),
    .X(_1103_));
 sky130_fd_sc_hd__o221a_1 _2589_ (.A1(_1100_),
    .A2(_1102_),
    .B1(_1103_),
    .B2(_0727_),
    .C1(_0729_),
    .X(_1104_));
 sky130_fd_sc_hd__nor3_1 _2590_ (.A(_0701_),
    .B(_1098_),
    .C(_1104_),
    .Y(_1105_));
 sky130_fd_sc_hd__a311o_1 _2591_ (.A1(_0701_),
    .A2(_1088_),
    .A3(_1092_),
    .B1(_1105_),
    .C1(_0663_),
    .X(_1106_));
 sky130_fd_sc_hd__mux2_1 _2592_ (.A0(\tms1x00.RAM[52][3] ),
    .A1(\tms1x00.RAM[53][3] ),
    .S(_0704_),
    .X(_1107_));
 sky130_fd_sc_hd__and2b_1 _2593_ (.A_N(_0703_),
    .B(_1107_),
    .X(_1108_));
 sky130_fd_sc_hd__mux2_1 _2594_ (.A0(\tms1x00.RAM[54][3] ),
    .A1(\tms1x00.RAM[55][3] ),
    .S(_0672_),
    .X(_1109_));
 sky130_fd_sc_hd__a21o_1 _2595_ (.A1(_0708_),
    .A2(_1109_),
    .B1(_0711_),
    .X(_1110_));
 sky130_fd_sc_hd__mux4_1 _2596_ (.A0(\tms1x00.RAM[48][3] ),
    .A1(\tms1x00.RAM[49][3] ),
    .A2(\tms1x00.RAM[50][3] ),
    .A3(\tms1x00.RAM[51][3] ),
    .S0(_0693_),
    .S1(_0694_),
    .X(_1111_));
 sky130_fd_sc_hd__o221a_1 _2597_ (.A1(_1108_),
    .A2(_1110_),
    .B1(_1111_),
    .B2(_0684_),
    .C1(_0697_),
    .X(_1112_));
 sky130_fd_sc_hd__mux4_1 _2598_ (.A0(\tms1x00.RAM[56][3] ),
    .A1(\tms1x00.RAM[57][3] ),
    .A2(\tms1x00.RAM[58][3] ),
    .A3(\tms1x00.RAM[59][3] ),
    .S0(_0724_),
    .S1(_0688_),
    .X(_1113_));
 sky130_fd_sc_hd__mux4_1 _2599_ (.A0(\tms1x00.RAM[60][3] ),
    .A1(\tms1x00.RAM[61][3] ),
    .A2(\tms1x00.RAM[62][3] ),
    .A3(\tms1x00.RAM[63][3] ),
    .S0(_0723_),
    .S1(_0687_),
    .X(_1114_));
 sky130_fd_sc_hd__or2_1 _2600_ (.A(_0758_),
    .B(_1114_),
    .X(_1115_));
 sky130_fd_sc_hd__o211a_1 _2601_ (.A1(_0727_),
    .A2(_1113_),
    .B1(_1115_),
    .C1(_0715_),
    .X(_1116_));
 sky130_fd_sc_hd__mux4_1 _2602_ (.A0(\tms1x00.RAM[44][3] ),
    .A1(\tms1x00.RAM[45][3] ),
    .A2(\tms1x00.RAM[46][3] ),
    .A3(\tms1x00.RAM[47][3] ),
    .S0(_0723_),
    .S1(_0687_),
    .X(_1117_));
 sky130_fd_sc_hd__or2_1 _2603_ (.A(_0758_),
    .B(_1117_),
    .X(_1118_));
 sky130_fd_sc_hd__mux4_2 _2604_ (.A0(\tms1x00.RAM[40][3] ),
    .A1(\tms1x00.RAM[41][3] ),
    .A2(\tms1x00.RAM[42][3] ),
    .A3(\tms1x00.RAM[43][3] ),
    .S0(_0755_),
    .S1(_0702_),
    .X(_1119_));
 sky130_fd_sc_hd__o21a_1 _2605_ (.A1(_0742_),
    .A2(_1119_),
    .B1(_0746_),
    .X(_1120_));
 sky130_fd_sc_hd__mux4_1 _2606_ (.A0(\tms1x00.RAM[32][3] ),
    .A1(\tms1x00.RAM[33][3] ),
    .A2(\tms1x00.RAM[34][3] ),
    .A3(\tms1x00.RAM[35][3] ),
    .S0(_0750_),
    .S1(_0687_),
    .X(_1121_));
 sky130_fd_sc_hd__or2_1 _2607_ (.A(_0726_),
    .B(_1121_),
    .X(_1122_));
 sky130_fd_sc_hd__mux4_1 _2608_ (.A0(\tms1x00.RAM[36][3] ),
    .A1(\tms1x00.RAM[37][3] ),
    .A2(\tms1x00.RAM[38][3] ),
    .A3(\tms1x00.RAM[39][3] ),
    .S0(_0755_),
    .S1(_0744_),
    .X(_1123_));
 sky130_fd_sc_hd__o21a_1 _2609_ (.A1(_0692_),
    .A2(_1123_),
    .B1(_0728_),
    .X(_1124_));
 sky130_fd_sc_hd__a221o_1 _2610_ (.A1(_1118_),
    .A2(_1120_),
    .B1(_1122_),
    .B2(_1124_),
    .C1(_0005_),
    .X(_1125_));
 sky130_fd_sc_hd__o311a_1 _2611_ (.A1(_0761_),
    .A2(_1112_),
    .A3(_1116_),
    .B1(_1125_),
    .C1(_0663_),
    .X(_1126_));
 sky130_fd_sc_hd__nor2_1 _2612_ (.A(_0007_),
    .B(_1126_),
    .Y(_1127_));
 sky130_fd_sc_hd__a22oi_4 _2613_ (.A1(_0007_),
    .A2(_1082_),
    .B1(_1106_),
    .B2(_1127_),
    .Y(_1128_));
 sky130_fd_sc_hd__nand2_1 _2614_ (.A(\tms1x00.ins_in[7] ),
    .B(\tms1x00.ins_in[6] ),
    .Y(_1129_));
 sky130_fd_sc_hd__and3_1 _2615_ (.A(\tms1x00.ins_in[7] ),
    .B(_0643_),
    .C(_0822_),
    .X(_1130_));
 sky130_fd_sc_hd__a221o_1 _2616_ (.A1(\tms1x00.A[3] ),
    .A2(_0824_),
    .B1(_1128_),
    .B2(_1129_),
    .C1(_1130_),
    .X(_1131_));
 sky130_fd_sc_hd__clkbuf_4 _2617_ (.A(_1131_),
    .X(_1132_));
 sky130_fd_sc_hd__clkbuf_4 _2618_ (.A(_1132_),
    .X(_1133_));
 sky130_fd_sc_hd__mux2_1 _2619_ (.A0(_1133_),
    .A1(\tms1x00.RAM[99][3] ),
    .S(_0834_),
    .X(_1134_));
 sky130_fd_sc_hd__clkbuf_1 _2620_ (.A(_1134_),
    .X(_0019_));
 sky130_fd_sc_hd__clkbuf_4 _2621_ (.A(_0826_),
    .X(_1135_));
 sky130_fd_sc_hd__nand3b_1 _2622_ (.A_N(\tms1x00.ram_addr_buff[5] ),
    .B(\tms1x00.ram_addr_buff[6] ),
    .C(\tms1x00.ram_addr_buff[4] ),
    .Y(_1136_));
 sky130_fd_sc_hd__clkbuf_8 _2623_ (.A(_1136_),
    .X(_1137_));
 sky130_fd_sc_hd__or3b_1 _2624_ (.A(\tms1x00.ram_addr_buff[2] ),
    .B(_0830_),
    .C_N(\tms1x00.ram_addr_buff[3] ),
    .X(_1138_));
 sky130_fd_sc_hd__or3b_1 _2625_ (.A(\tms1x00.ram_addr_buff[1] ),
    .B(_1138_),
    .C_N(_0620_),
    .X(_1139_));
 sky130_fd_sc_hd__clkbuf_8 _2626_ (.A(_1139_),
    .X(_1140_));
 sky130_fd_sc_hd__nor2_2 _2627_ (.A(_1137_),
    .B(_1140_),
    .Y(_1141_));
 sky130_fd_sc_hd__mux2_1 _2628_ (.A0(\tms1x00.RAM[89][0] ),
    .A1(_1135_),
    .S(_1141_),
    .X(_1142_));
 sky130_fd_sc_hd__clkbuf_1 _2629_ (.A(_1142_),
    .X(_0020_));
 sky130_fd_sc_hd__buf_2 _2630_ (.A(_0934_),
    .X(_1143_));
 sky130_fd_sc_hd__mux2_1 _2631_ (.A0(\tms1x00.RAM[89][1] ),
    .A1(_1143_),
    .S(_1141_),
    .X(_1144_));
 sky130_fd_sc_hd__clkbuf_1 _2632_ (.A(_1144_),
    .X(_0021_));
 sky130_fd_sc_hd__clkbuf_4 _2633_ (.A(_1034_),
    .X(_1145_));
 sky130_fd_sc_hd__mux2_1 _2634_ (.A0(\tms1x00.RAM[89][2] ),
    .A1(_1145_),
    .S(_1141_),
    .X(_1146_));
 sky130_fd_sc_hd__clkbuf_1 _2635_ (.A(_1146_),
    .X(_0022_));
 sky130_fd_sc_hd__clkbuf_4 _2636_ (.A(_1132_),
    .X(_1147_));
 sky130_fd_sc_hd__mux2_1 _2637_ (.A0(\tms1x00.RAM[89][3] ),
    .A1(_1147_),
    .S(_1141_),
    .X(_1148_));
 sky130_fd_sc_hd__clkbuf_1 _2638_ (.A(_1148_),
    .X(_0023_));
 sky130_fd_sc_hd__nand2_1 _2639_ (.A(\tms1x00.ram_addr_buff[4] ),
    .B(\tms1x00.ram_addr_buff[5] ),
    .Y(_1149_));
 sky130_fd_sc_hd__or2_1 _2640_ (.A(\tms1x00.ram_addr_buff[6] ),
    .B(_1149_),
    .X(_1150_));
 sky130_fd_sc_hd__buf_6 _2641_ (.A(_1150_),
    .X(_1151_));
 sky130_fd_sc_hd__or2_1 _2642_ (.A(_0832_),
    .B(_1138_),
    .X(_1152_));
 sky130_fd_sc_hd__buf_6 _2643_ (.A(_1152_),
    .X(_1153_));
 sky130_fd_sc_hd__nor2_2 _2644_ (.A(_1151_),
    .B(_1153_),
    .Y(_1154_));
 sky130_fd_sc_hd__mux2_1 _2645_ (.A0(\tms1x00.RAM[59][0] ),
    .A1(_1135_),
    .S(_1154_),
    .X(_1155_));
 sky130_fd_sc_hd__clkbuf_1 _2646_ (.A(_1155_),
    .X(_0024_));
 sky130_fd_sc_hd__mux2_1 _2647_ (.A0(\tms1x00.RAM[59][1] ),
    .A1(_1143_),
    .S(_1154_),
    .X(_1156_));
 sky130_fd_sc_hd__clkbuf_1 _2648_ (.A(_1156_),
    .X(_0025_));
 sky130_fd_sc_hd__mux2_1 _2649_ (.A0(\tms1x00.RAM[59][2] ),
    .A1(_1145_),
    .S(_1154_),
    .X(_1157_));
 sky130_fd_sc_hd__clkbuf_1 _2650_ (.A(_1157_),
    .X(_0026_));
 sky130_fd_sc_hd__mux2_1 _2651_ (.A0(\tms1x00.RAM[59][3] ),
    .A1(_1147_),
    .S(_1154_),
    .X(_1158_));
 sky130_fd_sc_hd__clkbuf_1 _2652_ (.A(_1158_),
    .X(_0027_));
 sky130_fd_sc_hd__and3b_2 _2653_ (.A_N(_0635_),
    .B(_0637_),
    .C(_0639_),
    .X(_1159_));
 sky130_fd_sc_hd__and3b_1 _2654_ (.A_N(_0830_),
    .B(\tms1x00.ram_addr_buff[3] ),
    .C(\tms1x00.ram_addr_buff[2] ),
    .X(_1160_));
 sky130_fd_sc_hd__and3b_1 _2655_ (.A_N(_0628_),
    .B(_1160_),
    .C(_0620_),
    .X(_1161_));
 sky130_fd_sc_hd__clkbuf_8 _2656_ (.A(_1161_),
    .X(_1162_));
 sky130_fd_sc_hd__nand2_2 _2657_ (.A(_1159_),
    .B(_1162_),
    .Y(_1163_));
 sky130_fd_sc_hd__mux2_1 _2658_ (.A0(_0827_),
    .A1(\tms1x00.RAM[109][0] ),
    .S(_1163_),
    .X(_1164_));
 sky130_fd_sc_hd__clkbuf_1 _2659_ (.A(_1164_),
    .X(_0028_));
 sky130_fd_sc_hd__mux2_1 _2660_ (.A0(_0935_),
    .A1(\tms1x00.RAM[109][1] ),
    .S(_1163_),
    .X(_1165_));
 sky130_fd_sc_hd__clkbuf_1 _2661_ (.A(_1165_),
    .X(_0029_));
 sky130_fd_sc_hd__mux2_1 _2662_ (.A0(_1035_),
    .A1(\tms1x00.RAM[109][2] ),
    .S(_1163_),
    .X(_1166_));
 sky130_fd_sc_hd__clkbuf_1 _2663_ (.A(_1166_),
    .X(_0030_));
 sky130_fd_sc_hd__mux2_1 _2664_ (.A0(_1133_),
    .A1(\tms1x00.RAM[109][3] ),
    .S(_1163_),
    .X(_1167_));
 sky130_fd_sc_hd__clkbuf_1 _2665_ (.A(_1167_),
    .X(_0031_));
 sky130_fd_sc_hd__nor3b_2 _2666_ (.A(_0635_),
    .B(_0637_),
    .C_N(_0639_),
    .Y(_1168_));
 sky130_fd_sc_hd__and3_1 _2667_ (.A(_0620_),
    .B(_0628_),
    .C(_1160_),
    .X(_1169_));
 sky130_fd_sc_hd__buf_4 _2668_ (.A(_1169_),
    .X(_1170_));
 sky130_fd_sc_hd__nand2_2 _2669_ (.A(_1168_),
    .B(_1170_),
    .Y(_1171_));
 sky130_fd_sc_hd__mux2_1 _2670_ (.A0(_0827_),
    .A1(\tms1x00.RAM[79][0] ),
    .S(_1171_),
    .X(_1172_));
 sky130_fd_sc_hd__clkbuf_1 _2671_ (.A(_1172_),
    .X(_0032_));
 sky130_fd_sc_hd__mux2_1 _2672_ (.A0(_0935_),
    .A1(\tms1x00.RAM[79][1] ),
    .S(_1171_),
    .X(_1173_));
 sky130_fd_sc_hd__clkbuf_1 _2673_ (.A(_1173_),
    .X(_0033_));
 sky130_fd_sc_hd__mux2_1 _2674_ (.A0(_1035_),
    .A1(\tms1x00.RAM[79][2] ),
    .S(_1171_),
    .X(_1174_));
 sky130_fd_sc_hd__clkbuf_1 _2675_ (.A(_1174_),
    .X(_0034_));
 sky130_fd_sc_hd__mux2_1 _2676_ (.A0(_1133_),
    .A1(\tms1x00.RAM[79][3] ),
    .S(_1171_),
    .X(_1175_));
 sky130_fd_sc_hd__clkbuf_1 _2677_ (.A(_1175_),
    .X(_0035_));
 sky130_fd_sc_hd__or3b_1 _2678_ (.A(\tms1x00.ram_addr_buff[4] ),
    .B(\tms1x00.ram_addr_buff[5] ),
    .C_N(\tms1x00.ram_addr_buff[6] ),
    .X(_1176_));
 sky130_fd_sc_hd__clkbuf_8 _2679_ (.A(_1176_),
    .X(_1177_));
 sky130_fd_sc_hd__or3b_1 _2680_ (.A(\tms1x00.ram_addr_buff[3] ),
    .B(_0830_),
    .C_N(\tms1x00.ram_addr_buff[2] ),
    .X(_1178_));
 sky130_fd_sc_hd__or3b_1 _2681_ (.A(\tms1x00.ram_addr_buff[1] ),
    .B(_1178_),
    .C_N(\tms1x00.ram_addr_buff[0] ),
    .X(_1179_));
 sky130_fd_sc_hd__buf_6 _2682_ (.A(_1179_),
    .X(_1180_));
 sky130_fd_sc_hd__nor2_2 _2683_ (.A(_1177_),
    .B(_1180_),
    .Y(_1181_));
 sky130_fd_sc_hd__mux2_1 _2684_ (.A0(\tms1x00.RAM[69][0] ),
    .A1(_1135_),
    .S(_1181_),
    .X(_1182_));
 sky130_fd_sc_hd__clkbuf_1 _2685_ (.A(_1182_),
    .X(_0036_));
 sky130_fd_sc_hd__mux2_1 _2686_ (.A0(\tms1x00.RAM[69][1] ),
    .A1(_1143_),
    .S(_1181_),
    .X(_1183_));
 sky130_fd_sc_hd__clkbuf_1 _2687_ (.A(_1183_),
    .X(_0037_));
 sky130_fd_sc_hd__mux2_1 _2688_ (.A0(\tms1x00.RAM[69][2] ),
    .A1(_1145_),
    .S(_1181_),
    .X(_1184_));
 sky130_fd_sc_hd__clkbuf_1 _2689_ (.A(_1184_),
    .X(_0038_));
 sky130_fd_sc_hd__mux2_1 _2690_ (.A0(\tms1x00.RAM[69][3] ),
    .A1(_1147_),
    .S(_1181_),
    .X(_1185_));
 sky130_fd_sc_hd__clkbuf_1 _2691_ (.A(_1185_),
    .X(_0039_));
 sky130_fd_sc_hd__and3_2 _2692_ (.A(_0635_),
    .B(_0637_),
    .C(_0639_),
    .X(_1186_));
 sky130_fd_sc_hd__nand2_2 _2693_ (.A(_1170_),
    .B(_1186_),
    .Y(_1187_));
 sky130_fd_sc_hd__mux2_1 _2694_ (.A0(_0827_),
    .A1(\tms1x00.RAM[127][0] ),
    .S(_1187_),
    .X(_1188_));
 sky130_fd_sc_hd__clkbuf_1 _2695_ (.A(_1188_),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_1 _2696_ (.A0(_0935_),
    .A1(\tms1x00.RAM[127][1] ),
    .S(_1187_),
    .X(_1189_));
 sky130_fd_sc_hd__clkbuf_1 _2697_ (.A(_1189_),
    .X(_0041_));
 sky130_fd_sc_hd__mux2_1 _2698_ (.A0(_1035_),
    .A1(\tms1x00.RAM[127][2] ),
    .S(_1187_),
    .X(_1190_));
 sky130_fd_sc_hd__clkbuf_1 _2699_ (.A(_1190_),
    .X(_0042_));
 sky130_fd_sc_hd__mux2_1 _2700_ (.A0(_1133_),
    .A1(\tms1x00.RAM[127][3] ),
    .S(_1187_),
    .X(_1191_));
 sky130_fd_sc_hd__clkbuf_1 _2701_ (.A(_1191_),
    .X(_0043_));
 sky130_fd_sc_hd__and2_1 _2702_ (.A(net20),
    .B(_0000_),
    .X(_1192_));
 sky130_fd_sc_hd__mux2_1 _2703_ (.A0(net56),
    .A1(net29),
    .S(_1192_),
    .X(_1193_));
 sky130_fd_sc_hd__clkbuf_1 _2704_ (.A(_1193_),
    .X(_0044_));
 sky130_fd_sc_hd__or3b_4 _2705_ (.A(_0628_),
    .B(_0831_),
    .C_N(_0620_),
    .X(_1194_));
 sky130_fd_sc_hd__or2_1 _2706_ (.A(_1151_),
    .B(_1194_),
    .X(_1195_));
 sky130_fd_sc_hd__mux2_1 _2707_ (.A0(_0827_),
    .A1(\tms1x00.RAM[49][0] ),
    .S(_1195_),
    .X(_1196_));
 sky130_fd_sc_hd__clkbuf_1 _2708_ (.A(_1196_),
    .X(_0045_));
 sky130_fd_sc_hd__mux2_1 _2709_ (.A0(_0935_),
    .A1(\tms1x00.RAM[49][1] ),
    .S(_1195_),
    .X(_1197_));
 sky130_fd_sc_hd__clkbuf_1 _2710_ (.A(_1197_),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_1 _2711_ (.A0(_1035_),
    .A1(\tms1x00.RAM[49][2] ),
    .S(_1195_),
    .X(_1198_));
 sky130_fd_sc_hd__clkbuf_1 _2712_ (.A(_1198_),
    .X(_0047_));
 sky130_fd_sc_hd__mux2_1 _2713_ (.A0(_1133_),
    .A1(\tms1x00.RAM[49][3] ),
    .S(_1195_),
    .X(_1199_));
 sky130_fd_sc_hd__clkbuf_1 _2714_ (.A(_1199_),
    .X(_0048_));
 sky130_fd_sc_hd__or3b_1 _2715_ (.A(\tms1x00.ram_addr_buff[5] ),
    .B(\tms1x00.ram_addr_buff[6] ),
    .C_N(\tms1x00.ram_addr_buff[4] ),
    .X(_1200_));
 sky130_fd_sc_hd__or2_2 _2716_ (.A(_0833_),
    .B(_1200_),
    .X(_1201_));
 sky130_fd_sc_hd__mux2_1 _2717_ (.A0(_0827_),
    .A1(\tms1x00.RAM[19][0] ),
    .S(_1201_),
    .X(_1202_));
 sky130_fd_sc_hd__clkbuf_1 _2718_ (.A(_1202_),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_1 _2719_ (.A0(_0935_),
    .A1(\tms1x00.RAM[19][1] ),
    .S(_1201_),
    .X(_1203_));
 sky130_fd_sc_hd__clkbuf_1 _2720_ (.A(_1203_),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _2721_ (.A0(_1035_),
    .A1(\tms1x00.RAM[19][2] ),
    .S(_1201_),
    .X(_1204_));
 sky130_fd_sc_hd__clkbuf_1 _2722_ (.A(_1204_),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _2723_ (.A0(_1133_),
    .A1(\tms1x00.RAM[19][3] ),
    .S(_1201_),
    .X(_1205_));
 sky130_fd_sc_hd__clkbuf_1 _2724_ (.A(_1205_),
    .X(_0052_));
 sky130_fd_sc_hd__and3b_2 _2725_ (.A_N(_0637_),
    .B(_0639_),
    .C(_0635_),
    .X(_1206_));
 sky130_fd_sc_hd__nand2_2 _2726_ (.A(_1206_),
    .B(_1170_),
    .Y(_1207_));
 sky130_fd_sc_hd__mux2_1 _2727_ (.A0(_0827_),
    .A1(\tms1x00.RAM[95][0] ),
    .S(_1207_),
    .X(_1208_));
 sky130_fd_sc_hd__clkbuf_1 _2728_ (.A(_1208_),
    .X(_0053_));
 sky130_fd_sc_hd__mux2_1 _2729_ (.A0(_0935_),
    .A1(\tms1x00.RAM[95][1] ),
    .S(_1207_),
    .X(_1209_));
 sky130_fd_sc_hd__clkbuf_1 _2730_ (.A(_1209_),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _2731_ (.A0(_1035_),
    .A1(\tms1x00.RAM[95][2] ),
    .S(_1207_),
    .X(_1210_));
 sky130_fd_sc_hd__clkbuf_1 _2732_ (.A(_1210_),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _2733_ (.A0(_1133_),
    .A1(\tms1x00.RAM[95][3] ),
    .S(_1207_),
    .X(_1211_));
 sky130_fd_sc_hd__clkbuf_1 _2734_ (.A(_1211_),
    .X(_0056_));
 sky130_fd_sc_hd__and3b_1 _2735_ (.A_N(_0620_),
    .B(_0628_),
    .C(_1160_),
    .X(_1212_));
 sky130_fd_sc_hd__buf_4 _2736_ (.A(_1212_),
    .X(_1213_));
 sky130_fd_sc_hd__nand2_2 _2737_ (.A(_1206_),
    .B(_1213_),
    .Y(_1214_));
 sky130_fd_sc_hd__mux2_1 _2738_ (.A0(_0827_),
    .A1(\tms1x00.RAM[94][0] ),
    .S(_1214_),
    .X(_1215_));
 sky130_fd_sc_hd__clkbuf_1 _2739_ (.A(_1215_),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _2740_ (.A0(_0935_),
    .A1(\tms1x00.RAM[94][1] ),
    .S(_1214_),
    .X(_1216_));
 sky130_fd_sc_hd__clkbuf_1 _2741_ (.A(_1216_),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_1 _2742_ (.A0(_1035_),
    .A1(\tms1x00.RAM[94][2] ),
    .S(_1214_),
    .X(_1217_));
 sky130_fd_sc_hd__clkbuf_1 _2743_ (.A(_1217_),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _2744_ (.A0(_1133_),
    .A1(\tms1x00.RAM[94][3] ),
    .S(_1214_),
    .X(_1218_));
 sky130_fd_sc_hd__clkbuf_1 _2745_ (.A(_1218_),
    .X(_0060_));
 sky130_fd_sc_hd__nand2_2 _2746_ (.A(_1206_),
    .B(_1162_),
    .Y(_1219_));
 sky130_fd_sc_hd__mux2_1 _2747_ (.A0(_0827_),
    .A1(\tms1x00.RAM[93][0] ),
    .S(_1219_),
    .X(_1220_));
 sky130_fd_sc_hd__clkbuf_1 _2748_ (.A(_1220_),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _2749_ (.A0(_0935_),
    .A1(\tms1x00.RAM[93][1] ),
    .S(_1219_),
    .X(_1221_));
 sky130_fd_sc_hd__clkbuf_1 _2750_ (.A(_1221_),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _2751_ (.A0(_1035_),
    .A1(\tms1x00.RAM[93][2] ),
    .S(_1219_),
    .X(_1222_));
 sky130_fd_sc_hd__clkbuf_1 _2752_ (.A(_1222_),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _2753_ (.A0(_1133_),
    .A1(\tms1x00.RAM[93][3] ),
    .S(_1219_),
    .X(_1223_));
 sky130_fd_sc_hd__clkbuf_1 _2754_ (.A(_1223_),
    .X(_0064_));
 sky130_fd_sc_hd__nor3b_4 _2755_ (.A(_0620_),
    .B(_0628_),
    .C_N(_1160_),
    .Y(_1224_));
 sky130_fd_sc_hd__nand2_2 _2756_ (.A(_1206_),
    .B(_1224_),
    .Y(_1225_));
 sky130_fd_sc_hd__mux2_1 _2757_ (.A0(_0827_),
    .A1(\tms1x00.RAM[92][0] ),
    .S(_1225_),
    .X(_1226_));
 sky130_fd_sc_hd__clkbuf_1 _2758_ (.A(_1226_),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _2759_ (.A0(_0935_),
    .A1(\tms1x00.RAM[92][1] ),
    .S(_1225_),
    .X(_1227_));
 sky130_fd_sc_hd__clkbuf_1 _2760_ (.A(_1227_),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_1 _2761_ (.A0(_1035_),
    .A1(\tms1x00.RAM[92][2] ),
    .S(_1225_),
    .X(_1228_));
 sky130_fd_sc_hd__clkbuf_1 _2762_ (.A(_1228_),
    .X(_0067_));
 sky130_fd_sc_hd__mux2_1 _2763_ (.A0(_1133_),
    .A1(\tms1x00.RAM[92][3] ),
    .S(_1225_),
    .X(_1229_));
 sky130_fd_sc_hd__clkbuf_1 _2764_ (.A(_1229_),
    .X(_0068_));
 sky130_fd_sc_hd__nor2_2 _2765_ (.A(_1137_),
    .B(_1153_),
    .Y(_1230_));
 sky130_fd_sc_hd__mux2_1 _2766_ (.A0(\tms1x00.RAM[91][0] ),
    .A1(_1135_),
    .S(_1230_),
    .X(_1231_));
 sky130_fd_sc_hd__clkbuf_1 _2767_ (.A(_1231_),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_1 _2768_ (.A0(\tms1x00.RAM[91][1] ),
    .A1(_1143_),
    .S(_1230_),
    .X(_1232_));
 sky130_fd_sc_hd__clkbuf_1 _2769_ (.A(_1232_),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _2770_ (.A0(\tms1x00.RAM[91][2] ),
    .A1(_1145_),
    .S(_1230_),
    .X(_1233_));
 sky130_fd_sc_hd__clkbuf_1 _2771_ (.A(_1233_),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _2772_ (.A0(\tms1x00.RAM[91][3] ),
    .A1(_1147_),
    .S(_1230_),
    .X(_1234_));
 sky130_fd_sc_hd__clkbuf_1 _2773_ (.A(_1234_),
    .X(_0072_));
 sky130_fd_sc_hd__or3b_1 _2774_ (.A(_1138_),
    .B(\tms1x00.ram_addr_buff[0] ),
    .C_N(_0628_),
    .X(_1235_));
 sky130_fd_sc_hd__buf_6 _2775_ (.A(_1235_),
    .X(_1236_));
 sky130_fd_sc_hd__nor2_2 _2776_ (.A(_1137_),
    .B(_1236_),
    .Y(_1237_));
 sky130_fd_sc_hd__mux2_1 _2777_ (.A0(\tms1x00.RAM[90][0] ),
    .A1(_1135_),
    .S(_1237_),
    .X(_1238_));
 sky130_fd_sc_hd__clkbuf_1 _2778_ (.A(_1238_),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _2779_ (.A0(\tms1x00.RAM[90][1] ),
    .A1(_1143_),
    .S(_1237_),
    .X(_1239_));
 sky130_fd_sc_hd__clkbuf_1 _2780_ (.A(_1239_),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _2781_ (.A0(\tms1x00.RAM[90][2] ),
    .A1(_1145_),
    .S(_1237_),
    .X(_1240_));
 sky130_fd_sc_hd__clkbuf_1 _2782_ (.A(_1240_),
    .X(_0075_));
 sky130_fd_sc_hd__mux2_1 _2783_ (.A0(\tms1x00.RAM[90][3] ),
    .A1(_1147_),
    .S(_1237_),
    .X(_1241_));
 sky130_fd_sc_hd__clkbuf_1 _2784_ (.A(_1241_),
    .X(_0076_));
 sky130_fd_sc_hd__or3_1 _2785_ (.A(\tms1x00.ram_addr_buff[4] ),
    .B(\tms1x00.ram_addr_buff[5] ),
    .C(\tms1x00.ram_addr_buff[6] ),
    .X(_1242_));
 sky130_fd_sc_hd__buf_6 _2786_ (.A(_1242_),
    .X(_1243_));
 sky130_fd_sc_hd__or3_1 _2787_ (.A(\tms1x00.ram_addr_buff[0] ),
    .B(\tms1x00.ram_addr_buff[1] ),
    .C(_1138_),
    .X(_1244_));
 sky130_fd_sc_hd__buf_6 _2788_ (.A(_1244_),
    .X(_1245_));
 sky130_fd_sc_hd__nor2_2 _2789_ (.A(_1243_),
    .B(_1245_),
    .Y(_1246_));
 sky130_fd_sc_hd__mux2_1 _2790_ (.A0(\tms1x00.RAM[8][0] ),
    .A1(_1135_),
    .S(_1246_),
    .X(_1247_));
 sky130_fd_sc_hd__clkbuf_1 _2791_ (.A(_1247_),
    .X(_0077_));
 sky130_fd_sc_hd__mux2_1 _2792_ (.A0(\tms1x00.RAM[8][1] ),
    .A1(_1143_),
    .S(_1246_),
    .X(_1248_));
 sky130_fd_sc_hd__clkbuf_1 _2793_ (.A(_1248_),
    .X(_0078_));
 sky130_fd_sc_hd__mux2_1 _2794_ (.A0(\tms1x00.RAM[8][2] ),
    .A1(_1145_),
    .S(_1246_),
    .X(_1249_));
 sky130_fd_sc_hd__clkbuf_1 _2795_ (.A(_1249_),
    .X(_0079_));
 sky130_fd_sc_hd__mux2_1 _2796_ (.A0(\tms1x00.RAM[8][3] ),
    .A1(_1147_),
    .S(_1246_),
    .X(_1250_));
 sky130_fd_sc_hd__clkbuf_1 _2797_ (.A(_1250_),
    .X(_0080_));
 sky130_fd_sc_hd__nor2_2 _2798_ (.A(_1137_),
    .B(_1245_),
    .Y(_1251_));
 sky130_fd_sc_hd__mux2_1 _2799_ (.A0(\tms1x00.RAM[88][0] ),
    .A1(_1135_),
    .S(_1251_),
    .X(_1252_));
 sky130_fd_sc_hd__clkbuf_1 _2800_ (.A(_1252_),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_1 _2801_ (.A0(\tms1x00.RAM[88][1] ),
    .A1(_1143_),
    .S(_1251_),
    .X(_1253_));
 sky130_fd_sc_hd__clkbuf_1 _2802_ (.A(_1253_),
    .X(_0082_));
 sky130_fd_sc_hd__mux2_1 _2803_ (.A0(\tms1x00.RAM[88][2] ),
    .A1(_1145_),
    .S(_1251_),
    .X(_1254_));
 sky130_fd_sc_hd__clkbuf_1 _2804_ (.A(_1254_),
    .X(_0083_));
 sky130_fd_sc_hd__mux2_1 _2805_ (.A0(\tms1x00.RAM[88][3] ),
    .A1(_1147_),
    .S(_1251_),
    .X(_1255_));
 sky130_fd_sc_hd__clkbuf_1 _2806_ (.A(_1255_),
    .X(_0084_));
 sky130_fd_sc_hd__or2_1 _2807_ (.A(_0832_),
    .B(_1178_),
    .X(_1256_));
 sky130_fd_sc_hd__buf_6 _2808_ (.A(_1256_),
    .X(_1257_));
 sky130_fd_sc_hd__nor2_2 _2809_ (.A(_1137_),
    .B(_1257_),
    .Y(_1258_));
 sky130_fd_sc_hd__mux2_1 _2810_ (.A0(\tms1x00.RAM[87][0] ),
    .A1(_1135_),
    .S(_1258_),
    .X(_1259_));
 sky130_fd_sc_hd__clkbuf_1 _2811_ (.A(_1259_),
    .X(_0085_));
 sky130_fd_sc_hd__mux2_1 _2812_ (.A0(\tms1x00.RAM[87][1] ),
    .A1(_1143_),
    .S(_1258_),
    .X(_1260_));
 sky130_fd_sc_hd__clkbuf_1 _2813_ (.A(_1260_),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_1 _2814_ (.A0(\tms1x00.RAM[87][2] ),
    .A1(_1145_),
    .S(_1258_),
    .X(_1261_));
 sky130_fd_sc_hd__clkbuf_1 _2815_ (.A(_1261_),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_1 _2816_ (.A0(\tms1x00.RAM[87][3] ),
    .A1(_1147_),
    .S(_1258_),
    .X(_1262_));
 sky130_fd_sc_hd__clkbuf_1 _2817_ (.A(_1262_),
    .X(_0088_));
 sky130_fd_sc_hd__clkbuf_4 _2818_ (.A(_0825_),
    .X(_1263_));
 sky130_fd_sc_hd__buf_2 _2819_ (.A(_1263_),
    .X(_1264_));
 sky130_fd_sc_hd__or3b_1 _2820_ (.A(_1178_),
    .B(\tms1x00.ram_addr_buff[0] ),
    .C_N(\tms1x00.ram_addr_buff[1] ),
    .X(_1265_));
 sky130_fd_sc_hd__buf_6 _2821_ (.A(_1265_),
    .X(_1266_));
 sky130_fd_sc_hd__nor2_2 _2822_ (.A(_1137_),
    .B(_1266_),
    .Y(_1267_));
 sky130_fd_sc_hd__mux2_1 _2823_ (.A0(\tms1x00.RAM[86][0] ),
    .A1(_1264_),
    .S(_1267_),
    .X(_1268_));
 sky130_fd_sc_hd__clkbuf_1 _2824_ (.A(_1268_),
    .X(_0089_));
 sky130_fd_sc_hd__clkbuf_4 _2825_ (.A(_0933_),
    .X(_1269_));
 sky130_fd_sc_hd__buf_2 _2826_ (.A(_1269_),
    .X(_1270_));
 sky130_fd_sc_hd__mux2_1 _2827_ (.A0(\tms1x00.RAM[86][1] ),
    .A1(_1270_),
    .S(_1267_),
    .X(_1271_));
 sky130_fd_sc_hd__clkbuf_1 _2828_ (.A(_1271_),
    .X(_0090_));
 sky130_fd_sc_hd__clkbuf_4 _2829_ (.A(_1033_),
    .X(_1272_));
 sky130_fd_sc_hd__buf_2 _2830_ (.A(_1272_),
    .X(_1273_));
 sky130_fd_sc_hd__mux2_1 _2831_ (.A0(\tms1x00.RAM[86][2] ),
    .A1(_1273_),
    .S(_1267_),
    .X(_1274_));
 sky130_fd_sc_hd__clkbuf_1 _2832_ (.A(_1274_),
    .X(_0091_));
 sky130_fd_sc_hd__clkbuf_4 _2833_ (.A(_1131_),
    .X(_1275_));
 sky130_fd_sc_hd__buf_2 _2834_ (.A(_1275_),
    .X(_1276_));
 sky130_fd_sc_hd__mux2_1 _2835_ (.A0(\tms1x00.RAM[86][3] ),
    .A1(_1276_),
    .S(_1267_),
    .X(_1277_));
 sky130_fd_sc_hd__clkbuf_1 _2836_ (.A(_1277_),
    .X(_0092_));
 sky130_fd_sc_hd__nor2_2 _2837_ (.A(_0829_),
    .B(_1140_),
    .Y(_1278_));
 sky130_fd_sc_hd__mux2_1 _2838_ (.A0(\tms1x00.RAM[105][0] ),
    .A1(_1264_),
    .S(_1278_),
    .X(_1279_));
 sky130_fd_sc_hd__clkbuf_1 _2839_ (.A(_1279_),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _2840_ (.A0(\tms1x00.RAM[105][1] ),
    .A1(_1270_),
    .S(_1278_),
    .X(_1280_));
 sky130_fd_sc_hd__clkbuf_1 _2841_ (.A(_1280_),
    .X(_0094_));
 sky130_fd_sc_hd__mux2_1 _2842_ (.A0(\tms1x00.RAM[105][2] ),
    .A1(_1273_),
    .S(_1278_),
    .X(_1281_));
 sky130_fd_sc_hd__clkbuf_1 _2843_ (.A(_1281_),
    .X(_0095_));
 sky130_fd_sc_hd__mux2_1 _2844_ (.A0(\tms1x00.RAM[105][3] ),
    .A1(_1276_),
    .S(_1278_),
    .X(_1282_));
 sky130_fd_sc_hd__clkbuf_1 _2845_ (.A(_1282_),
    .X(_0096_));
 sky130_fd_sc_hd__nor2_2 _2846_ (.A(_0829_),
    .B(_1245_),
    .Y(_1283_));
 sky130_fd_sc_hd__mux2_1 _2847_ (.A0(\tms1x00.RAM[104][0] ),
    .A1(_1264_),
    .S(_1283_),
    .X(_1284_));
 sky130_fd_sc_hd__clkbuf_1 _2848_ (.A(_1284_),
    .X(_0097_));
 sky130_fd_sc_hd__mux2_1 _2849_ (.A0(\tms1x00.RAM[104][1] ),
    .A1(_1270_),
    .S(_1283_),
    .X(_1285_));
 sky130_fd_sc_hd__clkbuf_1 _2850_ (.A(_1285_),
    .X(_0098_));
 sky130_fd_sc_hd__mux2_1 _2851_ (.A0(\tms1x00.RAM[104][2] ),
    .A1(_1273_),
    .S(_1283_),
    .X(_1286_));
 sky130_fd_sc_hd__clkbuf_1 _2852_ (.A(_1286_),
    .X(_0099_));
 sky130_fd_sc_hd__mux2_1 _2853_ (.A0(\tms1x00.RAM[104][3] ),
    .A1(_1276_),
    .S(_1283_),
    .X(_1287_));
 sky130_fd_sc_hd__clkbuf_1 _2854_ (.A(_1287_),
    .X(_0100_));
 sky130_fd_sc_hd__nor2_2 _2855_ (.A(_0829_),
    .B(_1257_),
    .Y(_1288_));
 sky130_fd_sc_hd__mux2_1 _2856_ (.A0(\tms1x00.RAM[103][0] ),
    .A1(_1264_),
    .S(_1288_),
    .X(_1289_));
 sky130_fd_sc_hd__clkbuf_1 _2857_ (.A(_1289_),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _2858_ (.A0(\tms1x00.RAM[103][1] ),
    .A1(_1270_),
    .S(_1288_),
    .X(_1290_));
 sky130_fd_sc_hd__clkbuf_1 _2859_ (.A(_1290_),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_1 _2860_ (.A0(\tms1x00.RAM[103][2] ),
    .A1(_1273_),
    .S(_1288_),
    .X(_1291_));
 sky130_fd_sc_hd__clkbuf_1 _2861_ (.A(_1291_),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _2862_ (.A0(\tms1x00.RAM[103][3] ),
    .A1(_1276_),
    .S(_1288_),
    .X(_1292_));
 sky130_fd_sc_hd__clkbuf_1 _2863_ (.A(_1292_),
    .X(_0104_));
 sky130_fd_sc_hd__nor2_2 _2864_ (.A(_0829_),
    .B(_1266_),
    .Y(_1293_));
 sky130_fd_sc_hd__mux2_1 _2865_ (.A0(\tms1x00.RAM[102][0] ),
    .A1(_1264_),
    .S(_1293_),
    .X(_1294_));
 sky130_fd_sc_hd__clkbuf_1 _2866_ (.A(_1294_),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _2867_ (.A0(\tms1x00.RAM[102][1] ),
    .A1(_1270_),
    .S(_1293_),
    .X(_1295_));
 sky130_fd_sc_hd__clkbuf_1 _2868_ (.A(_1295_),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _2869_ (.A0(\tms1x00.RAM[102][2] ),
    .A1(_1273_),
    .S(_1293_),
    .X(_1296_));
 sky130_fd_sc_hd__clkbuf_1 _2870_ (.A(_1296_),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _2871_ (.A0(\tms1x00.RAM[102][3] ),
    .A1(_1276_),
    .S(_1293_),
    .X(_1297_));
 sky130_fd_sc_hd__clkbuf_1 _2872_ (.A(_1297_),
    .X(_0108_));
 sky130_fd_sc_hd__nor2_2 _2873_ (.A(_0829_),
    .B(_1180_),
    .Y(_1298_));
 sky130_fd_sc_hd__mux2_1 _2874_ (.A0(\tms1x00.RAM[101][0] ),
    .A1(_1264_),
    .S(_1298_),
    .X(_1299_));
 sky130_fd_sc_hd__clkbuf_1 _2875_ (.A(_1299_),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _2876_ (.A0(\tms1x00.RAM[101][1] ),
    .A1(_1270_),
    .S(_1298_),
    .X(_1300_));
 sky130_fd_sc_hd__clkbuf_1 _2877_ (.A(_1300_),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_1 _2878_ (.A0(\tms1x00.RAM[101][2] ),
    .A1(_1273_),
    .S(_1298_),
    .X(_1301_));
 sky130_fd_sc_hd__clkbuf_1 _2879_ (.A(_1301_),
    .X(_0111_));
 sky130_fd_sc_hd__mux2_1 _2880_ (.A0(\tms1x00.RAM[101][3] ),
    .A1(_1276_),
    .S(_1298_),
    .X(_1302_));
 sky130_fd_sc_hd__clkbuf_1 _2881_ (.A(_1302_),
    .X(_0112_));
 sky130_fd_sc_hd__or3_1 _2882_ (.A(\tms1x00.ram_addr_buff[0] ),
    .B(\tms1x00.ram_addr_buff[1] ),
    .C(_1178_),
    .X(_1303_));
 sky130_fd_sc_hd__buf_6 _2883_ (.A(_1303_),
    .X(_1304_));
 sky130_fd_sc_hd__nor2_2 _2884_ (.A(_0829_),
    .B(_1304_),
    .Y(_1305_));
 sky130_fd_sc_hd__mux2_1 _2885_ (.A0(\tms1x00.RAM[100][0] ),
    .A1(_1264_),
    .S(_1305_),
    .X(_1306_));
 sky130_fd_sc_hd__clkbuf_1 _2886_ (.A(_1306_),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _2887_ (.A0(\tms1x00.RAM[100][1] ),
    .A1(_1270_),
    .S(_1305_),
    .X(_1307_));
 sky130_fd_sc_hd__clkbuf_1 _2888_ (.A(_1307_),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_1 _2889_ (.A0(\tms1x00.RAM[100][2] ),
    .A1(_1273_),
    .S(_1305_),
    .X(_1308_));
 sky130_fd_sc_hd__clkbuf_1 _2890_ (.A(_1308_),
    .X(_0115_));
 sky130_fd_sc_hd__mux2_1 _2891_ (.A0(\tms1x00.RAM[100][3] ),
    .A1(_1276_),
    .S(_1305_),
    .X(_1309_));
 sky130_fd_sc_hd__clkbuf_1 _2892_ (.A(_1309_),
    .X(_0116_));
 sky130_fd_sc_hd__buf_2 _2893_ (.A(_0826_),
    .X(_1310_));
 sky130_fd_sc_hd__or3_4 _2894_ (.A(_0620_),
    .B(_0628_),
    .C(_0831_),
    .X(_1311_));
 sky130_fd_sc_hd__or2_2 _2895_ (.A(_1243_),
    .B(_1311_),
    .X(_1312_));
 sky130_fd_sc_hd__mux2_1 _2896_ (.A0(_1310_),
    .A1(\tms1x00.RAM[0][0] ),
    .S(_1312_),
    .X(_1313_));
 sky130_fd_sc_hd__clkbuf_1 _2897_ (.A(_1313_),
    .X(_0117_));
 sky130_fd_sc_hd__buf_2 _2898_ (.A(_0934_),
    .X(_1314_));
 sky130_fd_sc_hd__mux2_1 _2899_ (.A0(_1314_),
    .A1(\tms1x00.RAM[0][1] ),
    .S(_1312_),
    .X(_1315_));
 sky130_fd_sc_hd__clkbuf_1 _2900_ (.A(_1315_),
    .X(_0118_));
 sky130_fd_sc_hd__buf_2 _2901_ (.A(_1034_),
    .X(_1316_));
 sky130_fd_sc_hd__mux2_1 _2902_ (.A0(_1316_),
    .A1(\tms1x00.RAM[0][2] ),
    .S(_1312_),
    .X(_1317_));
 sky130_fd_sc_hd__clkbuf_1 _2903_ (.A(_1317_),
    .X(_0119_));
 sky130_fd_sc_hd__buf_2 _2904_ (.A(_1132_),
    .X(_1318_));
 sky130_fd_sc_hd__mux2_1 _2905_ (.A0(_1318_),
    .A1(\tms1x00.RAM[0][3] ),
    .S(_1312_),
    .X(_1319_));
 sky130_fd_sc_hd__clkbuf_1 _2906_ (.A(_1319_),
    .X(_0120_));
 sky130_fd_sc_hd__or3b_4 _2907_ (.A(_0831_),
    .B(_0620_),
    .C_N(_0628_),
    .X(_1320_));
 sky130_fd_sc_hd__or2_2 _2908_ (.A(_0829_),
    .B(_1320_),
    .X(_1321_));
 sky130_fd_sc_hd__mux2_1 _2909_ (.A0(_1310_),
    .A1(\tms1x00.RAM[98][0] ),
    .S(_1321_),
    .X(_1322_));
 sky130_fd_sc_hd__clkbuf_1 _2910_ (.A(_1322_),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _2911_ (.A0(_1314_),
    .A1(\tms1x00.RAM[98][1] ),
    .S(_1321_),
    .X(_1323_));
 sky130_fd_sc_hd__clkbuf_1 _2912_ (.A(_1323_),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _2913_ (.A0(_1316_),
    .A1(\tms1x00.RAM[98][2] ),
    .S(_1321_),
    .X(_1324_));
 sky130_fd_sc_hd__clkbuf_1 _2914_ (.A(_1324_),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _2915_ (.A0(_1318_),
    .A1(\tms1x00.RAM[98][3] ),
    .S(_1321_),
    .X(_1325_));
 sky130_fd_sc_hd__clkbuf_1 _2916_ (.A(_1325_),
    .X(_0124_));
 sky130_fd_sc_hd__or2_2 _2917_ (.A(_0828_),
    .B(_1194_),
    .X(_1326_));
 sky130_fd_sc_hd__mux2_1 _2918_ (.A0(_1310_),
    .A1(\tms1x00.RAM[97][0] ),
    .S(_1326_),
    .X(_1327_));
 sky130_fd_sc_hd__clkbuf_1 _2919_ (.A(_1327_),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_1 _2920_ (.A0(_1314_),
    .A1(\tms1x00.RAM[97][1] ),
    .S(_1326_),
    .X(_1328_));
 sky130_fd_sc_hd__clkbuf_1 _2921_ (.A(_1328_),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_1 _2922_ (.A0(_1316_),
    .A1(\tms1x00.RAM[97][2] ),
    .S(_1326_),
    .X(_1329_));
 sky130_fd_sc_hd__clkbuf_1 _2923_ (.A(_1329_),
    .X(_0127_));
 sky130_fd_sc_hd__mux2_1 _2924_ (.A0(_1318_),
    .A1(\tms1x00.RAM[97][3] ),
    .S(_1326_),
    .X(_1330_));
 sky130_fd_sc_hd__clkbuf_1 _2925_ (.A(_1330_),
    .X(_0128_));
 sky130_fd_sc_hd__or2_2 _2926_ (.A(_0828_),
    .B(_1311_),
    .X(_1331_));
 sky130_fd_sc_hd__mux2_1 _2927_ (.A0(_1310_),
    .A1(\tms1x00.RAM[96][0] ),
    .S(_1331_),
    .X(_1332_));
 sky130_fd_sc_hd__clkbuf_1 _2928_ (.A(_1332_),
    .X(_0129_));
 sky130_fd_sc_hd__mux2_1 _2929_ (.A0(_1314_),
    .A1(\tms1x00.RAM[96][1] ),
    .S(_1331_),
    .X(_1333_));
 sky130_fd_sc_hd__clkbuf_1 _2930_ (.A(_1333_),
    .X(_0130_));
 sky130_fd_sc_hd__mux2_1 _2931_ (.A0(_1316_),
    .A1(\tms1x00.RAM[96][2] ),
    .S(_1331_),
    .X(_1334_));
 sky130_fd_sc_hd__clkbuf_1 _2932_ (.A(_1334_),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_1 _2933_ (.A0(_1318_),
    .A1(\tms1x00.RAM[96][3] ),
    .S(_1331_),
    .X(_1335_));
 sky130_fd_sc_hd__clkbuf_1 _2934_ (.A(_1335_),
    .X(_0132_));
 sky130_fd_sc_hd__nand3_1 _2935_ (.A(_0635_),
    .B(_0637_),
    .C(\tms1x00.ram_addr_buff[6] ),
    .Y(_1336_));
 sky130_fd_sc_hd__buf_2 _2936_ (.A(_1336_),
    .X(_1337_));
 sky130_fd_sc_hd__or2_2 _2937_ (.A(_0833_),
    .B(_1337_),
    .X(_1338_));
 sky130_fd_sc_hd__mux2_1 _2938_ (.A0(_1310_),
    .A1(\tms1x00.RAM[115][0] ),
    .S(_1338_),
    .X(_1339_));
 sky130_fd_sc_hd__clkbuf_1 _2939_ (.A(_1339_),
    .X(_0133_));
 sky130_fd_sc_hd__mux2_1 _2940_ (.A0(_1314_),
    .A1(\tms1x00.RAM[115][1] ),
    .S(_1338_),
    .X(_1340_));
 sky130_fd_sc_hd__clkbuf_1 _2941_ (.A(_1340_),
    .X(_0134_));
 sky130_fd_sc_hd__mux2_1 _2942_ (.A0(_1316_),
    .A1(\tms1x00.RAM[115][2] ),
    .S(_1338_),
    .X(_1341_));
 sky130_fd_sc_hd__clkbuf_1 _2943_ (.A(_1341_),
    .X(_0135_));
 sky130_fd_sc_hd__mux2_1 _2944_ (.A0(_1318_),
    .A1(\tms1x00.RAM[115][3] ),
    .S(_1338_),
    .X(_1342_));
 sky130_fd_sc_hd__clkbuf_1 _2945_ (.A(_1342_),
    .X(_0136_));
 sky130_fd_sc_hd__or2_2 _2946_ (.A(_1337_),
    .B(_1320_),
    .X(_1343_));
 sky130_fd_sc_hd__mux2_1 _2947_ (.A0(_1310_),
    .A1(\tms1x00.RAM[114][0] ),
    .S(_1343_),
    .X(_1344_));
 sky130_fd_sc_hd__clkbuf_1 _2948_ (.A(_1344_),
    .X(_0137_));
 sky130_fd_sc_hd__mux2_1 _2949_ (.A0(_1314_),
    .A1(\tms1x00.RAM[114][1] ),
    .S(_1343_),
    .X(_1345_));
 sky130_fd_sc_hd__clkbuf_1 _2950_ (.A(_1345_),
    .X(_0138_));
 sky130_fd_sc_hd__mux2_1 _2951_ (.A0(_1316_),
    .A1(\tms1x00.RAM[114][2] ),
    .S(_1343_),
    .X(_1346_));
 sky130_fd_sc_hd__clkbuf_1 _2952_ (.A(_1346_),
    .X(_0139_));
 sky130_fd_sc_hd__mux2_1 _2953_ (.A0(_1318_),
    .A1(\tms1x00.RAM[114][3] ),
    .S(_1343_),
    .X(_1347_));
 sky130_fd_sc_hd__clkbuf_1 _2954_ (.A(_1347_),
    .X(_0140_));
 sky130_fd_sc_hd__or2_2 _2955_ (.A(_1337_),
    .B(_1194_),
    .X(_1348_));
 sky130_fd_sc_hd__mux2_1 _2956_ (.A0(_1310_),
    .A1(\tms1x00.RAM[113][0] ),
    .S(_1348_),
    .X(_1349_));
 sky130_fd_sc_hd__clkbuf_1 _2957_ (.A(_1349_),
    .X(_0141_));
 sky130_fd_sc_hd__mux2_1 _2958_ (.A0(_1314_),
    .A1(\tms1x00.RAM[113][1] ),
    .S(_1348_),
    .X(_1350_));
 sky130_fd_sc_hd__clkbuf_1 _2959_ (.A(_1350_),
    .X(_0142_));
 sky130_fd_sc_hd__mux2_1 _2960_ (.A0(_1316_),
    .A1(\tms1x00.RAM[113][2] ),
    .S(_1348_),
    .X(_1351_));
 sky130_fd_sc_hd__clkbuf_1 _2961_ (.A(_1351_),
    .X(_0143_));
 sky130_fd_sc_hd__mux2_1 _2962_ (.A0(_1318_),
    .A1(\tms1x00.RAM[113][3] ),
    .S(_1348_),
    .X(_1352_));
 sky130_fd_sc_hd__clkbuf_1 _2963_ (.A(_1352_),
    .X(_0144_));
 sky130_fd_sc_hd__or2_2 _2964_ (.A(_1337_),
    .B(_1311_),
    .X(_1353_));
 sky130_fd_sc_hd__mux2_1 _2965_ (.A0(_1310_),
    .A1(\tms1x00.RAM[112][0] ),
    .S(_1353_),
    .X(_1354_));
 sky130_fd_sc_hd__clkbuf_1 _2966_ (.A(_1354_),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _2967_ (.A0(_1314_),
    .A1(\tms1x00.RAM[112][1] ),
    .S(_1353_),
    .X(_1355_));
 sky130_fd_sc_hd__clkbuf_1 _2968_ (.A(_1355_),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_1 _2969_ (.A0(_1316_),
    .A1(\tms1x00.RAM[112][2] ),
    .S(_1353_),
    .X(_1356_));
 sky130_fd_sc_hd__clkbuf_1 _2970_ (.A(_1356_),
    .X(_0147_));
 sky130_fd_sc_hd__mux2_1 _2971_ (.A0(_1318_),
    .A1(\tms1x00.RAM[112][3] ),
    .S(_1353_),
    .X(_1357_));
 sky130_fd_sc_hd__clkbuf_1 _2972_ (.A(_1357_),
    .X(_0148_));
 sky130_fd_sc_hd__nand2_2 _2973_ (.A(_1159_),
    .B(_1170_),
    .Y(_1358_));
 sky130_fd_sc_hd__mux2_1 _2974_ (.A0(_1310_),
    .A1(\tms1x00.RAM[111][0] ),
    .S(_1358_),
    .X(_1359_));
 sky130_fd_sc_hd__clkbuf_1 _2975_ (.A(_1359_),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_1 _2976_ (.A0(_1314_),
    .A1(\tms1x00.RAM[111][1] ),
    .S(_1358_),
    .X(_1360_));
 sky130_fd_sc_hd__clkbuf_1 _2977_ (.A(_1360_),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_1 _2978_ (.A0(_1316_),
    .A1(\tms1x00.RAM[111][2] ),
    .S(_1358_),
    .X(_1361_));
 sky130_fd_sc_hd__clkbuf_1 _2979_ (.A(_1361_),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _2980_ (.A0(_1318_),
    .A1(\tms1x00.RAM[111][3] ),
    .S(_1358_),
    .X(_1362_));
 sky130_fd_sc_hd__clkbuf_1 _2981_ (.A(_1362_),
    .X(_0152_));
 sky130_fd_sc_hd__nand2_2 _2982_ (.A(_1159_),
    .B(_1213_),
    .Y(_1363_));
 sky130_fd_sc_hd__mux2_1 _2983_ (.A0(_1310_),
    .A1(\tms1x00.RAM[110][0] ),
    .S(_1363_),
    .X(_1364_));
 sky130_fd_sc_hd__clkbuf_1 _2984_ (.A(_1364_),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _2985_ (.A0(_1314_),
    .A1(\tms1x00.RAM[110][1] ),
    .S(_1363_),
    .X(_1365_));
 sky130_fd_sc_hd__clkbuf_1 _2986_ (.A(_1365_),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_1 _2987_ (.A0(_1316_),
    .A1(\tms1x00.RAM[110][2] ),
    .S(_1363_),
    .X(_1366_));
 sky130_fd_sc_hd__clkbuf_1 _2988_ (.A(_1366_),
    .X(_0155_));
 sky130_fd_sc_hd__mux2_1 _2989_ (.A0(_1318_),
    .A1(\tms1x00.RAM[110][3] ),
    .S(_1363_),
    .X(_1367_));
 sky130_fd_sc_hd__clkbuf_1 _2990_ (.A(_1367_),
    .X(_0156_));
 sky130_fd_sc_hd__nor2_2 _2991_ (.A(_1236_),
    .B(_1243_),
    .Y(_1368_));
 sky130_fd_sc_hd__mux2_1 _2992_ (.A0(\tms1x00.RAM[10][0] ),
    .A1(_1264_),
    .S(_1368_),
    .X(_1369_));
 sky130_fd_sc_hd__clkbuf_1 _2993_ (.A(_1369_),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_1 _2994_ (.A0(\tms1x00.RAM[10][1] ),
    .A1(_1270_),
    .S(_1368_),
    .X(_1370_));
 sky130_fd_sc_hd__clkbuf_1 _2995_ (.A(_1370_),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_1 _2996_ (.A0(\tms1x00.RAM[10][2] ),
    .A1(_1273_),
    .S(_1368_),
    .X(_1371_));
 sky130_fd_sc_hd__clkbuf_1 _2997_ (.A(_1371_),
    .X(_0159_));
 sky130_fd_sc_hd__mux2_1 _2998_ (.A0(\tms1x00.RAM[10][3] ),
    .A1(_1276_),
    .S(_1368_),
    .X(_1372_));
 sky130_fd_sc_hd__clkbuf_1 _2999_ (.A(_1372_),
    .X(_0160_));
 sky130_fd_sc_hd__buf_2 _3000_ (.A(_0826_),
    .X(_1373_));
 sky130_fd_sc_hd__nand2_2 _3001_ (.A(_1159_),
    .B(_1224_),
    .Y(_1374_));
 sky130_fd_sc_hd__mux2_1 _3002_ (.A0(_1373_),
    .A1(\tms1x00.RAM[108][0] ),
    .S(_1374_),
    .X(_1375_));
 sky130_fd_sc_hd__clkbuf_1 _3003_ (.A(_1375_),
    .X(_0161_));
 sky130_fd_sc_hd__buf_2 _3004_ (.A(_0934_),
    .X(_1376_));
 sky130_fd_sc_hd__mux2_1 _3005_ (.A0(_1376_),
    .A1(\tms1x00.RAM[108][1] ),
    .S(_1374_),
    .X(_1377_));
 sky130_fd_sc_hd__clkbuf_1 _3006_ (.A(_1377_),
    .X(_0162_));
 sky130_fd_sc_hd__buf_2 _3007_ (.A(_1034_),
    .X(_1378_));
 sky130_fd_sc_hd__mux2_1 _3008_ (.A0(_1378_),
    .A1(\tms1x00.RAM[108][2] ),
    .S(_1374_),
    .X(_1379_));
 sky130_fd_sc_hd__clkbuf_1 _3009_ (.A(_1379_),
    .X(_0163_));
 sky130_fd_sc_hd__clkbuf_4 _3010_ (.A(_1132_),
    .X(_1380_));
 sky130_fd_sc_hd__mux2_1 _3011_ (.A0(_1380_),
    .A1(\tms1x00.RAM[108][3] ),
    .S(_1374_),
    .X(_1381_));
 sky130_fd_sc_hd__clkbuf_1 _3012_ (.A(_1381_),
    .X(_0164_));
 sky130_fd_sc_hd__nor2_2 _3013_ (.A(_0829_),
    .B(_1153_),
    .Y(_1382_));
 sky130_fd_sc_hd__mux2_1 _3014_ (.A0(\tms1x00.RAM[107][0] ),
    .A1(_1264_),
    .S(_1382_),
    .X(_1383_));
 sky130_fd_sc_hd__clkbuf_1 _3015_ (.A(_1383_),
    .X(_0165_));
 sky130_fd_sc_hd__mux2_1 _3016_ (.A0(\tms1x00.RAM[107][1] ),
    .A1(_1270_),
    .S(_1382_),
    .X(_1384_));
 sky130_fd_sc_hd__clkbuf_1 _3017_ (.A(_1384_),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_1 _3018_ (.A0(\tms1x00.RAM[107][2] ),
    .A1(_1273_),
    .S(_1382_),
    .X(_1385_));
 sky130_fd_sc_hd__clkbuf_1 _3019_ (.A(_1385_),
    .X(_0167_));
 sky130_fd_sc_hd__mux2_1 _3020_ (.A0(\tms1x00.RAM[107][3] ),
    .A1(_1276_),
    .S(_1382_),
    .X(_1386_));
 sky130_fd_sc_hd__clkbuf_1 _3021_ (.A(_1386_),
    .X(_0168_));
 sky130_fd_sc_hd__nor2_2 _3022_ (.A(_0829_),
    .B(_1236_),
    .Y(_1387_));
 sky130_fd_sc_hd__mux2_1 _3023_ (.A0(\tms1x00.RAM[106][0] ),
    .A1(_1264_),
    .S(_1387_),
    .X(_1388_));
 sky130_fd_sc_hd__clkbuf_1 _3024_ (.A(_1388_),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_1 _3025_ (.A0(\tms1x00.RAM[106][1] ),
    .A1(_1270_),
    .S(_1387_),
    .X(_1389_));
 sky130_fd_sc_hd__clkbuf_1 _3026_ (.A(_1389_),
    .X(_0170_));
 sky130_fd_sc_hd__mux2_1 _3027_ (.A0(\tms1x00.RAM[106][2] ),
    .A1(_1273_),
    .S(_1387_),
    .X(_1390_));
 sky130_fd_sc_hd__clkbuf_1 _3028_ (.A(_1390_),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _3029_ (.A0(\tms1x00.RAM[106][3] ),
    .A1(_1276_),
    .S(_1387_),
    .X(_1391_));
 sky130_fd_sc_hd__clkbuf_1 _3030_ (.A(_1391_),
    .X(_0172_));
 sky130_fd_sc_hd__nand2_2 _3031_ (.A(_1162_),
    .B(_1186_),
    .Y(_1392_));
 sky130_fd_sc_hd__mux2_1 _3032_ (.A0(_1373_),
    .A1(\tms1x00.RAM[125][0] ),
    .S(_1392_),
    .X(_1393_));
 sky130_fd_sc_hd__clkbuf_1 _3033_ (.A(_1393_),
    .X(_0173_));
 sky130_fd_sc_hd__mux2_1 _3034_ (.A0(_1376_),
    .A1(\tms1x00.RAM[125][1] ),
    .S(_1392_),
    .X(_1394_));
 sky130_fd_sc_hd__clkbuf_1 _3035_ (.A(_1394_),
    .X(_0174_));
 sky130_fd_sc_hd__mux2_1 _3036_ (.A0(_1378_),
    .A1(\tms1x00.RAM[125][2] ),
    .S(_1392_),
    .X(_1395_));
 sky130_fd_sc_hd__clkbuf_1 _3037_ (.A(_1395_),
    .X(_0175_));
 sky130_fd_sc_hd__mux2_1 _3038_ (.A0(_1380_),
    .A1(\tms1x00.RAM[125][3] ),
    .S(_1392_),
    .X(_1396_));
 sky130_fd_sc_hd__clkbuf_1 _3039_ (.A(_1396_),
    .X(_0176_));
 sky130_fd_sc_hd__nand2_2 _3040_ (.A(_1186_),
    .B(_1224_),
    .Y(_1397_));
 sky130_fd_sc_hd__mux2_1 _3041_ (.A0(_1373_),
    .A1(\tms1x00.RAM[124][0] ),
    .S(_1397_),
    .X(_1398_));
 sky130_fd_sc_hd__clkbuf_1 _3042_ (.A(_1398_),
    .X(_0177_));
 sky130_fd_sc_hd__mux2_1 _3043_ (.A0(_1376_),
    .A1(\tms1x00.RAM[124][1] ),
    .S(_1397_),
    .X(_1399_));
 sky130_fd_sc_hd__clkbuf_1 _3044_ (.A(_1399_),
    .X(_0178_));
 sky130_fd_sc_hd__mux2_1 _3045_ (.A0(_1378_),
    .A1(\tms1x00.RAM[124][2] ),
    .S(_1397_),
    .X(_1400_));
 sky130_fd_sc_hd__clkbuf_1 _3046_ (.A(_1400_),
    .X(_0179_));
 sky130_fd_sc_hd__mux2_1 _3047_ (.A0(_1380_),
    .A1(\tms1x00.RAM[124][3] ),
    .S(_1397_),
    .X(_1401_));
 sky130_fd_sc_hd__clkbuf_1 _3048_ (.A(_1401_),
    .X(_0180_));
 sky130_fd_sc_hd__or2_2 _3049_ (.A(_1153_),
    .B(_1337_),
    .X(_1402_));
 sky130_fd_sc_hd__mux2_1 _3050_ (.A0(_1373_),
    .A1(\tms1x00.RAM[123][0] ),
    .S(_1402_),
    .X(_1403_));
 sky130_fd_sc_hd__clkbuf_1 _3051_ (.A(_1403_),
    .X(_0181_));
 sky130_fd_sc_hd__mux2_1 _3052_ (.A0(_1376_),
    .A1(\tms1x00.RAM[123][1] ),
    .S(_1402_),
    .X(_1404_));
 sky130_fd_sc_hd__clkbuf_1 _3053_ (.A(_1404_),
    .X(_0182_));
 sky130_fd_sc_hd__mux2_1 _3054_ (.A0(_1378_),
    .A1(\tms1x00.RAM[123][2] ),
    .S(_1402_),
    .X(_1405_));
 sky130_fd_sc_hd__clkbuf_1 _3055_ (.A(_1405_),
    .X(_0183_));
 sky130_fd_sc_hd__mux2_1 _3056_ (.A0(_1380_),
    .A1(\tms1x00.RAM[123][3] ),
    .S(_1402_),
    .X(_1406_));
 sky130_fd_sc_hd__clkbuf_1 _3057_ (.A(_1406_),
    .X(_0184_));
 sky130_fd_sc_hd__or2_2 _3058_ (.A(_1337_),
    .B(_1236_),
    .X(_1407_));
 sky130_fd_sc_hd__mux2_1 _3059_ (.A0(_1373_),
    .A1(\tms1x00.RAM[122][0] ),
    .S(_1407_),
    .X(_1408_));
 sky130_fd_sc_hd__clkbuf_1 _3060_ (.A(_1408_),
    .X(_0185_));
 sky130_fd_sc_hd__mux2_1 _3061_ (.A0(_1376_),
    .A1(\tms1x00.RAM[122][1] ),
    .S(_1407_),
    .X(_1409_));
 sky130_fd_sc_hd__clkbuf_1 _3062_ (.A(_1409_),
    .X(_0186_));
 sky130_fd_sc_hd__mux2_1 _3063_ (.A0(_1378_),
    .A1(\tms1x00.RAM[122][2] ),
    .S(_1407_),
    .X(_1410_));
 sky130_fd_sc_hd__clkbuf_1 _3064_ (.A(_1410_),
    .X(_0187_));
 sky130_fd_sc_hd__mux2_1 _3065_ (.A0(_1380_),
    .A1(\tms1x00.RAM[122][3] ),
    .S(_1407_),
    .X(_1411_));
 sky130_fd_sc_hd__clkbuf_1 _3066_ (.A(_1411_),
    .X(_0188_));
 sky130_fd_sc_hd__or2_2 _3067_ (.A(_1140_),
    .B(_1336_),
    .X(_1412_));
 sky130_fd_sc_hd__mux2_1 _3068_ (.A0(_1373_),
    .A1(\tms1x00.RAM[121][0] ),
    .S(_1412_),
    .X(_1413_));
 sky130_fd_sc_hd__clkbuf_1 _3069_ (.A(_1413_),
    .X(_0189_));
 sky130_fd_sc_hd__mux2_1 _3070_ (.A0(_1376_),
    .A1(\tms1x00.RAM[121][1] ),
    .S(_1412_),
    .X(_1414_));
 sky130_fd_sc_hd__clkbuf_1 _3071_ (.A(_1414_),
    .X(_0190_));
 sky130_fd_sc_hd__mux2_1 _3072_ (.A0(_1378_),
    .A1(\tms1x00.RAM[121][2] ),
    .S(_1412_),
    .X(_1415_));
 sky130_fd_sc_hd__clkbuf_1 _3073_ (.A(_1415_),
    .X(_0191_));
 sky130_fd_sc_hd__mux2_1 _3074_ (.A0(_1380_),
    .A1(\tms1x00.RAM[121][3] ),
    .S(_1412_),
    .X(_1416_));
 sky130_fd_sc_hd__clkbuf_1 _3075_ (.A(_1416_),
    .X(_0192_));
 sky130_fd_sc_hd__or2_2 _3076_ (.A(_1337_),
    .B(_1245_),
    .X(_1417_));
 sky130_fd_sc_hd__mux2_1 _3077_ (.A0(_1373_),
    .A1(\tms1x00.RAM[120][0] ),
    .S(_1417_),
    .X(_1418_));
 sky130_fd_sc_hd__clkbuf_1 _3078_ (.A(_1418_),
    .X(_0193_));
 sky130_fd_sc_hd__mux2_1 _3079_ (.A0(_1376_),
    .A1(\tms1x00.RAM[120][1] ),
    .S(_1417_),
    .X(_1419_));
 sky130_fd_sc_hd__clkbuf_1 _3080_ (.A(_1419_),
    .X(_0194_));
 sky130_fd_sc_hd__mux2_1 _3081_ (.A0(_1378_),
    .A1(\tms1x00.RAM[120][2] ),
    .S(_1417_),
    .X(_1420_));
 sky130_fd_sc_hd__clkbuf_1 _3082_ (.A(_1420_),
    .X(_0195_));
 sky130_fd_sc_hd__mux2_1 _3083_ (.A0(_1380_),
    .A1(\tms1x00.RAM[120][3] ),
    .S(_1417_),
    .X(_1421_));
 sky130_fd_sc_hd__clkbuf_1 _3084_ (.A(_1421_),
    .X(_0196_));
 sky130_fd_sc_hd__clkbuf_4 _3085_ (.A(_1263_),
    .X(_1422_));
 sky130_fd_sc_hd__nor2_2 _3086_ (.A(_1153_),
    .B(_1243_),
    .Y(_1423_));
 sky130_fd_sc_hd__mux2_1 _3087_ (.A0(\tms1x00.RAM[11][0] ),
    .A1(_1422_),
    .S(_1423_),
    .X(_1424_));
 sky130_fd_sc_hd__clkbuf_1 _3088_ (.A(_1424_),
    .X(_0197_));
 sky130_fd_sc_hd__clkbuf_4 _3089_ (.A(_1269_),
    .X(_1425_));
 sky130_fd_sc_hd__mux2_1 _3090_ (.A0(\tms1x00.RAM[11][1] ),
    .A1(_1425_),
    .S(_1423_),
    .X(_1426_));
 sky130_fd_sc_hd__clkbuf_1 _3091_ (.A(_1426_),
    .X(_0198_));
 sky130_fd_sc_hd__clkbuf_4 _3092_ (.A(_1272_),
    .X(_1427_));
 sky130_fd_sc_hd__mux2_1 _3093_ (.A0(\tms1x00.RAM[11][2] ),
    .A1(_1427_),
    .S(_1423_),
    .X(_1428_));
 sky130_fd_sc_hd__clkbuf_1 _3094_ (.A(_1428_),
    .X(_0199_));
 sky130_fd_sc_hd__clkbuf_4 _3095_ (.A(_1275_),
    .X(_1429_));
 sky130_fd_sc_hd__mux2_1 _3096_ (.A0(\tms1x00.RAM[11][3] ),
    .A1(_1429_),
    .S(_1423_),
    .X(_1430_));
 sky130_fd_sc_hd__clkbuf_1 _3097_ (.A(_1430_),
    .X(_0200_));
 sky130_fd_sc_hd__or2_2 _3098_ (.A(_1337_),
    .B(_1266_),
    .X(_1431_));
 sky130_fd_sc_hd__mux2_1 _3099_ (.A0(_1373_),
    .A1(\tms1x00.RAM[118][0] ),
    .S(_1431_),
    .X(_1432_));
 sky130_fd_sc_hd__clkbuf_1 _3100_ (.A(_1432_),
    .X(_0201_));
 sky130_fd_sc_hd__mux2_1 _3101_ (.A0(_1376_),
    .A1(\tms1x00.RAM[118][1] ),
    .S(_1431_),
    .X(_1433_));
 sky130_fd_sc_hd__clkbuf_1 _3102_ (.A(_1433_),
    .X(_0202_));
 sky130_fd_sc_hd__mux2_1 _3103_ (.A0(_1378_),
    .A1(\tms1x00.RAM[118][2] ),
    .S(_1431_),
    .X(_1434_));
 sky130_fd_sc_hd__clkbuf_1 _3104_ (.A(_1434_),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_1 _3105_ (.A0(_1380_),
    .A1(\tms1x00.RAM[118][3] ),
    .S(_1431_),
    .X(_1435_));
 sky130_fd_sc_hd__clkbuf_1 _3106_ (.A(_1435_),
    .X(_0204_));
 sky130_fd_sc_hd__or2_2 _3107_ (.A(_1180_),
    .B(_1336_),
    .X(_1436_));
 sky130_fd_sc_hd__mux2_1 _3108_ (.A0(_1373_),
    .A1(\tms1x00.RAM[117][0] ),
    .S(_1436_),
    .X(_1437_));
 sky130_fd_sc_hd__clkbuf_1 _3109_ (.A(_1437_),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _3110_ (.A0(_1376_),
    .A1(\tms1x00.RAM[117][1] ),
    .S(_1436_),
    .X(_1438_));
 sky130_fd_sc_hd__clkbuf_1 _3111_ (.A(_1438_),
    .X(_0206_));
 sky130_fd_sc_hd__mux2_1 _3112_ (.A0(_1378_),
    .A1(\tms1x00.RAM[117][2] ),
    .S(_1436_),
    .X(_1439_));
 sky130_fd_sc_hd__clkbuf_1 _3113_ (.A(_1439_),
    .X(_0207_));
 sky130_fd_sc_hd__mux2_1 _3114_ (.A0(_1380_),
    .A1(\tms1x00.RAM[117][3] ),
    .S(_1436_),
    .X(_1440_));
 sky130_fd_sc_hd__clkbuf_1 _3115_ (.A(_1440_),
    .X(_0208_));
 sky130_fd_sc_hd__or2_2 _3116_ (.A(_1337_),
    .B(_1304_),
    .X(_1441_));
 sky130_fd_sc_hd__mux2_1 _3117_ (.A0(_1373_),
    .A1(\tms1x00.RAM[116][0] ),
    .S(_1441_),
    .X(_1442_));
 sky130_fd_sc_hd__clkbuf_1 _3118_ (.A(_1442_),
    .X(_0209_));
 sky130_fd_sc_hd__mux2_1 _3119_ (.A0(_1376_),
    .A1(\tms1x00.RAM[116][1] ),
    .S(_1441_),
    .X(_1443_));
 sky130_fd_sc_hd__clkbuf_1 _3120_ (.A(_1443_),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_1 _3121_ (.A0(_1378_),
    .A1(\tms1x00.RAM[116][2] ),
    .S(_1441_),
    .X(_1444_));
 sky130_fd_sc_hd__clkbuf_1 _3122_ (.A(_1444_),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_1 _3123_ (.A0(_1380_),
    .A1(\tms1x00.RAM[116][3] ),
    .S(_1441_),
    .X(_1445_));
 sky130_fd_sc_hd__clkbuf_1 _3124_ (.A(_1445_),
    .X(_0212_));
 sky130_fd_sc_hd__buf_2 _3125_ (.A(_0826_),
    .X(_1446_));
 sky130_fd_sc_hd__nand2_2 _3126_ (.A(_1186_),
    .B(_1213_),
    .Y(_1447_));
 sky130_fd_sc_hd__mux2_1 _3127_ (.A0(_1446_),
    .A1(\tms1x00.RAM[126][0] ),
    .S(_1447_),
    .X(_1448_));
 sky130_fd_sc_hd__clkbuf_1 _3128_ (.A(_1448_),
    .X(_0213_));
 sky130_fd_sc_hd__clkbuf_4 _3129_ (.A(_0934_),
    .X(_1449_));
 sky130_fd_sc_hd__mux2_1 _3130_ (.A0(_1449_),
    .A1(\tms1x00.RAM[126][1] ),
    .S(_1447_),
    .X(_1450_));
 sky130_fd_sc_hd__clkbuf_1 _3131_ (.A(_1450_),
    .X(_0214_));
 sky130_fd_sc_hd__clkbuf_4 _3132_ (.A(_1034_),
    .X(_1451_));
 sky130_fd_sc_hd__mux2_1 _3133_ (.A0(_1451_),
    .A1(\tms1x00.RAM[126][2] ),
    .S(_1447_),
    .X(_1452_));
 sky130_fd_sc_hd__clkbuf_1 _3134_ (.A(_1452_),
    .X(_0215_));
 sky130_fd_sc_hd__clkbuf_4 _3135_ (.A(_1132_),
    .X(_1453_));
 sky130_fd_sc_hd__mux2_1 _3136_ (.A0(_1453_),
    .A1(\tms1x00.RAM[126][3] ),
    .S(_1447_),
    .X(_1454_));
 sky130_fd_sc_hd__clkbuf_1 _3137_ (.A(_1454_),
    .X(_0216_));
 sky130_fd_sc_hd__or2_2 _3138_ (.A(_1194_),
    .B(_1242_),
    .X(_1455_));
 sky130_fd_sc_hd__mux2_1 _3139_ (.A0(_1446_),
    .A1(\tms1x00.RAM[1][0] ),
    .S(_1455_),
    .X(_1456_));
 sky130_fd_sc_hd__clkbuf_1 _3140_ (.A(_1456_),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _3141_ (.A0(_1449_),
    .A1(\tms1x00.RAM[1][1] ),
    .S(_1455_),
    .X(_1457_));
 sky130_fd_sc_hd__clkbuf_1 _3142_ (.A(_1457_),
    .X(_0218_));
 sky130_fd_sc_hd__mux2_1 _3143_ (.A0(_1451_),
    .A1(\tms1x00.RAM[1][2] ),
    .S(_1455_),
    .X(_1458_));
 sky130_fd_sc_hd__clkbuf_1 _3144_ (.A(_1458_),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _3145_ (.A0(_1453_),
    .A1(\tms1x00.RAM[1][3] ),
    .S(_1455_),
    .X(_1459_));
 sky130_fd_sc_hd__clkbuf_1 _3146_ (.A(_1459_),
    .X(_0220_));
 sky130_fd_sc_hd__buf_4 _3147_ (.A(_1200_),
    .X(_1460_));
 sky130_fd_sc_hd__nor2_2 _3148_ (.A(_1460_),
    .B(_1257_),
    .Y(_1461_));
 sky130_fd_sc_hd__mux2_1 _3149_ (.A0(\tms1x00.RAM[23][0] ),
    .A1(_1422_),
    .S(_1461_),
    .X(_1462_));
 sky130_fd_sc_hd__clkbuf_1 _3150_ (.A(_1462_),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _3151_ (.A0(\tms1x00.RAM[23][1] ),
    .A1(_1425_),
    .S(_1461_),
    .X(_1463_));
 sky130_fd_sc_hd__clkbuf_1 _3152_ (.A(_1463_),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _3153_ (.A0(\tms1x00.RAM[23][2] ),
    .A1(_1427_),
    .S(_1461_),
    .X(_1464_));
 sky130_fd_sc_hd__clkbuf_1 _3154_ (.A(_1464_),
    .X(_0223_));
 sky130_fd_sc_hd__mux2_1 _3155_ (.A0(\tms1x00.RAM[23][3] ),
    .A1(_1429_),
    .S(_1461_),
    .X(_1465_));
 sky130_fd_sc_hd__clkbuf_1 _3156_ (.A(_1465_),
    .X(_0224_));
 sky130_fd_sc_hd__nor2_2 _3157_ (.A(_1460_),
    .B(_1266_),
    .Y(_1466_));
 sky130_fd_sc_hd__mux2_1 _3158_ (.A0(\tms1x00.RAM[22][0] ),
    .A1(_1422_),
    .S(_1466_),
    .X(_1467_));
 sky130_fd_sc_hd__clkbuf_1 _3159_ (.A(_1467_),
    .X(_0225_));
 sky130_fd_sc_hd__mux2_1 _3160_ (.A0(\tms1x00.RAM[22][1] ),
    .A1(_1425_),
    .S(_1466_),
    .X(_1468_));
 sky130_fd_sc_hd__clkbuf_1 _3161_ (.A(_1468_),
    .X(_0226_));
 sky130_fd_sc_hd__mux2_1 _3162_ (.A0(\tms1x00.RAM[22][2] ),
    .A1(_1427_),
    .S(_1466_),
    .X(_1469_));
 sky130_fd_sc_hd__clkbuf_1 _3163_ (.A(_1469_),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_1 _3164_ (.A0(\tms1x00.RAM[22][3] ),
    .A1(_1429_),
    .S(_1466_),
    .X(_1470_));
 sky130_fd_sc_hd__clkbuf_1 _3165_ (.A(_1470_),
    .X(_0228_));
 sky130_fd_sc_hd__nor2_2 _3166_ (.A(_1180_),
    .B(_1460_),
    .Y(_1471_));
 sky130_fd_sc_hd__mux2_1 _3167_ (.A0(\tms1x00.RAM[21][0] ),
    .A1(_1422_),
    .S(_1471_),
    .X(_1472_));
 sky130_fd_sc_hd__clkbuf_1 _3168_ (.A(_1472_),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_1 _3169_ (.A0(\tms1x00.RAM[21][1] ),
    .A1(_1425_),
    .S(_1471_),
    .X(_1473_));
 sky130_fd_sc_hd__clkbuf_1 _3170_ (.A(_1473_),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_1 _3171_ (.A0(\tms1x00.RAM[21][2] ),
    .A1(_1427_),
    .S(_1471_),
    .X(_1474_));
 sky130_fd_sc_hd__clkbuf_1 _3172_ (.A(_1474_),
    .X(_0231_));
 sky130_fd_sc_hd__mux2_1 _3173_ (.A0(\tms1x00.RAM[21][3] ),
    .A1(_1429_),
    .S(_1471_),
    .X(_1475_));
 sky130_fd_sc_hd__clkbuf_1 _3174_ (.A(_1475_),
    .X(_0232_));
 sky130_fd_sc_hd__nor2_2 _3175_ (.A(_1460_),
    .B(_1304_),
    .Y(_1476_));
 sky130_fd_sc_hd__mux2_1 _3176_ (.A0(\tms1x00.RAM[20][0] ),
    .A1(_1422_),
    .S(_1476_),
    .X(_1477_));
 sky130_fd_sc_hd__clkbuf_1 _3177_ (.A(_1477_),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_1 _3178_ (.A0(\tms1x00.RAM[20][1] ),
    .A1(_1425_),
    .S(_1476_),
    .X(_1478_));
 sky130_fd_sc_hd__clkbuf_1 _3179_ (.A(_1478_),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _3180_ (.A0(\tms1x00.RAM[20][2] ),
    .A1(_1427_),
    .S(_1476_),
    .X(_1479_));
 sky130_fd_sc_hd__clkbuf_1 _3181_ (.A(_1479_),
    .X(_0235_));
 sky130_fd_sc_hd__mux2_1 _3182_ (.A0(\tms1x00.RAM[20][3] ),
    .A1(_1429_),
    .S(_1476_),
    .X(_1480_));
 sky130_fd_sc_hd__clkbuf_1 _3183_ (.A(_1480_),
    .X(_0236_));
 sky130_fd_sc_hd__nor3b_4 _3184_ (.A(_0637_),
    .B(_0639_),
    .C_N(_0635_),
    .Y(_1481_));
 sky130_fd_sc_hd__nand2_2 _3185_ (.A(_1481_),
    .B(_1224_),
    .Y(_1482_));
 sky130_fd_sc_hd__mux2_1 _3186_ (.A0(_1446_),
    .A1(\tms1x00.RAM[28][0] ),
    .S(_1482_),
    .X(_1483_));
 sky130_fd_sc_hd__clkbuf_1 _3187_ (.A(_1483_),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _3188_ (.A0(_1449_),
    .A1(\tms1x00.RAM[28][1] ),
    .S(_1482_),
    .X(_1484_));
 sky130_fd_sc_hd__clkbuf_1 _3189_ (.A(_1484_),
    .X(_0238_));
 sky130_fd_sc_hd__mux2_1 _3190_ (.A0(_1451_),
    .A1(\tms1x00.RAM[28][2] ),
    .S(_1482_),
    .X(_1485_));
 sky130_fd_sc_hd__clkbuf_1 _3191_ (.A(_1485_),
    .X(_0239_));
 sky130_fd_sc_hd__mux2_1 _3192_ (.A0(_1453_),
    .A1(\tms1x00.RAM[28][3] ),
    .S(_1482_),
    .X(_1486_));
 sky130_fd_sc_hd__clkbuf_1 _3193_ (.A(_1486_),
    .X(_0240_));
 sky130_fd_sc_hd__nor2_2 _3194_ (.A(_1153_),
    .B(_1460_),
    .Y(_1487_));
 sky130_fd_sc_hd__mux2_1 _3195_ (.A0(\tms1x00.RAM[27][0] ),
    .A1(_1422_),
    .S(_1487_),
    .X(_1488_));
 sky130_fd_sc_hd__clkbuf_1 _3196_ (.A(_1488_),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_1 _3197_ (.A0(\tms1x00.RAM[27][1] ),
    .A1(_1425_),
    .S(_1487_),
    .X(_1489_));
 sky130_fd_sc_hd__clkbuf_1 _3198_ (.A(_1489_),
    .X(_0242_));
 sky130_fd_sc_hd__mux2_1 _3199_ (.A0(\tms1x00.RAM[27][2] ),
    .A1(_1427_),
    .S(_1487_),
    .X(_1490_));
 sky130_fd_sc_hd__clkbuf_1 _3200_ (.A(_1490_),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _3201_ (.A0(\tms1x00.RAM[27][3] ),
    .A1(_1429_),
    .S(_1487_),
    .X(_1491_));
 sky130_fd_sc_hd__clkbuf_1 _3202_ (.A(_1491_),
    .X(_0244_));
 sky130_fd_sc_hd__nor2_2 _3203_ (.A(_1460_),
    .B(_1236_),
    .Y(_1492_));
 sky130_fd_sc_hd__mux2_1 _3204_ (.A0(\tms1x00.RAM[26][0] ),
    .A1(_1422_),
    .S(_1492_),
    .X(_1493_));
 sky130_fd_sc_hd__clkbuf_1 _3205_ (.A(_1493_),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _3206_ (.A0(\tms1x00.RAM[26][1] ),
    .A1(_1425_),
    .S(_1492_),
    .X(_1494_));
 sky130_fd_sc_hd__clkbuf_1 _3207_ (.A(_1494_),
    .X(_0246_));
 sky130_fd_sc_hd__mux2_1 _3208_ (.A0(\tms1x00.RAM[26][2] ),
    .A1(_1427_),
    .S(_1492_),
    .X(_1495_));
 sky130_fd_sc_hd__clkbuf_1 _3209_ (.A(_1495_),
    .X(_0247_));
 sky130_fd_sc_hd__mux2_1 _3210_ (.A0(\tms1x00.RAM[26][3] ),
    .A1(_1429_),
    .S(_1492_),
    .X(_1496_));
 sky130_fd_sc_hd__clkbuf_1 _3211_ (.A(_1496_),
    .X(_0248_));
 sky130_fd_sc_hd__nor2_2 _3212_ (.A(_1140_),
    .B(_1460_),
    .Y(_1497_));
 sky130_fd_sc_hd__mux2_1 _3213_ (.A0(\tms1x00.RAM[25][0] ),
    .A1(_1422_),
    .S(_1497_),
    .X(_1498_));
 sky130_fd_sc_hd__clkbuf_1 _3214_ (.A(_1498_),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _3215_ (.A0(\tms1x00.RAM[25][1] ),
    .A1(_1425_),
    .S(_1497_),
    .X(_1499_));
 sky130_fd_sc_hd__clkbuf_1 _3216_ (.A(_1499_),
    .X(_0250_));
 sky130_fd_sc_hd__mux2_1 _3217_ (.A0(\tms1x00.RAM[25][2] ),
    .A1(_1427_),
    .S(_1497_),
    .X(_1500_));
 sky130_fd_sc_hd__clkbuf_1 _3218_ (.A(_1500_),
    .X(_0251_));
 sky130_fd_sc_hd__mux2_1 _3219_ (.A0(\tms1x00.RAM[25][3] ),
    .A1(_1429_),
    .S(_1497_),
    .X(_1501_));
 sky130_fd_sc_hd__clkbuf_1 _3220_ (.A(_1501_),
    .X(_0252_));
 sky130_fd_sc_hd__nor2_2 _3221_ (.A(_1460_),
    .B(_1245_),
    .Y(_1502_));
 sky130_fd_sc_hd__mux2_1 _3222_ (.A0(\tms1x00.RAM[24][0] ),
    .A1(_1422_),
    .S(_1502_),
    .X(_1503_));
 sky130_fd_sc_hd__clkbuf_1 _3223_ (.A(_1503_),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _3224_ (.A0(\tms1x00.RAM[24][1] ),
    .A1(_1425_),
    .S(_1502_),
    .X(_1504_));
 sky130_fd_sc_hd__clkbuf_1 _3225_ (.A(_1504_),
    .X(_0254_));
 sky130_fd_sc_hd__mux2_1 _3226_ (.A0(\tms1x00.RAM[24][2] ),
    .A1(_1427_),
    .S(_1502_),
    .X(_1505_));
 sky130_fd_sc_hd__clkbuf_1 _3227_ (.A(_1505_),
    .X(_0255_));
 sky130_fd_sc_hd__mux2_1 _3228_ (.A0(\tms1x00.RAM[24][3] ),
    .A1(_1429_),
    .S(_1502_),
    .X(_1506_));
 sky130_fd_sc_hd__clkbuf_1 _3229_ (.A(_1506_),
    .X(_0256_));
 sky130_fd_sc_hd__or3b_1 _3230_ (.A(\tms1x00.ram_addr_buff[4] ),
    .B(\tms1x00.ram_addr_buff[6] ),
    .C_N(\tms1x00.ram_addr_buff[5] ),
    .X(_1507_));
 sky130_fd_sc_hd__buf_4 _3231_ (.A(_1507_),
    .X(_1508_));
 sky130_fd_sc_hd__or2_2 _3232_ (.A(_1311_),
    .B(_1508_),
    .X(_1509_));
 sky130_fd_sc_hd__mux2_1 _3233_ (.A0(_1446_),
    .A1(\tms1x00.RAM[32][0] ),
    .S(_1509_),
    .X(_1510_));
 sky130_fd_sc_hd__clkbuf_1 _3234_ (.A(_1510_),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _3235_ (.A0(_1449_),
    .A1(\tms1x00.RAM[32][1] ),
    .S(_1509_),
    .X(_1511_));
 sky130_fd_sc_hd__clkbuf_1 _3236_ (.A(_1511_),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_1 _3237_ (.A0(_1451_),
    .A1(\tms1x00.RAM[32][2] ),
    .S(_1509_),
    .X(_1512_));
 sky130_fd_sc_hd__clkbuf_1 _3238_ (.A(_1512_),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _3239_ (.A0(_1453_),
    .A1(\tms1x00.RAM[32][3] ),
    .S(_1509_),
    .X(_1513_));
 sky130_fd_sc_hd__clkbuf_1 _3240_ (.A(_1513_),
    .X(_0260_));
 sky130_fd_sc_hd__nand2_2 _3241_ (.A(_1170_),
    .B(_1481_),
    .Y(_1514_));
 sky130_fd_sc_hd__mux2_1 _3242_ (.A0(_1446_),
    .A1(\tms1x00.RAM[31][0] ),
    .S(_1514_),
    .X(_1515_));
 sky130_fd_sc_hd__clkbuf_1 _3243_ (.A(_1515_),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _3244_ (.A0(_1449_),
    .A1(\tms1x00.RAM[31][1] ),
    .S(_1514_),
    .X(_1516_));
 sky130_fd_sc_hd__clkbuf_1 _3245_ (.A(_1516_),
    .X(_0262_));
 sky130_fd_sc_hd__mux2_1 _3246_ (.A0(_1451_),
    .A1(\tms1x00.RAM[31][2] ),
    .S(_1514_),
    .X(_1517_));
 sky130_fd_sc_hd__clkbuf_1 _3247_ (.A(_1517_),
    .X(_0263_));
 sky130_fd_sc_hd__mux2_1 _3248_ (.A0(_1453_),
    .A1(\tms1x00.RAM[31][3] ),
    .S(_1514_),
    .X(_1518_));
 sky130_fd_sc_hd__clkbuf_1 _3249_ (.A(_1518_),
    .X(_0264_));
 sky130_fd_sc_hd__nand2_2 _3250_ (.A(_1481_),
    .B(_1213_),
    .Y(_1519_));
 sky130_fd_sc_hd__mux2_1 _3251_ (.A0(_1446_),
    .A1(\tms1x00.RAM[30][0] ),
    .S(_1519_),
    .X(_1520_));
 sky130_fd_sc_hd__clkbuf_1 _3252_ (.A(_1520_),
    .X(_0265_));
 sky130_fd_sc_hd__mux2_1 _3253_ (.A0(_1449_),
    .A1(\tms1x00.RAM[30][1] ),
    .S(_1519_),
    .X(_1521_));
 sky130_fd_sc_hd__clkbuf_1 _3254_ (.A(_1521_),
    .X(_0266_));
 sky130_fd_sc_hd__mux2_1 _3255_ (.A0(_1451_),
    .A1(\tms1x00.RAM[30][2] ),
    .S(_1519_),
    .X(_1522_));
 sky130_fd_sc_hd__clkbuf_1 _3256_ (.A(_1522_),
    .X(_0267_));
 sky130_fd_sc_hd__mux2_1 _3257_ (.A0(_1453_),
    .A1(\tms1x00.RAM[30][3] ),
    .S(_1519_),
    .X(_1523_));
 sky130_fd_sc_hd__clkbuf_1 _3258_ (.A(_1523_),
    .X(_0268_));
 sky130_fd_sc_hd__or2_2 _3259_ (.A(_1243_),
    .B(_1320_),
    .X(_1524_));
 sky130_fd_sc_hd__mux2_1 _3260_ (.A0(_1446_),
    .A1(\tms1x00.RAM[2][0] ),
    .S(_1524_),
    .X(_1525_));
 sky130_fd_sc_hd__clkbuf_1 _3261_ (.A(_1525_),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _3262_ (.A0(_1449_),
    .A1(\tms1x00.RAM[2][1] ),
    .S(_1524_),
    .X(_1526_));
 sky130_fd_sc_hd__clkbuf_1 _3263_ (.A(_1526_),
    .X(_0270_));
 sky130_fd_sc_hd__mux2_1 _3264_ (.A0(_1451_),
    .A1(\tms1x00.RAM[2][2] ),
    .S(_1524_),
    .X(_1527_));
 sky130_fd_sc_hd__clkbuf_1 _3265_ (.A(_1527_),
    .X(_0271_));
 sky130_fd_sc_hd__mux2_1 _3266_ (.A0(_1453_),
    .A1(\tms1x00.RAM[2][3] ),
    .S(_1524_),
    .X(_1528_));
 sky130_fd_sc_hd__clkbuf_1 _3267_ (.A(_1528_),
    .X(_0272_));
 sky130_fd_sc_hd__nor2_2 _3268_ (.A(_1304_),
    .B(_1508_),
    .Y(_1529_));
 sky130_fd_sc_hd__mux2_1 _3269_ (.A0(\tms1x00.RAM[36][0] ),
    .A1(_1422_),
    .S(_1529_),
    .X(_1530_));
 sky130_fd_sc_hd__clkbuf_1 _3270_ (.A(_1530_),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _3271_ (.A0(\tms1x00.RAM[36][1] ),
    .A1(_1425_),
    .S(_1529_),
    .X(_1531_));
 sky130_fd_sc_hd__clkbuf_1 _3272_ (.A(_1531_),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_1 _3273_ (.A0(\tms1x00.RAM[36][2] ),
    .A1(_1427_),
    .S(_1529_),
    .X(_1532_));
 sky130_fd_sc_hd__clkbuf_1 _3274_ (.A(_1532_),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_1 _3275_ (.A0(\tms1x00.RAM[36][3] ),
    .A1(_1429_),
    .S(_1529_),
    .X(_1533_));
 sky130_fd_sc_hd__clkbuf_1 _3276_ (.A(_1533_),
    .X(_0276_));
 sky130_fd_sc_hd__or2_2 _3277_ (.A(_0833_),
    .B(_1508_),
    .X(_1534_));
 sky130_fd_sc_hd__mux2_1 _3278_ (.A0(_1446_),
    .A1(\tms1x00.RAM[35][0] ),
    .S(_1534_),
    .X(_1535_));
 sky130_fd_sc_hd__clkbuf_1 _3279_ (.A(_1535_),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_1 _3280_ (.A0(_1449_),
    .A1(\tms1x00.RAM[35][1] ),
    .S(_1534_),
    .X(_1536_));
 sky130_fd_sc_hd__clkbuf_1 _3281_ (.A(_1536_),
    .X(_0278_));
 sky130_fd_sc_hd__mux2_1 _3282_ (.A0(_1451_),
    .A1(\tms1x00.RAM[35][2] ),
    .S(_1534_),
    .X(_1537_));
 sky130_fd_sc_hd__clkbuf_1 _3283_ (.A(_1537_),
    .X(_0279_));
 sky130_fd_sc_hd__mux2_1 _3284_ (.A0(_1453_),
    .A1(\tms1x00.RAM[35][3] ),
    .S(_1534_),
    .X(_1538_));
 sky130_fd_sc_hd__clkbuf_1 _3285_ (.A(_1538_),
    .X(_0280_));
 sky130_fd_sc_hd__or2_2 _3286_ (.A(_1320_),
    .B(_1507_),
    .X(_1539_));
 sky130_fd_sc_hd__mux2_1 _3287_ (.A0(_1446_),
    .A1(\tms1x00.RAM[34][0] ),
    .S(_1539_),
    .X(_1540_));
 sky130_fd_sc_hd__clkbuf_1 _3288_ (.A(_1540_),
    .X(_0281_));
 sky130_fd_sc_hd__mux2_1 _3289_ (.A0(_1449_),
    .A1(\tms1x00.RAM[34][1] ),
    .S(_1539_),
    .X(_1541_));
 sky130_fd_sc_hd__clkbuf_1 _3290_ (.A(_1541_),
    .X(_0282_));
 sky130_fd_sc_hd__mux2_1 _3291_ (.A0(_1451_),
    .A1(\tms1x00.RAM[34][2] ),
    .S(_1539_),
    .X(_1542_));
 sky130_fd_sc_hd__clkbuf_1 _3292_ (.A(_1542_),
    .X(_0283_));
 sky130_fd_sc_hd__mux2_1 _3293_ (.A0(_1453_),
    .A1(\tms1x00.RAM[34][3] ),
    .S(_1539_),
    .X(_1543_));
 sky130_fd_sc_hd__clkbuf_1 _3294_ (.A(_1543_),
    .X(_0284_));
 sky130_fd_sc_hd__or2_2 _3295_ (.A(_1194_),
    .B(_1507_),
    .X(_1544_));
 sky130_fd_sc_hd__mux2_1 _3296_ (.A0(_1446_),
    .A1(\tms1x00.RAM[33][0] ),
    .S(_1544_),
    .X(_1545_));
 sky130_fd_sc_hd__clkbuf_1 _3297_ (.A(_1545_),
    .X(_0285_));
 sky130_fd_sc_hd__mux2_1 _3298_ (.A0(_1449_),
    .A1(\tms1x00.RAM[33][1] ),
    .S(_1544_),
    .X(_1546_));
 sky130_fd_sc_hd__clkbuf_1 _3299_ (.A(_1546_),
    .X(_0286_));
 sky130_fd_sc_hd__mux2_1 _3300_ (.A0(_1451_),
    .A1(\tms1x00.RAM[33][2] ),
    .S(_1544_),
    .X(_1547_));
 sky130_fd_sc_hd__clkbuf_1 _3301_ (.A(_1547_),
    .X(_0287_));
 sky130_fd_sc_hd__mux2_1 _3302_ (.A0(_1453_),
    .A1(\tms1x00.RAM[33][3] ),
    .S(_1544_),
    .X(_1548_));
 sky130_fd_sc_hd__clkbuf_1 _3303_ (.A(_1548_),
    .X(_0288_));
 sky130_fd_sc_hd__buf_2 _3304_ (.A(_0826_),
    .X(_1549_));
 sky130_fd_sc_hd__nor2_2 _3305_ (.A(_1140_),
    .B(_1508_),
    .Y(_1550_));
 sky130_fd_sc_hd__mux2_1 _3306_ (.A0(\tms1x00.RAM[41][0] ),
    .A1(_1549_),
    .S(_1550_),
    .X(_1551_));
 sky130_fd_sc_hd__clkbuf_1 _3307_ (.A(_1551_),
    .X(_0289_));
 sky130_fd_sc_hd__buf_2 _3308_ (.A(_0934_),
    .X(_1552_));
 sky130_fd_sc_hd__mux2_1 _3309_ (.A0(\tms1x00.RAM[41][1] ),
    .A1(_1552_),
    .S(_1550_),
    .X(_1553_));
 sky130_fd_sc_hd__clkbuf_1 _3310_ (.A(_1553_),
    .X(_0290_));
 sky130_fd_sc_hd__buf_2 _3311_ (.A(_1034_),
    .X(_1554_));
 sky130_fd_sc_hd__mux2_1 _3312_ (.A0(\tms1x00.RAM[41][2] ),
    .A1(_1554_),
    .S(_1550_),
    .X(_1555_));
 sky130_fd_sc_hd__clkbuf_1 _3313_ (.A(_1555_),
    .X(_0291_));
 sky130_fd_sc_hd__buf_2 _3314_ (.A(_1132_),
    .X(_1556_));
 sky130_fd_sc_hd__mux2_1 _3315_ (.A0(\tms1x00.RAM[41][3] ),
    .A1(_1556_),
    .S(_1550_),
    .X(_1557_));
 sky130_fd_sc_hd__clkbuf_1 _3316_ (.A(_1557_),
    .X(_0292_));
 sky130_fd_sc_hd__nor2_2 _3317_ (.A(_1245_),
    .B(_1508_),
    .Y(_1558_));
 sky130_fd_sc_hd__mux2_1 _3318_ (.A0(\tms1x00.RAM[40][0] ),
    .A1(_1549_),
    .S(_1558_),
    .X(_1559_));
 sky130_fd_sc_hd__clkbuf_1 _3319_ (.A(_1559_),
    .X(_0293_));
 sky130_fd_sc_hd__mux2_1 _3320_ (.A0(\tms1x00.RAM[40][1] ),
    .A1(_1552_),
    .S(_1558_),
    .X(_1560_));
 sky130_fd_sc_hd__clkbuf_1 _3321_ (.A(_1560_),
    .X(_0294_));
 sky130_fd_sc_hd__mux2_1 _3322_ (.A0(\tms1x00.RAM[40][2] ),
    .A1(_1554_),
    .S(_1558_),
    .X(_1561_));
 sky130_fd_sc_hd__clkbuf_1 _3323_ (.A(_1561_),
    .X(_0295_));
 sky130_fd_sc_hd__mux2_1 _3324_ (.A0(\tms1x00.RAM[40][3] ),
    .A1(_1556_),
    .S(_1558_),
    .X(_1562_));
 sky130_fd_sc_hd__clkbuf_1 _3325_ (.A(_1562_),
    .X(_0296_));
 sky130_fd_sc_hd__buf_2 _3326_ (.A(_0826_),
    .X(_1563_));
 sky130_fd_sc_hd__or2_2 _3327_ (.A(_0833_),
    .B(_1242_),
    .X(_1564_));
 sky130_fd_sc_hd__mux2_1 _3328_ (.A0(_1563_),
    .A1(\tms1x00.RAM[3][0] ),
    .S(_1564_),
    .X(_1565_));
 sky130_fd_sc_hd__clkbuf_1 _3329_ (.A(_1565_),
    .X(_0297_));
 sky130_fd_sc_hd__buf_2 _3330_ (.A(_0934_),
    .X(_1566_));
 sky130_fd_sc_hd__mux2_1 _3331_ (.A0(_1566_),
    .A1(\tms1x00.RAM[3][1] ),
    .S(_1564_),
    .X(_1567_));
 sky130_fd_sc_hd__clkbuf_1 _3332_ (.A(_1567_),
    .X(_0298_));
 sky130_fd_sc_hd__buf_2 _3333_ (.A(_1034_),
    .X(_1568_));
 sky130_fd_sc_hd__mux2_1 _3334_ (.A0(_1568_),
    .A1(\tms1x00.RAM[3][2] ),
    .S(_1564_),
    .X(_1569_));
 sky130_fd_sc_hd__clkbuf_1 _3335_ (.A(_1569_),
    .X(_0299_));
 sky130_fd_sc_hd__buf_2 _3336_ (.A(_1132_),
    .X(_1570_));
 sky130_fd_sc_hd__mux2_1 _3337_ (.A0(_1570_),
    .A1(\tms1x00.RAM[3][3] ),
    .S(_1564_),
    .X(_1571_));
 sky130_fd_sc_hd__clkbuf_1 _3338_ (.A(_1571_),
    .X(_0300_));
 sky130_fd_sc_hd__nor2_2 _3339_ (.A(_1266_),
    .B(_1508_),
    .Y(_1572_));
 sky130_fd_sc_hd__mux2_1 _3340_ (.A0(\tms1x00.RAM[38][0] ),
    .A1(_1549_),
    .S(_1572_),
    .X(_1573_));
 sky130_fd_sc_hd__clkbuf_1 _3341_ (.A(_1573_),
    .X(_0301_));
 sky130_fd_sc_hd__mux2_1 _3342_ (.A0(\tms1x00.RAM[38][1] ),
    .A1(_1552_),
    .S(_1572_),
    .X(_1574_));
 sky130_fd_sc_hd__clkbuf_1 _3343_ (.A(_1574_),
    .X(_0302_));
 sky130_fd_sc_hd__mux2_1 _3344_ (.A0(\tms1x00.RAM[38][2] ),
    .A1(_1554_),
    .S(_1572_),
    .X(_1575_));
 sky130_fd_sc_hd__clkbuf_1 _3345_ (.A(_1575_),
    .X(_0303_));
 sky130_fd_sc_hd__mux2_1 _3346_ (.A0(\tms1x00.RAM[38][3] ),
    .A1(_1556_),
    .S(_1572_),
    .X(_1576_));
 sky130_fd_sc_hd__clkbuf_1 _3347_ (.A(_1576_),
    .X(_0304_));
 sky130_fd_sc_hd__nor2_2 _3348_ (.A(_1180_),
    .B(_1508_),
    .Y(_1577_));
 sky130_fd_sc_hd__mux2_1 _3349_ (.A0(\tms1x00.RAM[37][0] ),
    .A1(_1549_),
    .S(_1577_),
    .X(_1578_));
 sky130_fd_sc_hd__clkbuf_1 _3350_ (.A(_1578_),
    .X(_0305_));
 sky130_fd_sc_hd__mux2_1 _3351_ (.A0(\tms1x00.RAM[37][1] ),
    .A1(_1552_),
    .S(_1577_),
    .X(_1579_));
 sky130_fd_sc_hd__clkbuf_1 _3352_ (.A(_1579_),
    .X(_0306_));
 sky130_fd_sc_hd__mux2_1 _3353_ (.A0(\tms1x00.RAM[37][2] ),
    .A1(_1554_),
    .S(_1577_),
    .X(_1580_));
 sky130_fd_sc_hd__clkbuf_1 _3354_ (.A(_1580_),
    .X(_0307_));
 sky130_fd_sc_hd__mux2_1 _3355_ (.A0(\tms1x00.RAM[37][3] ),
    .A1(_1556_),
    .S(_1577_),
    .X(_1581_));
 sky130_fd_sc_hd__clkbuf_1 _3356_ (.A(_1581_),
    .X(_0308_));
 sky130_fd_sc_hd__nor3b_2 _3357_ (.A(_0635_),
    .B(_0639_),
    .C_N(_0637_),
    .Y(_1582_));
 sky130_fd_sc_hd__nand2_2 _3358_ (.A(_1162_),
    .B(_1582_),
    .Y(_1583_));
 sky130_fd_sc_hd__mux2_1 _3359_ (.A0(_1563_),
    .A1(\tms1x00.RAM[45][0] ),
    .S(_1583_),
    .X(_1584_));
 sky130_fd_sc_hd__clkbuf_1 _3360_ (.A(_1584_),
    .X(_0309_));
 sky130_fd_sc_hd__mux2_1 _3361_ (.A0(_1566_),
    .A1(\tms1x00.RAM[45][1] ),
    .S(_1583_),
    .X(_1585_));
 sky130_fd_sc_hd__clkbuf_1 _3362_ (.A(_1585_),
    .X(_0310_));
 sky130_fd_sc_hd__mux2_1 _3363_ (.A0(_1568_),
    .A1(\tms1x00.RAM[45][2] ),
    .S(_1583_),
    .X(_1586_));
 sky130_fd_sc_hd__clkbuf_1 _3364_ (.A(_1586_),
    .X(_0311_));
 sky130_fd_sc_hd__mux2_1 _3365_ (.A0(_1570_),
    .A1(\tms1x00.RAM[45][3] ),
    .S(_1583_),
    .X(_1587_));
 sky130_fd_sc_hd__clkbuf_1 _3366_ (.A(_1587_),
    .X(_0312_));
 sky130_fd_sc_hd__nand2_2 _3367_ (.A(_1224_),
    .B(_1582_),
    .Y(_1588_));
 sky130_fd_sc_hd__mux2_1 _3368_ (.A0(_1563_),
    .A1(\tms1x00.RAM[44][0] ),
    .S(_1588_),
    .X(_1589_));
 sky130_fd_sc_hd__clkbuf_1 _3369_ (.A(_1589_),
    .X(_0313_));
 sky130_fd_sc_hd__mux2_1 _3370_ (.A0(_1566_),
    .A1(\tms1x00.RAM[44][1] ),
    .S(_1588_),
    .X(_1590_));
 sky130_fd_sc_hd__clkbuf_1 _3371_ (.A(_1590_),
    .X(_0314_));
 sky130_fd_sc_hd__mux2_1 _3372_ (.A0(_1568_),
    .A1(\tms1x00.RAM[44][2] ),
    .S(_1588_),
    .X(_1591_));
 sky130_fd_sc_hd__clkbuf_1 _3373_ (.A(_1591_),
    .X(_0315_));
 sky130_fd_sc_hd__mux2_1 _3374_ (.A0(_1570_),
    .A1(\tms1x00.RAM[44][3] ),
    .S(_1588_),
    .X(_1592_));
 sky130_fd_sc_hd__clkbuf_1 _3375_ (.A(_1592_),
    .X(_0316_));
 sky130_fd_sc_hd__nor2_2 _3376_ (.A(_1153_),
    .B(_1508_),
    .Y(_1593_));
 sky130_fd_sc_hd__mux2_1 _3377_ (.A0(\tms1x00.RAM[43][0] ),
    .A1(_1549_),
    .S(_1593_),
    .X(_1594_));
 sky130_fd_sc_hd__clkbuf_1 _3378_ (.A(_1594_),
    .X(_0317_));
 sky130_fd_sc_hd__mux2_1 _3379_ (.A0(\tms1x00.RAM[43][1] ),
    .A1(_1552_),
    .S(_1593_),
    .X(_1595_));
 sky130_fd_sc_hd__clkbuf_1 _3380_ (.A(_1595_),
    .X(_0318_));
 sky130_fd_sc_hd__mux2_1 _3381_ (.A0(\tms1x00.RAM[43][2] ),
    .A1(_1554_),
    .S(_1593_),
    .X(_1596_));
 sky130_fd_sc_hd__clkbuf_1 _3382_ (.A(_1596_),
    .X(_0319_));
 sky130_fd_sc_hd__mux2_1 _3383_ (.A0(\tms1x00.RAM[43][3] ),
    .A1(_1556_),
    .S(_1593_),
    .X(_1597_));
 sky130_fd_sc_hd__clkbuf_1 _3384_ (.A(_1597_),
    .X(_0320_));
 sky130_fd_sc_hd__nor2_2 _3385_ (.A(_1236_),
    .B(_1508_),
    .Y(_1598_));
 sky130_fd_sc_hd__mux2_1 _3386_ (.A0(\tms1x00.RAM[42][0] ),
    .A1(_1549_),
    .S(_1598_),
    .X(_1599_));
 sky130_fd_sc_hd__clkbuf_1 _3387_ (.A(_1599_),
    .X(_0321_));
 sky130_fd_sc_hd__mux2_1 _3388_ (.A0(\tms1x00.RAM[42][1] ),
    .A1(_1552_),
    .S(_1598_),
    .X(_1600_));
 sky130_fd_sc_hd__clkbuf_1 _3389_ (.A(_1600_),
    .X(_0322_));
 sky130_fd_sc_hd__mux2_1 _3390_ (.A0(\tms1x00.RAM[42][2] ),
    .A1(_1554_),
    .S(_1598_),
    .X(_1601_));
 sky130_fd_sc_hd__clkbuf_1 _3391_ (.A(_1601_),
    .X(_0323_));
 sky130_fd_sc_hd__mux2_1 _3392_ (.A0(\tms1x00.RAM[42][3] ),
    .A1(_1556_),
    .S(_1598_),
    .X(_1602_));
 sky130_fd_sc_hd__clkbuf_1 _3393_ (.A(_1602_),
    .X(_0324_));
 sky130_fd_sc_hd__or2_2 _3394_ (.A(_1151_),
    .B(_1320_),
    .X(_1603_));
 sky130_fd_sc_hd__mux2_1 _3395_ (.A0(_1563_),
    .A1(\tms1x00.RAM[50][0] ),
    .S(_1603_),
    .X(_1604_));
 sky130_fd_sc_hd__clkbuf_1 _3396_ (.A(_1604_),
    .X(_0325_));
 sky130_fd_sc_hd__mux2_1 _3397_ (.A0(_1566_),
    .A1(\tms1x00.RAM[50][1] ),
    .S(_1603_),
    .X(_1605_));
 sky130_fd_sc_hd__clkbuf_1 _3398_ (.A(_1605_),
    .X(_0326_));
 sky130_fd_sc_hd__mux2_1 _3399_ (.A0(_1568_),
    .A1(\tms1x00.RAM[50][2] ),
    .S(_1603_),
    .X(_1606_));
 sky130_fd_sc_hd__clkbuf_1 _3400_ (.A(_1606_),
    .X(_0327_));
 sky130_fd_sc_hd__mux2_1 _3401_ (.A0(_1570_),
    .A1(\tms1x00.RAM[50][3] ),
    .S(_1603_),
    .X(_1607_));
 sky130_fd_sc_hd__clkbuf_1 _3402_ (.A(_1607_),
    .X(_0328_));
 sky130_fd_sc_hd__nor2_2 _3403_ (.A(_1243_),
    .B(_1304_),
    .Y(_1608_));
 sky130_fd_sc_hd__mux2_1 _3404_ (.A0(\tms1x00.RAM[4][0] ),
    .A1(_1549_),
    .S(_1608_),
    .X(_1609_));
 sky130_fd_sc_hd__clkbuf_1 _3405_ (.A(_1609_),
    .X(_0329_));
 sky130_fd_sc_hd__mux2_1 _3406_ (.A0(\tms1x00.RAM[4][1] ),
    .A1(_1552_),
    .S(_1608_),
    .X(_1610_));
 sky130_fd_sc_hd__clkbuf_1 _3407_ (.A(_1610_),
    .X(_0330_));
 sky130_fd_sc_hd__mux2_1 _3408_ (.A0(\tms1x00.RAM[4][2] ),
    .A1(_1554_),
    .S(_1608_),
    .X(_1611_));
 sky130_fd_sc_hd__clkbuf_1 _3409_ (.A(_1611_),
    .X(_0331_));
 sky130_fd_sc_hd__mux2_1 _3410_ (.A0(\tms1x00.RAM[4][3] ),
    .A1(_1556_),
    .S(_1608_),
    .X(_1612_));
 sky130_fd_sc_hd__clkbuf_1 _3411_ (.A(_1612_),
    .X(_0332_));
 sky130_fd_sc_hd__or2_2 _3412_ (.A(_1150_),
    .B(_1311_),
    .X(_1613_));
 sky130_fd_sc_hd__mux2_1 _3413_ (.A0(_1563_),
    .A1(\tms1x00.RAM[48][0] ),
    .S(_1613_),
    .X(_1614_));
 sky130_fd_sc_hd__clkbuf_1 _3414_ (.A(_1614_),
    .X(_0333_));
 sky130_fd_sc_hd__mux2_1 _3415_ (.A0(_1566_),
    .A1(\tms1x00.RAM[48][1] ),
    .S(_1613_),
    .X(_1615_));
 sky130_fd_sc_hd__clkbuf_1 _3416_ (.A(_1615_),
    .X(_0334_));
 sky130_fd_sc_hd__mux2_1 _3417_ (.A0(_1568_),
    .A1(\tms1x00.RAM[48][2] ),
    .S(_1613_),
    .X(_1616_));
 sky130_fd_sc_hd__clkbuf_1 _3418_ (.A(_1616_),
    .X(_0335_));
 sky130_fd_sc_hd__mux2_1 _3419_ (.A0(_1570_),
    .A1(\tms1x00.RAM[48][3] ),
    .S(_1613_),
    .X(_1617_));
 sky130_fd_sc_hd__clkbuf_1 _3420_ (.A(_1617_),
    .X(_0336_));
 sky130_fd_sc_hd__nand2_2 _3421_ (.A(_1170_),
    .B(_1582_),
    .Y(_1618_));
 sky130_fd_sc_hd__mux2_1 _3422_ (.A0(_1563_),
    .A1(\tms1x00.RAM[47][0] ),
    .S(_1618_),
    .X(_1619_));
 sky130_fd_sc_hd__clkbuf_1 _3423_ (.A(_1619_),
    .X(_0337_));
 sky130_fd_sc_hd__mux2_1 _3424_ (.A0(_1566_),
    .A1(\tms1x00.RAM[47][1] ),
    .S(_1618_),
    .X(_1620_));
 sky130_fd_sc_hd__clkbuf_1 _3425_ (.A(_1620_),
    .X(_0338_));
 sky130_fd_sc_hd__mux2_1 _3426_ (.A0(_1568_),
    .A1(\tms1x00.RAM[47][2] ),
    .S(_1618_),
    .X(_1621_));
 sky130_fd_sc_hd__clkbuf_1 _3427_ (.A(_1621_),
    .X(_0339_));
 sky130_fd_sc_hd__mux2_1 _3428_ (.A0(_1570_),
    .A1(\tms1x00.RAM[47][3] ),
    .S(_1618_),
    .X(_1622_));
 sky130_fd_sc_hd__clkbuf_1 _3429_ (.A(_1622_),
    .X(_0340_));
 sky130_fd_sc_hd__nand2_2 _3430_ (.A(_1213_),
    .B(_1582_),
    .Y(_1623_));
 sky130_fd_sc_hd__mux2_1 _3431_ (.A0(_1563_),
    .A1(\tms1x00.RAM[46][0] ),
    .S(_1623_),
    .X(_1624_));
 sky130_fd_sc_hd__clkbuf_1 _3432_ (.A(_1624_),
    .X(_0341_));
 sky130_fd_sc_hd__mux2_1 _3433_ (.A0(_1566_),
    .A1(\tms1x00.RAM[46][1] ),
    .S(_1623_),
    .X(_1625_));
 sky130_fd_sc_hd__clkbuf_1 _3434_ (.A(_1625_),
    .X(_0342_));
 sky130_fd_sc_hd__mux2_1 _3435_ (.A0(_1568_),
    .A1(\tms1x00.RAM[46][2] ),
    .S(_1623_),
    .X(_1626_));
 sky130_fd_sc_hd__clkbuf_1 _3436_ (.A(_1626_),
    .X(_0343_));
 sky130_fd_sc_hd__mux2_1 _3437_ (.A0(_1570_),
    .A1(\tms1x00.RAM[46][3] ),
    .S(_1623_),
    .X(_1627_));
 sky130_fd_sc_hd__clkbuf_1 _3438_ (.A(_1627_),
    .X(_0344_));
 sky130_fd_sc_hd__nor2_2 _3439_ (.A(_1151_),
    .B(_1266_),
    .Y(_1628_));
 sky130_fd_sc_hd__mux2_1 _3440_ (.A0(\tms1x00.RAM[54][0] ),
    .A1(_1549_),
    .S(_1628_),
    .X(_1629_));
 sky130_fd_sc_hd__clkbuf_1 _3441_ (.A(_1629_),
    .X(_0345_));
 sky130_fd_sc_hd__mux2_1 _3442_ (.A0(\tms1x00.RAM[54][1] ),
    .A1(_1552_),
    .S(_1628_),
    .X(_1630_));
 sky130_fd_sc_hd__clkbuf_1 _3443_ (.A(_1630_),
    .X(_0346_));
 sky130_fd_sc_hd__mux2_1 _3444_ (.A0(\tms1x00.RAM[54][2] ),
    .A1(_1554_),
    .S(_1628_),
    .X(_1631_));
 sky130_fd_sc_hd__clkbuf_1 _3445_ (.A(_1631_),
    .X(_0347_));
 sky130_fd_sc_hd__mux2_1 _3446_ (.A0(\tms1x00.RAM[54][3] ),
    .A1(_1556_),
    .S(_1628_),
    .X(_1632_));
 sky130_fd_sc_hd__clkbuf_1 _3447_ (.A(_1632_),
    .X(_0348_));
 sky130_fd_sc_hd__nor2_2 _3448_ (.A(_1151_),
    .B(_1180_),
    .Y(_1633_));
 sky130_fd_sc_hd__mux2_1 _3449_ (.A0(\tms1x00.RAM[53][0] ),
    .A1(_1549_),
    .S(_1633_),
    .X(_1634_));
 sky130_fd_sc_hd__clkbuf_1 _3450_ (.A(_1634_),
    .X(_0349_));
 sky130_fd_sc_hd__mux2_1 _3451_ (.A0(\tms1x00.RAM[53][1] ),
    .A1(_1552_),
    .S(_1633_),
    .X(_1635_));
 sky130_fd_sc_hd__clkbuf_1 _3452_ (.A(_1635_),
    .X(_0350_));
 sky130_fd_sc_hd__mux2_1 _3453_ (.A0(\tms1x00.RAM[53][2] ),
    .A1(_1554_),
    .S(_1633_),
    .X(_1636_));
 sky130_fd_sc_hd__clkbuf_1 _3454_ (.A(_1636_),
    .X(_0351_));
 sky130_fd_sc_hd__mux2_1 _3455_ (.A0(\tms1x00.RAM[53][3] ),
    .A1(_1556_),
    .S(_1633_),
    .X(_1637_));
 sky130_fd_sc_hd__clkbuf_1 _3456_ (.A(_1637_),
    .X(_0352_));
 sky130_fd_sc_hd__nor2_2 _3457_ (.A(_1151_),
    .B(_1304_),
    .Y(_1638_));
 sky130_fd_sc_hd__mux2_1 _3458_ (.A0(\tms1x00.RAM[52][0] ),
    .A1(_1549_),
    .S(_1638_),
    .X(_1639_));
 sky130_fd_sc_hd__clkbuf_1 _3459_ (.A(_1639_),
    .X(_0353_));
 sky130_fd_sc_hd__mux2_1 _3460_ (.A0(\tms1x00.RAM[52][1] ),
    .A1(_1552_),
    .S(_1638_),
    .X(_1640_));
 sky130_fd_sc_hd__clkbuf_1 _3461_ (.A(_1640_),
    .X(_0354_));
 sky130_fd_sc_hd__mux2_1 _3462_ (.A0(\tms1x00.RAM[52][2] ),
    .A1(_1554_),
    .S(_1638_),
    .X(_1641_));
 sky130_fd_sc_hd__clkbuf_1 _3463_ (.A(_1641_),
    .X(_0355_));
 sky130_fd_sc_hd__mux2_1 _3464_ (.A0(\tms1x00.RAM[52][3] ),
    .A1(_1556_),
    .S(_1638_),
    .X(_1642_));
 sky130_fd_sc_hd__clkbuf_1 _3465_ (.A(_1642_),
    .X(_0356_));
 sky130_fd_sc_hd__or2_2 _3466_ (.A(_0833_),
    .B(_1150_),
    .X(_1643_));
 sky130_fd_sc_hd__mux2_1 _3467_ (.A0(_1563_),
    .A1(\tms1x00.RAM[51][0] ),
    .S(_1643_),
    .X(_1644_));
 sky130_fd_sc_hd__clkbuf_1 _3468_ (.A(_1644_),
    .X(_0357_));
 sky130_fd_sc_hd__mux2_1 _3469_ (.A0(_1566_),
    .A1(\tms1x00.RAM[51][1] ),
    .S(_1643_),
    .X(_1645_));
 sky130_fd_sc_hd__clkbuf_1 _3470_ (.A(_1645_),
    .X(_0358_));
 sky130_fd_sc_hd__mux2_1 _3471_ (.A0(_1568_),
    .A1(\tms1x00.RAM[51][2] ),
    .S(_1643_),
    .X(_1646_));
 sky130_fd_sc_hd__clkbuf_1 _3472_ (.A(_1646_),
    .X(_0359_));
 sky130_fd_sc_hd__mux2_1 _3473_ (.A0(_1570_),
    .A1(\tms1x00.RAM[51][3] ),
    .S(_1643_),
    .X(_1647_));
 sky130_fd_sc_hd__clkbuf_1 _3474_ (.A(_1647_),
    .X(_0360_));
 sky130_fd_sc_hd__clkbuf_4 _3475_ (.A(_0826_),
    .X(_1648_));
 sky130_fd_sc_hd__nor2_2 _3476_ (.A(_1151_),
    .B(_1236_),
    .Y(_1649_));
 sky130_fd_sc_hd__mux2_1 _3477_ (.A0(\tms1x00.RAM[58][0] ),
    .A1(_1648_),
    .S(_1649_),
    .X(_1650_));
 sky130_fd_sc_hd__clkbuf_1 _3478_ (.A(_1650_),
    .X(_0361_));
 sky130_fd_sc_hd__clkbuf_4 _3479_ (.A(_0934_),
    .X(_1651_));
 sky130_fd_sc_hd__mux2_1 _3480_ (.A0(\tms1x00.RAM[58][1] ),
    .A1(_1651_),
    .S(_1649_),
    .X(_1652_));
 sky130_fd_sc_hd__clkbuf_1 _3481_ (.A(_1652_),
    .X(_0362_));
 sky130_fd_sc_hd__clkbuf_4 _3482_ (.A(_1034_),
    .X(_1653_));
 sky130_fd_sc_hd__mux2_1 _3483_ (.A0(\tms1x00.RAM[58][2] ),
    .A1(_1653_),
    .S(_1649_),
    .X(_1654_));
 sky130_fd_sc_hd__clkbuf_1 _3484_ (.A(_1654_),
    .X(_0363_));
 sky130_fd_sc_hd__clkbuf_4 _3485_ (.A(_1132_),
    .X(_1655_));
 sky130_fd_sc_hd__mux2_1 _3486_ (.A0(\tms1x00.RAM[58][3] ),
    .A1(_1655_),
    .S(_1649_),
    .X(_1656_));
 sky130_fd_sc_hd__clkbuf_1 _3487_ (.A(_1656_),
    .X(_0364_));
 sky130_fd_sc_hd__nor2_2 _3488_ (.A(_1140_),
    .B(_1151_),
    .Y(_1657_));
 sky130_fd_sc_hd__mux2_1 _3489_ (.A0(\tms1x00.RAM[57][0] ),
    .A1(_1648_),
    .S(_1657_),
    .X(_1658_));
 sky130_fd_sc_hd__clkbuf_1 _3490_ (.A(_1658_),
    .X(_0365_));
 sky130_fd_sc_hd__mux2_1 _3491_ (.A0(\tms1x00.RAM[57][1] ),
    .A1(_1651_),
    .S(_1657_),
    .X(_1659_));
 sky130_fd_sc_hd__clkbuf_1 _3492_ (.A(_1659_),
    .X(_0366_));
 sky130_fd_sc_hd__mux2_1 _3493_ (.A0(\tms1x00.RAM[57][2] ),
    .A1(_1653_),
    .S(_1657_),
    .X(_1660_));
 sky130_fd_sc_hd__clkbuf_1 _3494_ (.A(_1660_),
    .X(_0367_));
 sky130_fd_sc_hd__mux2_1 _3495_ (.A0(\tms1x00.RAM[57][3] ),
    .A1(_1655_),
    .S(_1657_),
    .X(_1661_));
 sky130_fd_sc_hd__clkbuf_1 _3496_ (.A(_1661_),
    .X(_0368_));
 sky130_fd_sc_hd__nor2_2 _3497_ (.A(_1151_),
    .B(_1245_),
    .Y(_1662_));
 sky130_fd_sc_hd__mux2_1 _3498_ (.A0(\tms1x00.RAM[56][0] ),
    .A1(_1648_),
    .S(_1662_),
    .X(_1663_));
 sky130_fd_sc_hd__clkbuf_1 _3499_ (.A(_1663_),
    .X(_0369_));
 sky130_fd_sc_hd__mux2_1 _3500_ (.A0(\tms1x00.RAM[56][1] ),
    .A1(_1651_),
    .S(_1662_),
    .X(_1664_));
 sky130_fd_sc_hd__clkbuf_1 _3501_ (.A(_1664_),
    .X(_0370_));
 sky130_fd_sc_hd__mux2_1 _3502_ (.A0(\tms1x00.RAM[56][2] ),
    .A1(_1653_),
    .S(_1662_),
    .X(_1665_));
 sky130_fd_sc_hd__clkbuf_1 _3503_ (.A(_1665_),
    .X(_0371_));
 sky130_fd_sc_hd__mux2_1 _3504_ (.A0(\tms1x00.RAM[56][3] ),
    .A1(_1655_),
    .S(_1662_),
    .X(_1666_));
 sky130_fd_sc_hd__clkbuf_1 _3505_ (.A(_1666_),
    .X(_0372_));
 sky130_fd_sc_hd__nor2_2 _3506_ (.A(_1151_),
    .B(_1257_),
    .Y(_1667_));
 sky130_fd_sc_hd__mux2_1 _3507_ (.A0(\tms1x00.RAM[55][0] ),
    .A1(_1648_),
    .S(_1667_),
    .X(_1668_));
 sky130_fd_sc_hd__clkbuf_1 _3508_ (.A(_1668_),
    .X(_0373_));
 sky130_fd_sc_hd__mux2_1 _3509_ (.A0(\tms1x00.RAM[55][1] ),
    .A1(_1651_),
    .S(_1667_),
    .X(_1669_));
 sky130_fd_sc_hd__clkbuf_1 _3510_ (.A(_1669_),
    .X(_0374_));
 sky130_fd_sc_hd__mux2_1 _3511_ (.A0(\tms1x00.RAM[55][2] ),
    .A1(_1653_),
    .S(_1667_),
    .X(_1670_));
 sky130_fd_sc_hd__clkbuf_1 _3512_ (.A(_1670_),
    .X(_0375_));
 sky130_fd_sc_hd__mux2_1 _3513_ (.A0(\tms1x00.RAM[55][3] ),
    .A1(_1655_),
    .S(_1667_),
    .X(_1671_));
 sky130_fd_sc_hd__clkbuf_1 _3514_ (.A(_1671_),
    .X(_0376_));
 sky130_fd_sc_hd__nor2_2 _3515_ (.A(_0639_),
    .B(_1149_),
    .Y(_1672_));
 sky130_fd_sc_hd__nand2_2 _3516_ (.A(_1672_),
    .B(_1170_),
    .Y(_1673_));
 sky130_fd_sc_hd__mux2_1 _3517_ (.A0(_1563_),
    .A1(\tms1x00.RAM[63][0] ),
    .S(_1673_),
    .X(_1674_));
 sky130_fd_sc_hd__clkbuf_1 _3518_ (.A(_1674_),
    .X(_0377_));
 sky130_fd_sc_hd__mux2_1 _3519_ (.A0(_1566_),
    .A1(\tms1x00.RAM[63][1] ),
    .S(_1673_),
    .X(_1675_));
 sky130_fd_sc_hd__clkbuf_1 _3520_ (.A(_1675_),
    .X(_0378_));
 sky130_fd_sc_hd__mux2_1 _3521_ (.A0(_1568_),
    .A1(\tms1x00.RAM[63][2] ),
    .S(_1673_),
    .X(_1676_));
 sky130_fd_sc_hd__clkbuf_1 _3522_ (.A(_1676_),
    .X(_0379_));
 sky130_fd_sc_hd__mux2_1 _3523_ (.A0(_1570_),
    .A1(\tms1x00.RAM[63][3] ),
    .S(_1673_),
    .X(_1677_));
 sky130_fd_sc_hd__clkbuf_1 _3524_ (.A(_1677_),
    .X(_0380_));
 sky130_fd_sc_hd__nand2_2 _3525_ (.A(_1672_),
    .B(_1213_),
    .Y(_1678_));
 sky130_fd_sc_hd__mux2_1 _3526_ (.A0(_1563_),
    .A1(\tms1x00.RAM[62][0] ),
    .S(_1678_),
    .X(_1679_));
 sky130_fd_sc_hd__clkbuf_1 _3527_ (.A(_1679_),
    .X(_0381_));
 sky130_fd_sc_hd__mux2_1 _3528_ (.A0(_1566_),
    .A1(\tms1x00.RAM[62][1] ),
    .S(_1678_),
    .X(_1680_));
 sky130_fd_sc_hd__clkbuf_1 _3529_ (.A(_1680_),
    .X(_0382_));
 sky130_fd_sc_hd__mux2_1 _3530_ (.A0(_1568_),
    .A1(\tms1x00.RAM[62][2] ),
    .S(_1678_),
    .X(_1681_));
 sky130_fd_sc_hd__clkbuf_1 _3531_ (.A(_1681_),
    .X(_0383_));
 sky130_fd_sc_hd__mux2_1 _3532_ (.A0(_1570_),
    .A1(\tms1x00.RAM[62][3] ),
    .S(_1678_),
    .X(_1682_));
 sky130_fd_sc_hd__clkbuf_1 _3533_ (.A(_1682_),
    .X(_0384_));
 sky130_fd_sc_hd__clkbuf_4 _3534_ (.A(_0826_),
    .X(_1683_));
 sky130_fd_sc_hd__nand2_2 _3535_ (.A(_1672_),
    .B(_1162_),
    .Y(_1684_));
 sky130_fd_sc_hd__mux2_1 _3536_ (.A0(_1683_),
    .A1(\tms1x00.RAM[61][0] ),
    .S(_1684_),
    .X(_1685_));
 sky130_fd_sc_hd__clkbuf_1 _3537_ (.A(_1685_),
    .X(_0385_));
 sky130_fd_sc_hd__clkbuf_4 _3538_ (.A(_0934_),
    .X(_1686_));
 sky130_fd_sc_hd__mux2_1 _3539_ (.A0(_1686_),
    .A1(\tms1x00.RAM[61][1] ),
    .S(_1684_),
    .X(_1687_));
 sky130_fd_sc_hd__clkbuf_1 _3540_ (.A(_1687_),
    .X(_0386_));
 sky130_fd_sc_hd__clkbuf_4 _3541_ (.A(_1034_),
    .X(_1688_));
 sky130_fd_sc_hd__mux2_1 _3542_ (.A0(_1688_),
    .A1(\tms1x00.RAM[61][2] ),
    .S(_1684_),
    .X(_1689_));
 sky130_fd_sc_hd__clkbuf_1 _3543_ (.A(_1689_),
    .X(_0387_));
 sky130_fd_sc_hd__buf_2 _3544_ (.A(_1132_),
    .X(_1690_));
 sky130_fd_sc_hd__mux2_1 _3545_ (.A0(_1690_),
    .A1(\tms1x00.RAM[61][3] ),
    .S(_1684_),
    .X(_1691_));
 sky130_fd_sc_hd__clkbuf_1 _3546_ (.A(_1691_),
    .X(_0388_));
 sky130_fd_sc_hd__nand2_1 _3547_ (.A(_1672_),
    .B(_1224_),
    .Y(_1692_));
 sky130_fd_sc_hd__mux2_1 _3548_ (.A0(_1683_),
    .A1(\tms1x00.RAM[60][0] ),
    .S(_1692_),
    .X(_1693_));
 sky130_fd_sc_hd__clkbuf_1 _3549_ (.A(_1693_),
    .X(_0389_));
 sky130_fd_sc_hd__mux2_1 _3550_ (.A0(_1686_),
    .A1(\tms1x00.RAM[60][1] ),
    .S(_1692_),
    .X(_1694_));
 sky130_fd_sc_hd__clkbuf_1 _3551_ (.A(_1694_),
    .X(_0390_));
 sky130_fd_sc_hd__mux2_1 _3552_ (.A0(_1688_),
    .A1(\tms1x00.RAM[60][2] ),
    .S(_1692_),
    .X(_1695_));
 sky130_fd_sc_hd__clkbuf_1 _3553_ (.A(_1695_),
    .X(_0391_));
 sky130_fd_sc_hd__mux2_1 _3554_ (.A0(_1690_),
    .A1(\tms1x00.RAM[60][3] ),
    .S(_1692_),
    .X(_1696_));
 sky130_fd_sc_hd__clkbuf_1 _3555_ (.A(_1696_),
    .X(_0392_));
 sky130_fd_sc_hd__nor2_2 _3556_ (.A(_1180_),
    .B(_1243_),
    .Y(_1697_));
 sky130_fd_sc_hd__mux2_1 _3557_ (.A0(\tms1x00.RAM[5][0] ),
    .A1(_1648_),
    .S(_1697_),
    .X(_1698_));
 sky130_fd_sc_hd__clkbuf_1 _3558_ (.A(_1698_),
    .X(_0393_));
 sky130_fd_sc_hd__mux2_1 _3559_ (.A0(\tms1x00.RAM[5][1] ),
    .A1(_1651_),
    .S(_1697_),
    .X(_1699_));
 sky130_fd_sc_hd__clkbuf_1 _3560_ (.A(_1699_),
    .X(_0394_));
 sky130_fd_sc_hd__mux2_1 _3561_ (.A0(\tms1x00.RAM[5][2] ),
    .A1(_1653_),
    .S(_1697_),
    .X(_1700_));
 sky130_fd_sc_hd__clkbuf_1 _3562_ (.A(_1700_),
    .X(_0395_));
 sky130_fd_sc_hd__mux2_1 _3563_ (.A0(\tms1x00.RAM[5][3] ),
    .A1(_1655_),
    .S(_1697_),
    .X(_1701_));
 sky130_fd_sc_hd__clkbuf_1 _3564_ (.A(_1701_),
    .X(_0396_));
 sky130_fd_sc_hd__or2_2 _3565_ (.A(_0833_),
    .B(_1176_),
    .X(_1702_));
 sky130_fd_sc_hd__mux2_1 _3566_ (.A0(_1683_),
    .A1(\tms1x00.RAM[67][0] ),
    .S(_1702_),
    .X(_1703_));
 sky130_fd_sc_hd__clkbuf_1 _3567_ (.A(_1703_),
    .X(_0397_));
 sky130_fd_sc_hd__mux2_1 _3568_ (.A0(_1686_),
    .A1(\tms1x00.RAM[67][1] ),
    .S(_1702_),
    .X(_1704_));
 sky130_fd_sc_hd__clkbuf_1 _3569_ (.A(_1704_),
    .X(_0398_));
 sky130_fd_sc_hd__mux2_1 _3570_ (.A0(_1688_),
    .A1(\tms1x00.RAM[67][2] ),
    .S(_1702_),
    .X(_1705_));
 sky130_fd_sc_hd__clkbuf_1 _3571_ (.A(_1705_),
    .X(_0399_));
 sky130_fd_sc_hd__mux2_1 _3572_ (.A0(_1690_),
    .A1(\tms1x00.RAM[67][3] ),
    .S(_1702_),
    .X(_1706_));
 sky130_fd_sc_hd__clkbuf_1 _3573_ (.A(_1706_),
    .X(_0400_));
 sky130_fd_sc_hd__or2_2 _3574_ (.A(_1177_),
    .B(_1320_),
    .X(_1707_));
 sky130_fd_sc_hd__mux2_1 _3575_ (.A0(_1683_),
    .A1(\tms1x00.RAM[66][0] ),
    .S(_1707_),
    .X(_1708_));
 sky130_fd_sc_hd__clkbuf_1 _3576_ (.A(_1708_),
    .X(_0401_));
 sky130_fd_sc_hd__mux2_1 _3577_ (.A0(_1686_),
    .A1(\tms1x00.RAM[66][1] ),
    .S(_1707_),
    .X(_1709_));
 sky130_fd_sc_hd__clkbuf_1 _3578_ (.A(_1709_),
    .X(_0402_));
 sky130_fd_sc_hd__mux2_1 _3579_ (.A0(_1688_),
    .A1(\tms1x00.RAM[66][2] ),
    .S(_1707_),
    .X(_1710_));
 sky130_fd_sc_hd__clkbuf_1 _3580_ (.A(_1710_),
    .X(_0403_));
 sky130_fd_sc_hd__mux2_1 _3581_ (.A0(_1690_),
    .A1(\tms1x00.RAM[66][3] ),
    .S(_1707_),
    .X(_1711_));
 sky130_fd_sc_hd__clkbuf_1 _3582_ (.A(_1711_),
    .X(_0404_));
 sky130_fd_sc_hd__or2_2 _3583_ (.A(_1177_),
    .B(_1194_),
    .X(_1712_));
 sky130_fd_sc_hd__mux2_1 _3584_ (.A0(_1683_),
    .A1(\tms1x00.RAM[65][0] ),
    .S(_1712_),
    .X(_1713_));
 sky130_fd_sc_hd__clkbuf_1 _3585_ (.A(_1713_),
    .X(_0405_));
 sky130_fd_sc_hd__mux2_1 _3586_ (.A0(_1686_),
    .A1(\tms1x00.RAM[65][1] ),
    .S(_1712_),
    .X(_1714_));
 sky130_fd_sc_hd__clkbuf_1 _3587_ (.A(_1714_),
    .X(_0406_));
 sky130_fd_sc_hd__mux2_1 _3588_ (.A0(_1688_),
    .A1(\tms1x00.RAM[65][2] ),
    .S(_1712_),
    .X(_1715_));
 sky130_fd_sc_hd__clkbuf_1 _3589_ (.A(_1715_),
    .X(_0407_));
 sky130_fd_sc_hd__mux2_1 _3590_ (.A0(_1690_),
    .A1(\tms1x00.RAM[65][3] ),
    .S(_1712_),
    .X(_1716_));
 sky130_fd_sc_hd__clkbuf_1 _3591_ (.A(_1716_),
    .X(_0408_));
 sky130_fd_sc_hd__or2_2 _3592_ (.A(_1176_),
    .B(_1311_),
    .X(_1717_));
 sky130_fd_sc_hd__mux2_1 _3593_ (.A0(_1683_),
    .A1(\tms1x00.RAM[64][0] ),
    .S(_1717_),
    .X(_1718_));
 sky130_fd_sc_hd__clkbuf_1 _3594_ (.A(_1718_),
    .X(_0409_));
 sky130_fd_sc_hd__mux2_1 _3595_ (.A0(_1686_),
    .A1(\tms1x00.RAM[64][1] ),
    .S(_1717_),
    .X(_1719_));
 sky130_fd_sc_hd__clkbuf_1 _3596_ (.A(_1719_),
    .X(_0410_));
 sky130_fd_sc_hd__mux2_1 _3597_ (.A0(_1688_),
    .A1(\tms1x00.RAM[64][2] ),
    .S(_1717_),
    .X(_1720_));
 sky130_fd_sc_hd__clkbuf_1 _3598_ (.A(_1720_),
    .X(_0411_));
 sky130_fd_sc_hd__mux2_1 _3599_ (.A0(_1690_),
    .A1(\tms1x00.RAM[64][3] ),
    .S(_1717_),
    .X(_1721_));
 sky130_fd_sc_hd__clkbuf_1 _3600_ (.A(_1721_),
    .X(_0412_));
 sky130_fd_sc_hd__nor2_2 _3601_ (.A(_1177_),
    .B(_1257_),
    .Y(_1722_));
 sky130_fd_sc_hd__mux2_1 _3602_ (.A0(\tms1x00.RAM[71][0] ),
    .A1(_1648_),
    .S(_1722_),
    .X(_1723_));
 sky130_fd_sc_hd__clkbuf_1 _3603_ (.A(_1723_),
    .X(_0413_));
 sky130_fd_sc_hd__mux2_1 _3604_ (.A0(\tms1x00.RAM[71][1] ),
    .A1(_1651_),
    .S(_1722_),
    .X(_1724_));
 sky130_fd_sc_hd__clkbuf_1 _3605_ (.A(_1724_),
    .X(_0414_));
 sky130_fd_sc_hd__mux2_1 _3606_ (.A0(\tms1x00.RAM[71][2] ),
    .A1(_1653_),
    .S(_1722_),
    .X(_1725_));
 sky130_fd_sc_hd__clkbuf_1 _3607_ (.A(_1725_),
    .X(_0415_));
 sky130_fd_sc_hd__mux2_1 _3608_ (.A0(\tms1x00.RAM[71][3] ),
    .A1(_1655_),
    .S(_1722_),
    .X(_1726_));
 sky130_fd_sc_hd__clkbuf_1 _3609_ (.A(_1726_),
    .X(_0416_));
 sky130_fd_sc_hd__nor2_2 _3610_ (.A(_1177_),
    .B(_1266_),
    .Y(_1727_));
 sky130_fd_sc_hd__mux2_1 _3611_ (.A0(\tms1x00.RAM[70][0] ),
    .A1(_1648_),
    .S(_1727_),
    .X(_1728_));
 sky130_fd_sc_hd__clkbuf_1 _3612_ (.A(_1728_),
    .X(_0417_));
 sky130_fd_sc_hd__mux2_1 _3613_ (.A0(\tms1x00.RAM[70][1] ),
    .A1(_1651_),
    .S(_1727_),
    .X(_1729_));
 sky130_fd_sc_hd__clkbuf_1 _3614_ (.A(_1729_),
    .X(_0418_));
 sky130_fd_sc_hd__mux2_1 _3615_ (.A0(\tms1x00.RAM[70][2] ),
    .A1(_1653_),
    .S(_1727_),
    .X(_1730_));
 sky130_fd_sc_hd__clkbuf_1 _3616_ (.A(_1730_),
    .X(_0419_));
 sky130_fd_sc_hd__mux2_1 _3617_ (.A0(\tms1x00.RAM[70][3] ),
    .A1(_1655_),
    .S(_1727_),
    .X(_1731_));
 sky130_fd_sc_hd__clkbuf_1 _3618_ (.A(_1731_),
    .X(_0420_));
 sky130_fd_sc_hd__nor2_2 _3619_ (.A(_1243_),
    .B(_1266_),
    .Y(_1732_));
 sky130_fd_sc_hd__mux2_1 _3620_ (.A0(\tms1x00.RAM[6][0] ),
    .A1(_1648_),
    .S(_1732_),
    .X(_1733_));
 sky130_fd_sc_hd__clkbuf_1 _3621_ (.A(_1733_),
    .X(_0421_));
 sky130_fd_sc_hd__mux2_1 _3622_ (.A0(\tms1x00.RAM[6][1] ),
    .A1(_1651_),
    .S(_1732_),
    .X(_1734_));
 sky130_fd_sc_hd__clkbuf_1 _3623_ (.A(_1734_),
    .X(_0422_));
 sky130_fd_sc_hd__mux2_1 _3624_ (.A0(\tms1x00.RAM[6][2] ),
    .A1(_1653_),
    .S(_1732_),
    .X(_1735_));
 sky130_fd_sc_hd__clkbuf_1 _3625_ (.A(_1735_),
    .X(_0423_));
 sky130_fd_sc_hd__mux2_1 _3626_ (.A0(\tms1x00.RAM[6][3] ),
    .A1(_1655_),
    .S(_1732_),
    .X(_1736_));
 sky130_fd_sc_hd__clkbuf_1 _3627_ (.A(_1736_),
    .X(_0424_));
 sky130_fd_sc_hd__nor2_2 _3628_ (.A(_1177_),
    .B(_1304_),
    .Y(_1737_));
 sky130_fd_sc_hd__mux2_1 _3629_ (.A0(\tms1x00.RAM[68][0] ),
    .A1(_1648_),
    .S(_1737_),
    .X(_1738_));
 sky130_fd_sc_hd__clkbuf_1 _3630_ (.A(_1738_),
    .X(_0425_));
 sky130_fd_sc_hd__mux2_1 _3631_ (.A0(\tms1x00.RAM[68][1] ),
    .A1(_1651_),
    .S(_1737_),
    .X(_1739_));
 sky130_fd_sc_hd__clkbuf_1 _3632_ (.A(_1739_),
    .X(_0426_));
 sky130_fd_sc_hd__mux2_1 _3633_ (.A0(\tms1x00.RAM[68][2] ),
    .A1(_1653_),
    .S(_1737_),
    .X(_1740_));
 sky130_fd_sc_hd__clkbuf_1 _3634_ (.A(_1740_),
    .X(_0427_));
 sky130_fd_sc_hd__mux2_1 _3635_ (.A0(\tms1x00.RAM[68][3] ),
    .A1(_1655_),
    .S(_1737_),
    .X(_1741_));
 sky130_fd_sc_hd__clkbuf_1 _3636_ (.A(_1741_),
    .X(_0428_));
 sky130_fd_sc_hd__nand2_2 _3637_ (.A(_1168_),
    .B(_1224_),
    .Y(_1742_));
 sky130_fd_sc_hd__mux2_1 _3638_ (.A0(_1683_),
    .A1(\tms1x00.RAM[76][0] ),
    .S(_1742_),
    .X(_1743_));
 sky130_fd_sc_hd__clkbuf_1 _3639_ (.A(_1743_),
    .X(_0429_));
 sky130_fd_sc_hd__mux2_1 _3640_ (.A0(_1686_),
    .A1(\tms1x00.RAM[76][1] ),
    .S(_1742_),
    .X(_1744_));
 sky130_fd_sc_hd__clkbuf_1 _3641_ (.A(_1744_),
    .X(_0430_));
 sky130_fd_sc_hd__mux2_1 _3642_ (.A0(_1688_),
    .A1(\tms1x00.RAM[76][2] ),
    .S(_1742_),
    .X(_1745_));
 sky130_fd_sc_hd__clkbuf_1 _3643_ (.A(_1745_),
    .X(_0431_));
 sky130_fd_sc_hd__mux2_1 _3644_ (.A0(_1690_),
    .A1(\tms1x00.RAM[76][3] ),
    .S(_1742_),
    .X(_1746_));
 sky130_fd_sc_hd__clkbuf_1 _3645_ (.A(_1746_),
    .X(_0432_));
 sky130_fd_sc_hd__nor2_1 _3646_ (.A(_1153_),
    .B(_1177_),
    .Y(_1747_));
 sky130_fd_sc_hd__mux2_1 _3647_ (.A0(\tms1x00.RAM[75][0] ),
    .A1(_1648_),
    .S(_1747_),
    .X(_1748_));
 sky130_fd_sc_hd__clkbuf_1 _3648_ (.A(_1748_),
    .X(_0433_));
 sky130_fd_sc_hd__mux2_1 _3649_ (.A0(\tms1x00.RAM[75][1] ),
    .A1(_1651_),
    .S(_1747_),
    .X(_1749_));
 sky130_fd_sc_hd__clkbuf_1 _3650_ (.A(_1749_),
    .X(_0434_));
 sky130_fd_sc_hd__mux2_1 _3651_ (.A0(\tms1x00.RAM[75][2] ),
    .A1(_1653_),
    .S(_1747_),
    .X(_1750_));
 sky130_fd_sc_hd__clkbuf_1 _3652_ (.A(_1750_),
    .X(_0435_));
 sky130_fd_sc_hd__mux2_1 _3653_ (.A0(\tms1x00.RAM[75][3] ),
    .A1(_1655_),
    .S(_1747_),
    .X(_1751_));
 sky130_fd_sc_hd__clkbuf_1 _3654_ (.A(_1751_),
    .X(_0436_));
 sky130_fd_sc_hd__nor2_2 _3655_ (.A(_1177_),
    .B(_1236_),
    .Y(_1752_));
 sky130_fd_sc_hd__mux2_1 _3656_ (.A0(\tms1x00.RAM[74][0] ),
    .A1(_1263_),
    .S(_1752_),
    .X(_1753_));
 sky130_fd_sc_hd__clkbuf_1 _3657_ (.A(_1753_),
    .X(_0437_));
 sky130_fd_sc_hd__mux2_1 _3658_ (.A0(\tms1x00.RAM[74][1] ),
    .A1(_1269_),
    .S(_1752_),
    .X(_1754_));
 sky130_fd_sc_hd__clkbuf_1 _3659_ (.A(_1754_),
    .X(_0438_));
 sky130_fd_sc_hd__mux2_1 _3660_ (.A0(\tms1x00.RAM[74][2] ),
    .A1(_1272_),
    .S(_1752_),
    .X(_1755_));
 sky130_fd_sc_hd__clkbuf_1 _3661_ (.A(_1755_),
    .X(_0439_));
 sky130_fd_sc_hd__mux2_1 _3662_ (.A0(\tms1x00.RAM[74][3] ),
    .A1(_1275_),
    .S(_1752_),
    .X(_1756_));
 sky130_fd_sc_hd__clkbuf_1 _3663_ (.A(_1756_),
    .X(_0440_));
 sky130_fd_sc_hd__nor2_2 _3664_ (.A(_1140_),
    .B(_1177_),
    .Y(_1757_));
 sky130_fd_sc_hd__mux2_1 _3665_ (.A0(\tms1x00.RAM[73][0] ),
    .A1(_1263_),
    .S(_1757_),
    .X(_1758_));
 sky130_fd_sc_hd__clkbuf_1 _3666_ (.A(_1758_),
    .X(_0441_));
 sky130_fd_sc_hd__mux2_1 _3667_ (.A0(\tms1x00.RAM[73][1] ),
    .A1(_1269_),
    .S(_1757_),
    .X(_1759_));
 sky130_fd_sc_hd__clkbuf_1 _3668_ (.A(_1759_),
    .X(_0442_));
 sky130_fd_sc_hd__mux2_1 _3669_ (.A0(\tms1x00.RAM[73][2] ),
    .A1(_1272_),
    .S(_1757_),
    .X(_1760_));
 sky130_fd_sc_hd__clkbuf_1 _3670_ (.A(_1760_),
    .X(_0443_));
 sky130_fd_sc_hd__mux2_1 _3671_ (.A0(\tms1x00.RAM[73][3] ),
    .A1(_1275_),
    .S(_1757_),
    .X(_1761_));
 sky130_fd_sc_hd__clkbuf_1 _3672_ (.A(_1761_),
    .X(_0444_));
 sky130_fd_sc_hd__nor2_2 _3673_ (.A(_1177_),
    .B(_1245_),
    .Y(_1762_));
 sky130_fd_sc_hd__mux2_1 _3674_ (.A0(\tms1x00.RAM[72][0] ),
    .A1(_1263_),
    .S(_1762_),
    .X(_1763_));
 sky130_fd_sc_hd__clkbuf_1 _3675_ (.A(_1763_),
    .X(_0445_));
 sky130_fd_sc_hd__mux2_1 _3676_ (.A0(\tms1x00.RAM[72][1] ),
    .A1(_1269_),
    .S(_1762_),
    .X(_1764_));
 sky130_fd_sc_hd__clkbuf_1 _3677_ (.A(_1764_),
    .X(_0446_));
 sky130_fd_sc_hd__mux2_1 _3678_ (.A0(\tms1x00.RAM[72][2] ),
    .A1(_1272_),
    .S(_1762_),
    .X(_1765_));
 sky130_fd_sc_hd__clkbuf_1 _3679_ (.A(_1765_),
    .X(_0447_));
 sky130_fd_sc_hd__mux2_1 _3680_ (.A0(\tms1x00.RAM[72][3] ),
    .A1(_1275_),
    .S(_1762_),
    .X(_1766_));
 sky130_fd_sc_hd__clkbuf_1 _3681_ (.A(_1766_),
    .X(_0448_));
 sky130_fd_sc_hd__nand2_2 _3682_ (.A(_1162_),
    .B(_1168_),
    .Y(_1767_));
 sky130_fd_sc_hd__mux2_1 _3683_ (.A0(_1683_),
    .A1(\tms1x00.RAM[77][0] ),
    .S(_1767_),
    .X(_1768_));
 sky130_fd_sc_hd__clkbuf_1 _3684_ (.A(_1768_),
    .X(_0449_));
 sky130_fd_sc_hd__mux2_1 _3685_ (.A0(_1686_),
    .A1(\tms1x00.RAM[77][1] ),
    .S(_1767_),
    .X(_1769_));
 sky130_fd_sc_hd__clkbuf_1 _3686_ (.A(_1769_),
    .X(_0450_));
 sky130_fd_sc_hd__mux2_1 _3687_ (.A0(_1688_),
    .A1(\tms1x00.RAM[77][2] ),
    .S(_1767_),
    .X(_1770_));
 sky130_fd_sc_hd__clkbuf_1 _3688_ (.A(_1770_),
    .X(_0451_));
 sky130_fd_sc_hd__mux2_1 _3689_ (.A0(_1690_),
    .A1(\tms1x00.RAM[77][3] ),
    .S(_1767_),
    .X(_1771_));
 sky130_fd_sc_hd__clkbuf_1 _3690_ (.A(_1771_),
    .X(_0452_));
 sky130_fd_sc_hd__or2_2 _3691_ (.A(_1137_),
    .B(_1311_),
    .X(_1772_));
 sky130_fd_sc_hd__mux2_1 _3692_ (.A0(_1683_),
    .A1(\tms1x00.RAM[80][0] ),
    .S(_1772_),
    .X(_1773_));
 sky130_fd_sc_hd__clkbuf_1 _3693_ (.A(_1773_),
    .X(_0453_));
 sky130_fd_sc_hd__mux2_1 _3694_ (.A0(_1686_),
    .A1(\tms1x00.RAM[80][1] ),
    .S(_1772_),
    .X(_1774_));
 sky130_fd_sc_hd__clkbuf_1 _3695_ (.A(_1774_),
    .X(_0454_));
 sky130_fd_sc_hd__mux2_1 _3696_ (.A0(_1688_),
    .A1(\tms1x00.RAM[80][2] ),
    .S(_1772_),
    .X(_1775_));
 sky130_fd_sc_hd__clkbuf_1 _3697_ (.A(_1775_),
    .X(_0455_));
 sky130_fd_sc_hd__mux2_1 _3698_ (.A0(_1690_),
    .A1(\tms1x00.RAM[80][3] ),
    .S(_1772_),
    .X(_1776_));
 sky130_fd_sc_hd__clkbuf_1 _3699_ (.A(_1776_),
    .X(_0456_));
 sky130_fd_sc_hd__nor2_2 _3700_ (.A(_1243_),
    .B(_1257_),
    .Y(_1777_));
 sky130_fd_sc_hd__mux2_1 _3701_ (.A0(\tms1x00.RAM[7][0] ),
    .A1(_1263_),
    .S(_1777_),
    .X(_1778_));
 sky130_fd_sc_hd__clkbuf_1 _3702_ (.A(_1778_),
    .X(_0457_));
 sky130_fd_sc_hd__mux2_1 _3703_ (.A0(\tms1x00.RAM[7][1] ),
    .A1(_1269_),
    .S(_1777_),
    .X(_1779_));
 sky130_fd_sc_hd__clkbuf_1 _3704_ (.A(_1779_),
    .X(_0458_));
 sky130_fd_sc_hd__mux2_1 _3705_ (.A0(\tms1x00.RAM[7][2] ),
    .A1(_1272_),
    .S(_1777_),
    .X(_1780_));
 sky130_fd_sc_hd__clkbuf_1 _3706_ (.A(_1780_),
    .X(_0459_));
 sky130_fd_sc_hd__mux2_1 _3707_ (.A0(\tms1x00.RAM[7][3] ),
    .A1(_1275_),
    .S(_1777_),
    .X(_1781_));
 sky130_fd_sc_hd__clkbuf_1 _3708_ (.A(_1781_),
    .X(_0460_));
 sky130_fd_sc_hd__nand2_1 _3709_ (.A(_1168_),
    .B(_1213_),
    .Y(_1782_));
 sky130_fd_sc_hd__mux2_1 _3710_ (.A0(_1683_),
    .A1(\tms1x00.RAM[78][0] ),
    .S(_1782_),
    .X(_1783_));
 sky130_fd_sc_hd__clkbuf_1 _3711_ (.A(_1783_),
    .X(_0461_));
 sky130_fd_sc_hd__mux2_1 _3712_ (.A0(_1686_),
    .A1(\tms1x00.RAM[78][1] ),
    .S(_1782_),
    .X(_1784_));
 sky130_fd_sc_hd__clkbuf_1 _3713_ (.A(_1784_),
    .X(_0462_));
 sky130_fd_sc_hd__mux2_1 _3714_ (.A0(_1688_),
    .A1(\tms1x00.RAM[78][2] ),
    .S(_1782_),
    .X(_1785_));
 sky130_fd_sc_hd__clkbuf_1 _3715_ (.A(_1785_),
    .X(_0463_));
 sky130_fd_sc_hd__mux2_1 _3716_ (.A0(_1690_),
    .A1(\tms1x00.RAM[78][3] ),
    .S(_1782_),
    .X(_1786_));
 sky130_fd_sc_hd__clkbuf_1 _3717_ (.A(_1786_),
    .X(_0464_));
 sky130_fd_sc_hd__nor2_2 _3718_ (.A(_1137_),
    .B(_1180_),
    .Y(_1787_));
 sky130_fd_sc_hd__mux2_1 _3719_ (.A0(\tms1x00.RAM[85][0] ),
    .A1(_1263_),
    .S(_1787_),
    .X(_1788_));
 sky130_fd_sc_hd__clkbuf_1 _3720_ (.A(_1788_),
    .X(_0465_));
 sky130_fd_sc_hd__mux2_1 _3721_ (.A0(\tms1x00.RAM[85][1] ),
    .A1(_1269_),
    .S(_1787_),
    .X(_1789_));
 sky130_fd_sc_hd__clkbuf_1 _3722_ (.A(_1789_),
    .X(_0466_));
 sky130_fd_sc_hd__mux2_1 _3723_ (.A0(\tms1x00.RAM[85][2] ),
    .A1(_1272_),
    .S(_1787_),
    .X(_1790_));
 sky130_fd_sc_hd__clkbuf_1 _3724_ (.A(_1790_),
    .X(_0467_));
 sky130_fd_sc_hd__mux2_1 _3725_ (.A0(\tms1x00.RAM[85][3] ),
    .A1(_1275_),
    .S(_1787_),
    .X(_1791_));
 sky130_fd_sc_hd__clkbuf_1 _3726_ (.A(_1791_),
    .X(_0468_));
 sky130_fd_sc_hd__nor2_2 _3727_ (.A(_1137_),
    .B(_1304_),
    .Y(_1792_));
 sky130_fd_sc_hd__mux2_1 _3728_ (.A0(\tms1x00.RAM[84][0] ),
    .A1(_1263_),
    .S(_1792_),
    .X(_1793_));
 sky130_fd_sc_hd__clkbuf_1 _3729_ (.A(_1793_),
    .X(_0469_));
 sky130_fd_sc_hd__mux2_1 _3730_ (.A0(\tms1x00.RAM[84][1] ),
    .A1(_1269_),
    .S(_1792_),
    .X(_1794_));
 sky130_fd_sc_hd__clkbuf_1 _3731_ (.A(_1794_),
    .X(_0470_));
 sky130_fd_sc_hd__mux2_1 _3732_ (.A0(\tms1x00.RAM[84][2] ),
    .A1(_1272_),
    .S(_1792_),
    .X(_1795_));
 sky130_fd_sc_hd__clkbuf_1 _3733_ (.A(_1795_),
    .X(_0471_));
 sky130_fd_sc_hd__mux2_1 _3734_ (.A0(\tms1x00.RAM[84][3] ),
    .A1(_1275_),
    .S(_1792_),
    .X(_1796_));
 sky130_fd_sc_hd__clkbuf_1 _3735_ (.A(_1796_),
    .X(_0472_));
 sky130_fd_sc_hd__clkbuf_4 _3736_ (.A(_0826_),
    .X(_1797_));
 sky130_fd_sc_hd__or2_2 _3737_ (.A(_0833_),
    .B(_1136_),
    .X(_1798_));
 sky130_fd_sc_hd__mux2_1 _3738_ (.A0(_1797_),
    .A1(\tms1x00.RAM[83][0] ),
    .S(_1798_),
    .X(_1799_));
 sky130_fd_sc_hd__clkbuf_1 _3739_ (.A(_1799_),
    .X(_0473_));
 sky130_fd_sc_hd__clkbuf_4 _3740_ (.A(_0934_),
    .X(_1800_));
 sky130_fd_sc_hd__mux2_1 _3741_ (.A0(_1800_),
    .A1(\tms1x00.RAM[83][1] ),
    .S(_1798_),
    .X(_1801_));
 sky130_fd_sc_hd__clkbuf_1 _3742_ (.A(_1801_),
    .X(_0474_));
 sky130_fd_sc_hd__clkbuf_4 _3743_ (.A(_1034_),
    .X(_1802_));
 sky130_fd_sc_hd__mux2_1 _3744_ (.A0(_1802_),
    .A1(\tms1x00.RAM[83][2] ),
    .S(_1798_),
    .X(_1803_));
 sky130_fd_sc_hd__clkbuf_1 _3745_ (.A(_1803_),
    .X(_0475_));
 sky130_fd_sc_hd__clkbuf_4 _3746_ (.A(_1132_),
    .X(_1804_));
 sky130_fd_sc_hd__mux2_1 _3747_ (.A0(_1804_),
    .A1(\tms1x00.RAM[83][3] ),
    .S(_1798_),
    .X(_1805_));
 sky130_fd_sc_hd__clkbuf_1 _3748_ (.A(_1805_),
    .X(_0476_));
 sky130_fd_sc_hd__or2_2 _3749_ (.A(_1137_),
    .B(_1320_),
    .X(_1806_));
 sky130_fd_sc_hd__mux2_1 _3750_ (.A0(_1797_),
    .A1(\tms1x00.RAM[82][0] ),
    .S(_1806_),
    .X(_1807_));
 sky130_fd_sc_hd__clkbuf_1 _3751_ (.A(_1807_),
    .X(_0477_));
 sky130_fd_sc_hd__mux2_1 _3752_ (.A0(_1800_),
    .A1(\tms1x00.RAM[82][1] ),
    .S(_1806_),
    .X(_1808_));
 sky130_fd_sc_hd__clkbuf_1 _3753_ (.A(_1808_),
    .X(_0478_));
 sky130_fd_sc_hd__mux2_1 _3754_ (.A0(_1802_),
    .A1(\tms1x00.RAM[82][2] ),
    .S(_1806_),
    .X(_1809_));
 sky130_fd_sc_hd__clkbuf_1 _3755_ (.A(_1809_),
    .X(_0479_));
 sky130_fd_sc_hd__mux2_1 _3756_ (.A0(_1804_),
    .A1(\tms1x00.RAM[82][3] ),
    .S(_1806_),
    .X(_1810_));
 sky130_fd_sc_hd__clkbuf_1 _3757_ (.A(_1810_),
    .X(_0480_));
 sky130_fd_sc_hd__or2_2 _3758_ (.A(_1136_),
    .B(_1194_),
    .X(_1811_));
 sky130_fd_sc_hd__mux2_1 _3759_ (.A0(_1797_),
    .A1(\tms1x00.RAM[81][0] ),
    .S(_1811_),
    .X(_1812_));
 sky130_fd_sc_hd__clkbuf_1 _3760_ (.A(_1812_),
    .X(_0481_));
 sky130_fd_sc_hd__mux2_1 _3761_ (.A0(_1800_),
    .A1(\tms1x00.RAM[81][1] ),
    .S(_1811_),
    .X(_1813_));
 sky130_fd_sc_hd__clkbuf_1 _3762_ (.A(_1813_),
    .X(_0482_));
 sky130_fd_sc_hd__mux2_1 _3763_ (.A0(_1802_),
    .A1(\tms1x00.RAM[81][2] ),
    .S(_1811_),
    .X(_1814_));
 sky130_fd_sc_hd__clkbuf_1 _3764_ (.A(_1814_),
    .X(_0483_));
 sky130_fd_sc_hd__mux2_1 _3765_ (.A0(_1804_),
    .A1(\tms1x00.RAM[81][3] ),
    .S(_1811_),
    .X(_1815_));
 sky130_fd_sc_hd__clkbuf_1 _3766_ (.A(_1815_),
    .X(_0484_));
 sky130_fd_sc_hd__mux2_1 _3767_ (.A0(_0619_),
    .A1(_0620_),
    .S(_0625_),
    .X(_1816_));
 sky130_fd_sc_hd__clkbuf_1 _3768_ (.A(_1816_),
    .X(_0485_));
 sky130_fd_sc_hd__mux2_1 _3769_ (.A0(_0627_),
    .A1(_0628_),
    .S(_0625_),
    .X(_1817_));
 sky130_fd_sc_hd__clkbuf_1 _3770_ (.A(_1817_),
    .X(_0486_));
 sky130_fd_sc_hd__mux2_1 _3771_ (.A0(_0630_),
    .A1(\tms1x00.ram_addr_buff[2] ),
    .S(_0625_),
    .X(_1818_));
 sky130_fd_sc_hd__clkbuf_1 _3772_ (.A(_1818_),
    .X(_0487_));
 sky130_fd_sc_hd__mux2_1 _3773_ (.A0(_0633_),
    .A1(\tms1x00.ram_addr_buff[3] ),
    .S(_0624_),
    .X(_1819_));
 sky130_fd_sc_hd__clkbuf_1 _3774_ (.A(_1819_),
    .X(_0488_));
 sky130_fd_sc_hd__mux2_1 _3775_ (.A0(\tms1x00.X[2] ),
    .A1(_0635_),
    .S(_0624_),
    .X(_1820_));
 sky130_fd_sc_hd__clkbuf_1 _3776_ (.A(_1820_),
    .X(_0489_));
 sky130_fd_sc_hd__mux2_1 _3777_ (.A0(\tms1x00.X[0] ),
    .A1(_0637_),
    .S(_0624_),
    .X(_1821_));
 sky130_fd_sc_hd__clkbuf_1 _3778_ (.A(_1821_),
    .X(_0490_));
 sky130_fd_sc_hd__mux2_1 _3779_ (.A0(\tms1x00.X[1] ),
    .A1(_0639_),
    .S(_0624_),
    .X(_1822_));
 sky130_fd_sc_hd__clkbuf_1 _3780_ (.A(_1822_),
    .X(_0491_));
 sky130_fd_sc_hd__buf_2 _3781_ (.A(net16),
    .X(_1823_));
 sky130_fd_sc_hd__clkbuf_4 _3782_ (.A(_1823_),
    .X(_1824_));
 sky130_fd_sc_hd__nor2_1 _3783_ (.A(net37),
    .B(_1824_),
    .Y(_0492_));
 sky130_fd_sc_hd__xnor2_1 _3784_ (.A(net37),
    .B(net38),
    .Y(_1825_));
 sky130_fd_sc_hd__and3b_1 _3785_ (.A_N(net38),
    .B(net37),
    .C(net39),
    .X(_1826_));
 sky130_fd_sc_hd__nor3_1 _3786_ (.A(_1824_),
    .B(_1825_),
    .C(_1826_),
    .Y(_0493_));
 sky130_fd_sc_hd__a21oi_1 _3787_ (.A1(_0622_),
    .A2(_0647_),
    .B1(_1824_),
    .Y(_0494_));
 sky130_fd_sc_hd__buf_2 _3788_ (.A(\tms1x00.rom_addr[1] ),
    .X(_1827_));
 sky130_fd_sc_hd__mux4_1 _3789_ (.A0(net5),
    .A1(net7),
    .A2(net8),
    .A3(net9),
    .S0(\tms1x00.rom_addr[0] ),
    .S1(_1827_),
    .X(_1828_));
 sky130_fd_sc_hd__mux2_1 _3790_ (.A0(\tms1x00.ins_in[0] ),
    .A1(_1828_),
    .S(_0623_),
    .X(_1829_));
 sky130_fd_sc_hd__or2_1 _3791_ (.A(_1824_),
    .B(_1829_),
    .X(_1830_));
 sky130_fd_sc_hd__clkbuf_1 _3792_ (.A(_1830_),
    .X(_0495_));
 sky130_fd_sc_hd__mux4_1 _3793_ (.A0(net7),
    .A1(net8),
    .A2(net9),
    .A3(net10),
    .S0(\tms1x00.rom_addr[0] ),
    .S1(_1827_),
    .X(_1831_));
 sky130_fd_sc_hd__mux2_1 _3794_ (.A0(\tms1x00.ins_in[1] ),
    .A1(_1831_),
    .S(_0623_),
    .X(_1832_));
 sky130_fd_sc_hd__or2_1 _3795_ (.A(_1824_),
    .B(_1832_),
    .X(_1833_));
 sky130_fd_sc_hd__clkbuf_1 _3796_ (.A(_1833_),
    .X(_0496_));
 sky130_fd_sc_hd__or2_1 _3797_ (.A(net38),
    .B(_0622_),
    .X(_1834_));
 sky130_fd_sc_hd__nor2_1 _3798_ (.A(_1823_),
    .B(_1834_),
    .Y(_1835_));
 sky130_fd_sc_hd__mux2_1 _3799_ (.A0(net10),
    .A1(net11),
    .S(\tms1x00.rom_addr[0] ),
    .X(_1836_));
 sky130_fd_sc_hd__or2b_1 _3800_ (.A(_1836_),
    .B_N(_1827_),
    .X(_1837_));
 sky130_fd_sc_hd__mux2_1 _3801_ (.A0(net8),
    .A1(net9),
    .S(\tms1x00.rom_addr[0] ),
    .X(_1838_));
 sky130_fd_sc_hd__or2_1 _3802_ (.A(_1827_),
    .B(_1838_),
    .X(_1839_));
 sky130_fd_sc_hd__nor2_2 _3803_ (.A(_1823_),
    .B(_0623_),
    .Y(_1840_));
 sky130_fd_sc_hd__a32o_1 _3804_ (.A1(_1835_),
    .A2(_1837_),
    .A3(_1839_),
    .B1(_1840_),
    .B2(\tms1x00.ins_in[2] ),
    .X(_0497_));
 sky130_fd_sc_hd__mux4_1 _3805_ (.A0(net9),
    .A1(net10),
    .A2(net11),
    .A3(net12),
    .S0(\tms1x00.rom_addr[0] ),
    .S1(_1827_),
    .X(_1841_));
 sky130_fd_sc_hd__or2_1 _3806_ (.A(_1834_),
    .B(_1841_),
    .X(_1842_));
 sky130_fd_sc_hd__clkbuf_4 _3807_ (.A(_0621_),
    .X(_1843_));
 sky130_fd_sc_hd__o211a_1 _3808_ (.A1(\tms1x00.ins_in[3] ),
    .A2(_0623_),
    .B1(_1842_),
    .C1(_1843_),
    .X(_0498_));
 sky130_fd_sc_hd__mux2_1 _3809_ (.A0(net12),
    .A1(net13),
    .S(\tms1x00.rom_addr[0] ),
    .X(_1844_));
 sky130_fd_sc_hd__or2b_1 _3810_ (.A(_1844_),
    .B_N(_1827_),
    .X(_1845_));
 sky130_fd_sc_hd__or2_1 _3811_ (.A(_1827_),
    .B(_1836_),
    .X(_1846_));
 sky130_fd_sc_hd__clkbuf_4 _3812_ (.A(\tms1x00.ins_in[4] ),
    .X(_1847_));
 sky130_fd_sc_hd__a32o_1 _3813_ (.A1(_1835_),
    .A2(_1845_),
    .A3(_1846_),
    .B1(_1840_),
    .B2(_1847_),
    .X(_0499_));
 sky130_fd_sc_hd__clkbuf_4 _3814_ (.A(\tms1x00.ins_in[5] ),
    .X(_1848_));
 sky130_fd_sc_hd__mux4_1 _3815_ (.A0(net11),
    .A1(net12),
    .A2(net13),
    .A3(net14),
    .S0(\tms1x00.rom_addr[0] ),
    .S1(\tms1x00.rom_addr[1] ),
    .X(_1849_));
 sky130_fd_sc_hd__mux2_1 _3816_ (.A0(_1848_),
    .A1(_1849_),
    .S(_0623_),
    .X(_1850_));
 sky130_fd_sc_hd__or2_1 _3817_ (.A(_1824_),
    .B(_1850_),
    .X(_1851_));
 sky130_fd_sc_hd__clkbuf_1 _3818_ (.A(_1851_),
    .X(_0500_));
 sky130_fd_sc_hd__mux4_1 _3819_ (.A0(net12),
    .A1(net13),
    .A2(net14),
    .A3(net15),
    .S0(\tms1x00.rom_addr[0] ),
    .S1(_1827_),
    .X(_1852_));
 sky130_fd_sc_hd__or2_1 _3820_ (.A(_1834_),
    .B(_1852_),
    .X(_1853_));
 sky130_fd_sc_hd__o211a_1 _3821_ (.A1(_0643_),
    .A2(_0623_),
    .B1(_1853_),
    .C1(_1843_),
    .X(_0501_));
 sky130_fd_sc_hd__mux4_1 _3822_ (.A0(net13),
    .A1(net14),
    .A2(net15),
    .A3(net6),
    .S0(\tms1x00.rom_addr[0] ),
    .S1(_1827_),
    .X(_1854_));
 sky130_fd_sc_hd__or2_1 _3823_ (.A(_1834_),
    .B(_1854_),
    .X(_1855_));
 sky130_fd_sc_hd__o211a_1 _3824_ (.A1(_0642_),
    .A2(_0623_),
    .B1(_1855_),
    .C1(_1843_),
    .X(_0502_));
 sky130_fd_sc_hd__or3b_1 _3825_ (.A(_0630_),
    .B(_0627_),
    .C_N(_0619_),
    .X(_1856_));
 sky130_fd_sc_hd__nor3b_1 _3826_ (.A(_0630_),
    .B(_0627_),
    .C_N(\tms1x00.Y[0] ),
    .Y(_1857_));
 sky130_fd_sc_hd__a31o_1 _3827_ (.A1(_0651_),
    .A2(_0656_),
    .A3(_1857_),
    .B1(net41),
    .X(_1858_));
 sky130_fd_sc_hd__o311a_1 _3828_ (.A1(_0633_),
    .A2(_0649_),
    .A3(_1856_),
    .B1(_1858_),
    .C1(_0658_),
    .X(_0503_));
 sky130_fd_sc_hd__or3b_1 _3829_ (.A(_0630_),
    .B(_0619_),
    .C_N(_0627_),
    .X(_1859_));
 sky130_fd_sc_hd__nor3b_1 _3830_ (.A(_0630_),
    .B(_0619_),
    .C_N(\tms1x00.Y[1] ),
    .Y(_1860_));
 sky130_fd_sc_hd__a31o_1 _3831_ (.A1(_0651_),
    .A2(_0656_),
    .A3(_1860_),
    .B1(net42),
    .X(_1861_));
 sky130_fd_sc_hd__buf_2 _3832_ (.A(_0621_),
    .X(_1862_));
 sky130_fd_sc_hd__o311a_1 _3833_ (.A1(_0633_),
    .A2(_0649_),
    .A3(_1859_),
    .B1(_1861_),
    .C1(_1862_),
    .X(_0504_));
 sky130_fd_sc_hd__and3b_1 _3834_ (.A_N(\tms1x00.Y[2] ),
    .B(\tms1x00.Y[1] ),
    .C(\tms1x00.Y[0] ),
    .X(_1863_));
 sky130_fd_sc_hd__a31o_1 _3835_ (.A1(_0651_),
    .A2(_0655_),
    .A3(_1863_),
    .B1(net43),
    .X(_1864_));
 sky130_fd_sc_hd__or3b_1 _3836_ (.A(\tms1x00.Y[3] ),
    .B(_0648_),
    .C_N(_1863_),
    .X(_1865_));
 sky130_fd_sc_hd__and3_1 _3837_ (.A(_1862_),
    .B(_1864_),
    .C(_1865_),
    .X(_1866_));
 sky130_fd_sc_hd__clkbuf_1 _3838_ (.A(_1866_),
    .X(_0505_));
 sky130_fd_sc_hd__or3b_1 _3839_ (.A(_0627_),
    .B(_0619_),
    .C_N(_0630_),
    .X(_1867_));
 sky130_fd_sc_hd__nor3b_1 _3840_ (.A(\tms1x00.Y[1] ),
    .B(\tms1x00.Y[0] ),
    .C_N(\tms1x00.Y[2] ),
    .Y(_1868_));
 sky130_fd_sc_hd__a31o_1 _3841_ (.A1(_0651_),
    .A2(_0656_),
    .A3(_1868_),
    .B1(net44),
    .X(_1869_));
 sky130_fd_sc_hd__o311a_1 _3842_ (.A1(_0633_),
    .A2(_0649_),
    .A3(_1867_),
    .B1(_1869_),
    .C1(_1862_),
    .X(_0506_));
 sky130_fd_sc_hd__and3b_1 _3843_ (.A_N(\tms1x00.Y[1] ),
    .B(\tms1x00.Y[0] ),
    .C(\tms1x00.Y[2] ),
    .X(_1870_));
 sky130_fd_sc_hd__a31o_1 _3844_ (.A1(_0651_),
    .A2(_0655_),
    .A3(_1870_),
    .B1(net45),
    .X(_1871_));
 sky130_fd_sc_hd__or3b_1 _3845_ (.A(\tms1x00.Y[3] ),
    .B(_0648_),
    .C_N(_1870_),
    .X(_1872_));
 sky130_fd_sc_hd__and3_1 _3846_ (.A(_1862_),
    .B(_1871_),
    .C(_1872_),
    .X(_1873_));
 sky130_fd_sc_hd__clkbuf_1 _3847_ (.A(_1873_),
    .X(_0507_));
 sky130_fd_sc_hd__and3b_1 _3848_ (.A_N(\tms1x00.Y[0] ),
    .B(\tms1x00.Y[1] ),
    .C(\tms1x00.Y[2] ),
    .X(_1874_));
 sky130_fd_sc_hd__a31o_1 _3849_ (.A1(_0650_),
    .A2(_0655_),
    .A3(_1874_),
    .B1(net46),
    .X(_1875_));
 sky130_fd_sc_hd__or3b_1 _3850_ (.A(\tms1x00.Y[3] ),
    .B(_0648_),
    .C_N(_1874_),
    .X(_1876_));
 sky130_fd_sc_hd__and3_1 _3851_ (.A(_1862_),
    .B(_1875_),
    .C(_1876_),
    .X(_1877_));
 sky130_fd_sc_hd__clkbuf_1 _3852_ (.A(_1877_),
    .X(_0508_));
 sky130_fd_sc_hd__and3_1 _3853_ (.A(\tms1x00.Y[2] ),
    .B(\tms1x00.Y[1] ),
    .C(\tms1x00.Y[0] ),
    .X(_1878_));
 sky130_fd_sc_hd__a31o_1 _3854_ (.A1(_0650_),
    .A2(_0655_),
    .A3(_1878_),
    .B1(net47),
    .X(_1879_));
 sky130_fd_sc_hd__or3b_1 _3855_ (.A(\tms1x00.Y[3] ),
    .B(_0648_),
    .C_N(_1878_),
    .X(_1880_));
 sky130_fd_sc_hd__and3_1 _3856_ (.A(_1862_),
    .B(_1879_),
    .C(_1880_),
    .X(_1881_));
 sky130_fd_sc_hd__clkbuf_1 _3857_ (.A(_1881_),
    .X(_0509_));
 sky130_fd_sc_hd__a31o_1 _3858_ (.A1(_0632_),
    .A2(_0652_),
    .A3(_0655_),
    .B1(net48),
    .X(_1882_));
 sky130_fd_sc_hd__o311a_1 _3859_ (.A1(_0651_),
    .A2(_0641_),
    .A3(_0649_),
    .B1(_1882_),
    .C1(_1862_),
    .X(_0510_));
 sky130_fd_sc_hd__a31o_1 _3860_ (.A1(_0632_),
    .A2(_0656_),
    .A3(_1857_),
    .B1(net49),
    .X(_1883_));
 sky130_fd_sc_hd__o311a_1 _3861_ (.A1(_0651_),
    .A2(_0649_),
    .A3(_1856_),
    .B1(_1883_),
    .C1(_1862_),
    .X(_0511_));
 sky130_fd_sc_hd__a31o_1 _3862_ (.A1(_0632_),
    .A2(_0656_),
    .A3(_1860_),
    .B1(net50),
    .X(_1884_));
 sky130_fd_sc_hd__o311a_1 _3863_ (.A1(_0651_),
    .A2(_0649_),
    .A3(_1859_),
    .B1(_1884_),
    .C1(_1862_),
    .X(_0512_));
 sky130_fd_sc_hd__a31o_1 _3864_ (.A1(_0632_),
    .A2(_0655_),
    .A3(_1863_),
    .B1(net51),
    .X(_1885_));
 sky130_fd_sc_hd__or3b_1 _3865_ (.A(_0650_),
    .B(_0648_),
    .C_N(_1863_),
    .X(_1886_));
 sky130_fd_sc_hd__and3_1 _3866_ (.A(_0621_),
    .B(_1885_),
    .C(_1886_),
    .X(_1887_));
 sky130_fd_sc_hd__clkbuf_1 _3867_ (.A(_1887_),
    .X(_0513_));
 sky130_fd_sc_hd__a31o_1 _3868_ (.A1(_0632_),
    .A2(_0656_),
    .A3(_1868_),
    .B1(net52),
    .X(_1888_));
 sky130_fd_sc_hd__o311a_1 _3869_ (.A1(_0651_),
    .A2(_0648_),
    .A3(_1867_),
    .B1(_1888_),
    .C1(_1862_),
    .X(_0514_));
 sky130_fd_sc_hd__nand2_1 _3870_ (.A(_0633_),
    .B(_1870_),
    .Y(_1889_));
 sky130_fd_sc_hd__a31o_1 _3871_ (.A1(_0632_),
    .A2(_0656_),
    .A3(_1870_),
    .B1(net53),
    .X(_1890_));
 sky130_fd_sc_hd__o211a_1 _3872_ (.A1(_0649_),
    .A2(_1889_),
    .B1(_1890_),
    .C1(_1843_),
    .X(_0515_));
 sky130_fd_sc_hd__nand2_1 _3873_ (.A(_0633_),
    .B(_1874_),
    .Y(_1891_));
 sky130_fd_sc_hd__a31o_1 _3874_ (.A1(_0632_),
    .A2(_0656_),
    .A3(_1874_),
    .B1(net54),
    .X(_1892_));
 sky130_fd_sc_hd__o211a_1 _3875_ (.A1(_0649_),
    .A2(_1891_),
    .B1(_1892_),
    .C1(_1843_),
    .X(_0516_));
 sky130_fd_sc_hd__nand2_1 _3876_ (.A(_0633_),
    .B(_1878_),
    .Y(_1893_));
 sky130_fd_sc_hd__a31o_1 _3877_ (.A1(_0632_),
    .A2(_0656_),
    .A3(_1878_),
    .B1(net55),
    .X(_1894_));
 sky130_fd_sc_hd__o211a_1 _3878_ (.A1(_0649_),
    .A2(_1893_),
    .B1(_1894_),
    .C1(_1843_),
    .X(_0517_));
 sky130_fd_sc_hd__nor2_1 _3879_ (.A(_0644_),
    .B(_0647_),
    .Y(_1895_));
 sky130_fd_sc_hd__and4b_1 _3880_ (.A_N(_1848_),
    .B(_1847_),
    .C(_1895_),
    .D(_0643_),
    .X(_1896_));
 sky130_fd_sc_hd__buf_2 _3881_ (.A(_1896_),
    .X(_1897_));
 sky130_fd_sc_hd__inv_2 _3882_ (.A(\tms1x00.A[0] ),
    .Y(_1898_));
 sky130_fd_sc_hd__o21ai_1 _3883_ (.A1(_0642_),
    .A2(_1898_),
    .B1(_1897_),
    .Y(_1899_));
 sky130_fd_sc_hd__o211a_1 _3884_ (.A1(net32),
    .A2(_1897_),
    .B1(_1899_),
    .C1(_1843_),
    .X(_0518_));
 sky130_fd_sc_hd__inv_2 _3885_ (.A(\tms1x00.A[1] ),
    .Y(_1900_));
 sky130_fd_sc_hd__o21ai_1 _3886_ (.A1(_0642_),
    .A2(_1900_),
    .B1(_1897_),
    .Y(_1901_));
 sky130_fd_sc_hd__o211a_1 _3887_ (.A1(net33),
    .A2(_1897_),
    .B1(_1901_),
    .C1(_1843_),
    .X(_0519_));
 sky130_fd_sc_hd__inv_2 _3888_ (.A(\tms1x00.A[2] ),
    .Y(_1902_));
 sky130_fd_sc_hd__o21ai_1 _3889_ (.A1(_0642_),
    .A2(_1902_),
    .B1(_1897_),
    .Y(_1903_));
 sky130_fd_sc_hd__o211a_1 _3890_ (.A1(net34),
    .A2(_1897_),
    .B1(_1903_),
    .C1(_1843_),
    .X(_0520_));
 sky130_fd_sc_hd__inv_2 _3891_ (.A(\tms1x00.A[3] ),
    .Y(_1904_));
 sky130_fd_sc_hd__o21ai_1 _3892_ (.A1(_0642_),
    .A2(_1904_),
    .B1(_1897_),
    .Y(_1905_));
 sky130_fd_sc_hd__o211a_1 _3893_ (.A1(net35),
    .A2(_1897_),
    .B1(_1905_),
    .C1(_1843_),
    .X(_0521_));
 sky130_fd_sc_hd__inv_2 _3894_ (.A(\tms1x00.status ),
    .Y(_1906_));
 sky130_fd_sc_hd__o21ai_1 _3895_ (.A1(_1906_),
    .A2(_0642_),
    .B1(_1897_),
    .Y(_1907_));
 sky130_fd_sc_hd__o211a_1 _3896_ (.A1(net36),
    .A2(_1897_),
    .B1(_1907_),
    .C1(_0658_),
    .X(_0522_));
 sky130_fd_sc_hd__inv_2 _3897_ (.A(\tms1x00.CL ),
    .Y(_1908_));
 sky130_fd_sc_hd__and3_1 _3898_ (.A(\tms1x00.status ),
    .B(\tms1x00.ins_in[0] ),
    .C(_1826_),
    .X(_1909_));
 sky130_fd_sc_hd__clkbuf_4 _3899_ (.A(_1909_),
    .X(_1910_));
 sky130_fd_sc_hd__nand2_2 _3900_ (.A(\tms1x00.ins_in[1] ),
    .B(_1910_),
    .Y(_1911_));
 sky130_fd_sc_hd__nor2_1 _3901_ (.A(_0646_),
    .B(_1129_),
    .Y(_1912_));
 sky130_fd_sc_hd__and3_1 _3902_ (.A(\tms1x00.CL ),
    .B(_1826_),
    .C(_1912_),
    .X(_1913_));
 sky130_fd_sc_hd__buf_2 _3903_ (.A(_1913_),
    .X(_1914_));
 sky130_fd_sc_hd__a211oi_1 _3904_ (.A1(_1908_),
    .A2(_1911_),
    .B1(_1914_),
    .C1(_1824_),
    .Y(_0523_));
 sky130_fd_sc_hd__or3_1 _3905_ (.A(\tms1x00.status ),
    .B(_1823_),
    .C(_1826_),
    .X(_1915_));
 sky130_fd_sc_hd__clkbuf_1 _3906_ (.A(_1915_),
    .X(_0524_));
 sky130_fd_sc_hd__inv_2 _3907_ (.A(_0647_),
    .Y(_1916_));
 sky130_fd_sc_hd__and3b_1 _3908_ (.A_N(\tms1x00.ins_in[2] ),
    .B(_0819_),
    .C(\tms1x00.ins_in[3] ),
    .X(_1917_));
 sky130_fd_sc_hd__nand2_1 _3909_ (.A(_1916_),
    .B(_1917_),
    .Y(_1918_));
 sky130_fd_sc_hd__mux2_1 _3910_ (.A0(\tms1x00.PA[0] ),
    .A1(\tms1x00.PB[0] ),
    .S(_1911_),
    .X(_1919_));
 sky130_fd_sc_hd__and3_1 _3911_ (.A(_1847_),
    .B(_1916_),
    .C(_1917_),
    .X(_1920_));
 sky130_fd_sc_hd__a211o_1 _3912_ (.A1(_1918_),
    .A2(_1919_),
    .B1(_1920_),
    .C1(_1824_),
    .X(_0525_));
 sky130_fd_sc_hd__mux2_1 _3913_ (.A0(\tms1x00.PA[1] ),
    .A1(\tms1x00.PB[1] ),
    .S(_1911_),
    .X(_1921_));
 sky130_fd_sc_hd__and3_1 _3914_ (.A(_1848_),
    .B(_1916_),
    .C(_1917_),
    .X(_1922_));
 sky130_fd_sc_hd__a211o_1 _3915_ (.A1(_1918_),
    .A2(_1921_),
    .B1(_1922_),
    .C1(_1824_),
    .X(_0526_));
 sky130_fd_sc_hd__mux2_1 _3916_ (.A0(\tms1x00.PA[2] ),
    .A1(\tms1x00.PB[2] ),
    .S(_1911_),
    .X(_1923_));
 sky130_fd_sc_hd__mux2_1 _3917_ (.A0(_0643_),
    .A1(_1923_),
    .S(_1918_),
    .X(_1924_));
 sky130_fd_sc_hd__or2_1 _3918_ (.A(_1823_),
    .B(_1924_),
    .X(_1925_));
 sky130_fd_sc_hd__clkbuf_1 _3919_ (.A(_1925_),
    .X(_0527_));
 sky130_fd_sc_hd__mux2_1 _3920_ (.A0(\tms1x00.PA[3] ),
    .A1(\tms1x00.PB[3] ),
    .S(_1911_),
    .X(_1926_));
 sky130_fd_sc_hd__mux2_1 _3921_ (.A0(_0642_),
    .A1(_1926_),
    .S(_1918_),
    .X(_1927_));
 sky130_fd_sc_hd__or2_1 _3922_ (.A(_1823_),
    .B(_1927_),
    .X(_1928_));
 sky130_fd_sc_hd__clkbuf_1 _3923_ (.A(_1928_),
    .X(_0528_));
 sky130_fd_sc_hd__and4_2 _3924_ (.A(_1908_),
    .B(\tms1x00.ins_in[1] ),
    .C(_0621_),
    .D(_1910_),
    .X(_1929_));
 sky130_fd_sc_hd__mux2_1 _3925_ (.A0(\tms1x00.SR[0] ),
    .A1(\tms1x00.PC[0] ),
    .S(_1929_),
    .X(_1930_));
 sky130_fd_sc_hd__clkbuf_1 _3926_ (.A(_1930_),
    .X(_0529_));
 sky130_fd_sc_hd__mux2_1 _3927_ (.A0(\tms1x00.SR[1] ),
    .A1(\tms1x00.PC[1] ),
    .S(_1929_),
    .X(_1931_));
 sky130_fd_sc_hd__clkbuf_1 _3928_ (.A(_1931_),
    .X(_0530_));
 sky130_fd_sc_hd__mux2_1 _3929_ (.A0(\tms1x00.SR[2] ),
    .A1(\tms1x00.PC[2] ),
    .S(_1929_),
    .X(_1932_));
 sky130_fd_sc_hd__clkbuf_1 _3930_ (.A(_1932_),
    .X(_0531_));
 sky130_fd_sc_hd__mux2_1 _3931_ (.A0(\tms1x00.SR[3] ),
    .A1(\tms1x00.PC[3] ),
    .S(_1929_),
    .X(_1933_));
 sky130_fd_sc_hd__clkbuf_1 _3932_ (.A(_1933_),
    .X(_0532_));
 sky130_fd_sc_hd__mux2_1 _3933_ (.A0(\tms1x00.SR[4] ),
    .A1(\tms1x00.PC[4] ),
    .S(_1929_),
    .X(_1934_));
 sky130_fd_sc_hd__clkbuf_1 _3934_ (.A(_1934_),
    .X(_0533_));
 sky130_fd_sc_hd__mux2_1 _3935_ (.A0(\tms1x00.SR[5] ),
    .A1(\tms1x00.PC[5] ),
    .S(_1929_),
    .X(_1935_));
 sky130_fd_sc_hd__clkbuf_1 _3936_ (.A(_1935_),
    .X(_0534_));
 sky130_fd_sc_hd__and3_1 _3937_ (.A(\tms1x00.status ),
    .B(_1908_),
    .C(\tms1x00.ins_in[0] ),
    .X(_1936_));
 sky130_fd_sc_hd__o21a_1 _3938_ (.A1(_1912_),
    .A2(_1936_),
    .B1(_1826_),
    .X(_1937_));
 sky130_fd_sc_hd__mux2_1 _3939_ (.A0(\tms1x00.PA[0] ),
    .A1(\tms1x00.PB[0] ),
    .S(_1937_),
    .X(_1938_));
 sky130_fd_sc_hd__or2_1 _3940_ (.A(_1823_),
    .B(_1938_),
    .X(_1939_));
 sky130_fd_sc_hd__clkbuf_1 _3941_ (.A(_1939_),
    .X(_0535_));
 sky130_fd_sc_hd__mux2_1 _3942_ (.A0(\tms1x00.PA[1] ),
    .A1(\tms1x00.PB[1] ),
    .S(_1937_),
    .X(_1940_));
 sky130_fd_sc_hd__or2_1 _3943_ (.A(_1823_),
    .B(_1940_),
    .X(_1941_));
 sky130_fd_sc_hd__clkbuf_1 _3944_ (.A(_1941_),
    .X(_0536_));
 sky130_fd_sc_hd__mux2_1 _3945_ (.A0(\tms1x00.PA[2] ),
    .A1(\tms1x00.PB[2] ),
    .S(_1937_),
    .X(_1942_));
 sky130_fd_sc_hd__or2_1 _3946_ (.A(_1823_),
    .B(_1942_),
    .X(_1943_));
 sky130_fd_sc_hd__clkbuf_1 _3947_ (.A(_1943_),
    .X(_0537_));
 sky130_fd_sc_hd__mux2_1 _3948_ (.A0(\tms1x00.PA[3] ),
    .A1(\tms1x00.PB[3] ),
    .S(_1937_),
    .X(_1944_));
 sky130_fd_sc_hd__or2_1 _3949_ (.A(_1823_),
    .B(_1944_),
    .X(_1945_));
 sky130_fd_sc_hd__clkbuf_1 _3950_ (.A(_1945_),
    .X(_0538_));
 sky130_fd_sc_hd__inv_2 _3951_ (.A(_1910_),
    .Y(_1946_));
 sky130_fd_sc_hd__inv_2 _3952_ (.A(_1914_),
    .Y(_1947_));
 sky130_fd_sc_hd__or3_1 _3953_ (.A(\tms1x00.PC[0] ),
    .B(_1910_),
    .C(_1914_),
    .X(_1948_));
 sky130_fd_sc_hd__o221a_1 _3954_ (.A1(\tms1x00.ins_in[2] ),
    .A2(_1946_),
    .B1(_1947_),
    .B2(\tms1x00.SR[0] ),
    .C1(_1948_),
    .X(_1949_));
 sky130_fd_sc_hd__a21oi_1 _3955_ (.A1(_0623_),
    .A2(_1949_),
    .B1(_1824_),
    .Y(_1950_));
 sky130_fd_sc_hd__o21a_1 _3956_ (.A1(_0623_),
    .A2(_1949_),
    .B1(_1950_),
    .X(_0539_));
 sky130_fd_sc_hd__nor2_1 _3957_ (.A(_1910_),
    .B(_1914_),
    .Y(_1951_));
 sky130_fd_sc_hd__and2_1 _3958_ (.A(\tms1x00.PC[1] ),
    .B(_1951_),
    .X(_1952_));
 sky130_fd_sc_hd__a22o_1 _3959_ (.A1(\tms1x00.ins_in[3] ),
    .A2(_1910_),
    .B1(_1914_),
    .B2(\tms1x00.SR[1] ),
    .X(_1953_));
 sky130_fd_sc_hd__o21a_1 _3960_ (.A1(_1952_),
    .A2(_1953_),
    .B1(_1840_),
    .X(_0540_));
 sky130_fd_sc_hd__and2_1 _3961_ (.A(\tms1x00.PC[2] ),
    .B(_1951_),
    .X(_1954_));
 sky130_fd_sc_hd__a22o_1 _3962_ (.A1(_1847_),
    .A2(_1910_),
    .B1(_1914_),
    .B2(\tms1x00.SR[2] ),
    .X(_1955_));
 sky130_fd_sc_hd__o21a_1 _3963_ (.A1(_1954_),
    .A2(_1955_),
    .B1(_1840_),
    .X(_0541_));
 sky130_fd_sc_hd__and2_1 _3964_ (.A(\tms1x00.PC[3] ),
    .B(_1951_),
    .X(_1956_));
 sky130_fd_sc_hd__a22o_1 _3965_ (.A1(_1848_),
    .A2(_1910_),
    .B1(_1914_),
    .B2(\tms1x00.SR[3] ),
    .X(_1957_));
 sky130_fd_sc_hd__o21a_1 _3966_ (.A1(_1956_),
    .A2(_1957_),
    .B1(_1840_),
    .X(_0542_));
 sky130_fd_sc_hd__and2_1 _3967_ (.A(\tms1x00.PC[4] ),
    .B(_1951_),
    .X(_1958_));
 sky130_fd_sc_hd__a22o_1 _3968_ (.A1(_0643_),
    .A2(_1910_),
    .B1(_1914_),
    .B2(\tms1x00.SR[4] ),
    .X(_1959_));
 sky130_fd_sc_hd__o21a_1 _3969_ (.A1(_1958_),
    .A2(_1959_),
    .B1(_1840_),
    .X(_0543_));
 sky130_fd_sc_hd__and2_1 _3970_ (.A(\tms1x00.PC[5] ),
    .B(_1951_),
    .X(_1960_));
 sky130_fd_sc_hd__a22o_1 _3971_ (.A1(_0642_),
    .A2(_1910_),
    .B1(_1914_),
    .B2(\tms1x00.SR[5] ),
    .X(_1961_));
 sky130_fd_sc_hd__o21a_1 _3972_ (.A1(_1960_),
    .A2(_1961_),
    .B1(_1840_),
    .X(_0544_));
 sky130_fd_sc_hd__or3_1 _3973_ (.A(net39),
    .B(net38),
    .C(net16),
    .X(_1962_));
 sky130_fd_sc_hd__nor2_2 _3974_ (.A(net37),
    .B(_1962_),
    .Y(_1963_));
 sky130_fd_sc_hd__and2_1 _3975_ (.A(_0659_),
    .B(_1917_),
    .X(_1964_));
 sky130_fd_sc_hd__nor3_1 _3976_ (.A(_0764_),
    .B(_0817_),
    .C(_1964_),
    .Y(_1965_));
 sky130_fd_sc_hd__nand2_1 _3977_ (.A(\tms1x00.ins_in[1] ),
    .B(\tms1x00.ins_in[0] ),
    .Y(_1966_));
 sky130_fd_sc_hd__or2_1 _3978_ (.A(_0660_),
    .B(_1966_),
    .X(_1967_));
 sky130_fd_sc_hd__nor4_1 _3979_ (.A(\tms1x00.ins_in[7] ),
    .B(_0643_),
    .C(_1848_),
    .D(_1847_),
    .Y(_1968_));
 sky130_fd_sc_hd__and2_1 _3980_ (.A(\tms1x00.ins_in[3] ),
    .B(_1968_),
    .X(_1969_));
 sky130_fd_sc_hd__or2_1 _3981_ (.A(net37),
    .B(_1962_),
    .X(_1970_));
 sky130_fd_sc_hd__a221o_1 _3982_ (.A1(_1847_),
    .A2(_0930_),
    .B1(_1969_),
    .B2(\tms1x00.K_latch[0] ),
    .C1(_1970_),
    .X(_1971_));
 sky130_fd_sc_hd__a21o_1 _3983_ (.A1(_0619_),
    .A2(_1967_),
    .B1(_1971_),
    .X(_1972_));
 sky130_fd_sc_hd__o22a_1 _3984_ (.A1(\tms1x00.P[0] ),
    .A2(_1963_),
    .B1(_1965_),
    .B2(_1972_),
    .X(_0545_));
 sky130_fd_sc_hd__nor3_1 _3985_ (.A(_0882_),
    .B(_0929_),
    .C(_1964_),
    .Y(_1973_));
 sky130_fd_sc_hd__a221o_1 _3986_ (.A1(_1848_),
    .A2(_0930_),
    .B1(_1969_),
    .B2(\tms1x00.K_latch[1] ),
    .C1(_1970_),
    .X(_1974_));
 sky130_fd_sc_hd__a21o_1 _3987_ (.A1(_0627_),
    .A2(_1967_),
    .B1(_1974_),
    .X(_1975_));
 sky130_fd_sc_hd__o22a_1 _3988_ (.A1(\tms1x00.P[1] ),
    .A2(_1963_),
    .B1(_1973_),
    .B2(_1975_),
    .X(_0546_));
 sky130_fd_sc_hd__nor2_1 _3989_ (.A(_0983_),
    .B(_1030_),
    .Y(_1976_));
 sky130_fd_sc_hd__nand2_1 _3990_ (.A(_0659_),
    .B(_1917_),
    .Y(_1977_));
 sky130_fd_sc_hd__a221o_1 _3991_ (.A1(\tms1x00.Y[2] ),
    .A2(_1967_),
    .B1(_1969_),
    .B2(\tms1x00.K_latch[2] ),
    .C1(_0930_),
    .X(_1978_));
 sky130_fd_sc_hd__a211o_1 _3992_ (.A1(_1976_),
    .A2(_1977_),
    .B1(_1978_),
    .C1(_1970_),
    .X(_1979_));
 sky130_fd_sc_hd__o21a_1 _3993_ (.A1(\tms1x00.P[2] ),
    .A2(_1963_),
    .B1(_1979_),
    .X(_0547_));
 sky130_fd_sc_hd__and2_1 _3994_ (.A(_1128_),
    .B(_1977_),
    .X(_1980_));
 sky130_fd_sc_hd__a221o_1 _3995_ (.A1(_0632_),
    .A2(_1967_),
    .B1(_1969_),
    .B2(\tms1x00.K_latch[3] ),
    .C1(_1970_),
    .X(_1981_));
 sky130_fd_sc_hd__o22a_1 _3996_ (.A1(\tms1x00.P[3] ),
    .A2(_1963_),
    .B1(_1980_),
    .B2(_1981_),
    .X(_0548_));
 sky130_fd_sc_hd__nor3b_4 _3997_ (.A(_1847_),
    .B(_0654_),
    .C_N(_1848_),
    .Y(_1982_));
 sky130_fd_sc_hd__o31a_1 _3998_ (.A1(\tms1x00.ins_in[5] ),
    .A2(_1847_),
    .A3(_0653_),
    .B1(\tms1x00.N[0] ),
    .X(_1983_));
 sky130_fd_sc_hd__or4_1 _3999_ (.A(\tms1x00.ins_in[5] ),
    .B(\tms1x00.ins_in[4] ),
    .C(\tms1x00.N[0] ),
    .D(_0653_),
    .X(_1984_));
 sky130_fd_sc_hd__and2b_1 _4000_ (.A_N(_1983_),
    .B(_1984_),
    .X(_1985_));
 sky130_fd_sc_hd__xnor2_1 _4001_ (.A(\tms1x00.P[0] ),
    .B(_1985_),
    .Y(_1986_));
 sky130_fd_sc_hd__nand2_1 _4002_ (.A(_1982_),
    .B(_1986_),
    .Y(_1987_));
 sky130_fd_sc_hd__o211a_1 _4003_ (.A1(_0619_),
    .A2(_1982_),
    .B1(_1987_),
    .C1(_0658_),
    .X(_0549_));
 sky130_fd_sc_hd__and2_1 _4004_ (.A(\tms1x00.P[1] ),
    .B(\tms1x00.N[1] ),
    .X(_1988_));
 sky130_fd_sc_hd__nor2_1 _4005_ (.A(\tms1x00.P[1] ),
    .B(\tms1x00.N[1] ),
    .Y(_1989_));
 sky130_fd_sc_hd__or2_1 _4006_ (.A(_1988_),
    .B(_1989_),
    .X(_1990_));
 sky130_fd_sc_hd__a21oi_1 _4007_ (.A1(\tms1x00.P[0] ),
    .A2(_1984_),
    .B1(_1983_),
    .Y(_1991_));
 sky130_fd_sc_hd__xnor2_1 _4008_ (.A(_1990_),
    .B(_1991_),
    .Y(_1992_));
 sky130_fd_sc_hd__nand2_1 _4009_ (.A(_1982_),
    .B(_1992_),
    .Y(_1993_));
 sky130_fd_sc_hd__o211a_1 _4010_ (.A1(_0627_),
    .A2(_1982_),
    .B1(_1993_),
    .C1(_0658_),
    .X(_0550_));
 sky130_fd_sc_hd__nand2_1 _4011_ (.A(\tms1x00.P[2] ),
    .B(\tms1x00.N[2] ),
    .Y(_1994_));
 sky130_fd_sc_hd__or2_1 _4012_ (.A(\tms1x00.P[2] ),
    .B(\tms1x00.N[2] ),
    .X(_1995_));
 sky130_fd_sc_hd__nand2_1 _4013_ (.A(_1994_),
    .B(_1995_),
    .Y(_1996_));
 sky130_fd_sc_hd__o21ba_1 _4014_ (.A1(_1989_),
    .A2(_1991_),
    .B1_N(_1988_),
    .X(_1997_));
 sky130_fd_sc_hd__xnor2_1 _4015_ (.A(_1996_),
    .B(_1997_),
    .Y(_1998_));
 sky130_fd_sc_hd__nand2_1 _4016_ (.A(_1982_),
    .B(_1998_),
    .Y(_1999_));
 sky130_fd_sc_hd__o211a_1 _4017_ (.A1(_0630_),
    .A2(_1982_),
    .B1(_1999_),
    .C1(_0658_),
    .X(_0551_));
 sky130_fd_sc_hd__o21a_1 _4018_ (.A1(_1996_),
    .A2(_1997_),
    .B1(_1994_),
    .X(_2000_));
 sky130_fd_sc_hd__xnor2_1 _4019_ (.A(\tms1x00.P[3] ),
    .B(\tms1x00.N[3] ),
    .Y(_2001_));
 sky130_fd_sc_hd__xnor2_1 _4020_ (.A(_2000_),
    .B(_2001_),
    .Y(_2002_));
 sky130_fd_sc_hd__nand2_1 _4021_ (.A(_1982_),
    .B(_2002_),
    .Y(_2003_));
 sky130_fd_sc_hd__o211a_1 _4022_ (.A1(_0633_),
    .A2(_1982_),
    .B1(_2003_),
    .C1(_0658_),
    .X(_0552_));
 sky130_fd_sc_hd__and3_1 _4023_ (.A(_1848_),
    .B(_1847_),
    .C(_0820_),
    .X(_2004_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _4024_ (.A(_2004_),
    .X(_2005_));
 sky130_fd_sc_hd__a22o_1 _4025_ (.A1(_1895_),
    .A2(_1968_),
    .B1(_2005_),
    .B2(_1916_),
    .X(_2006_));
 sky130_fd_sc_hd__nand2_1 _4026_ (.A(_0643_),
    .B(_2005_),
    .Y(_2007_));
 sky130_fd_sc_hd__o211ai_1 _4027_ (.A1(\tms1x00.X[0] ),
    .A2(_2005_),
    .B1(_2006_),
    .C1(_2007_),
    .Y(_2008_));
 sky130_fd_sc_hd__o211a_1 _4028_ (.A1(\tms1x00.X[0] ),
    .A2(_2006_),
    .B1(_2008_),
    .C1(_0658_),
    .X(_0553_));
 sky130_fd_sc_hd__nand2_1 _4029_ (.A(_0642_),
    .B(_2005_),
    .Y(_2009_));
 sky130_fd_sc_hd__o211ai_1 _4030_ (.A1(\tms1x00.X[1] ),
    .A2(_2005_),
    .B1(_2006_),
    .C1(_2009_),
    .Y(_2010_));
 sky130_fd_sc_hd__o211a_1 _4031_ (.A1(\tms1x00.X[1] ),
    .A2(_2006_),
    .B1(_2010_),
    .C1(_0658_),
    .X(_0554_));
 sky130_fd_sc_hd__o21ai_1 _4032_ (.A1(\tms1x00.X[2] ),
    .A2(_1848_),
    .B1(_2006_),
    .Y(_2011_));
 sky130_fd_sc_hd__o211a_1 _4033_ (.A1(\tms1x00.X[2] ),
    .A2(_2006_),
    .B1(_2011_),
    .C1(_0658_),
    .X(_0555_));
 sky130_fd_sc_hd__or2_1 _4034_ (.A(\tms1x00.N[0] ),
    .B(_1963_),
    .X(_2012_));
 sky130_fd_sc_hd__clkbuf_1 _4035_ (.A(_2012_),
    .X(_0556_));
 sky130_fd_sc_hd__or2_1 _4036_ (.A(\tms1x00.N[1] ),
    .B(_1963_),
    .X(_2013_));
 sky130_fd_sc_hd__clkbuf_1 _4037_ (.A(_2013_),
    .X(_0557_));
 sky130_fd_sc_hd__or2_1 _4038_ (.A(\tms1x00.N[2] ),
    .B(_1963_),
    .X(_2014_));
 sky130_fd_sc_hd__clkbuf_1 _4039_ (.A(_2014_),
    .X(_0558_));
 sky130_fd_sc_hd__or2_1 _4040_ (.A(\tms1x00.N[3] ),
    .B(_1963_),
    .X(_2015_));
 sky130_fd_sc_hd__clkbuf_1 _4041_ (.A(_2015_),
    .X(_0559_));
 sky130_fd_sc_hd__or4b_1 _4042_ (.A(_1848_),
    .B(net16),
    .C(_0654_),
    .D_N(_1847_),
    .X(_2016_));
 sky130_fd_sc_hd__buf_2 _4043_ (.A(_2016_),
    .X(_2017_));
 sky130_fd_sc_hd__nand2_1 _4044_ (.A(\tms1x00.A[0] ),
    .B(_2017_),
    .Y(_2018_));
 sky130_fd_sc_hd__o21ai_1 _4045_ (.A1(_1986_),
    .A2(_2017_),
    .B1(_2018_),
    .Y(_0560_));
 sky130_fd_sc_hd__nand2_1 _4046_ (.A(\tms1x00.A[1] ),
    .B(_2017_),
    .Y(_2019_));
 sky130_fd_sc_hd__o21ai_1 _4047_ (.A1(_1992_),
    .A2(_2017_),
    .B1(_2019_),
    .Y(_0561_));
 sky130_fd_sc_hd__nand2_1 _4048_ (.A(\tms1x00.A[2] ),
    .B(_2017_),
    .Y(_2020_));
 sky130_fd_sc_hd__o21ai_1 _4049_ (.A1(_1998_),
    .A2(_2017_),
    .B1(_2020_),
    .Y(_0562_));
 sky130_fd_sc_hd__nand2_1 _4050_ (.A(\tms1x00.A[3] ),
    .B(_2017_),
    .Y(_2021_));
 sky130_fd_sc_hd__o21ai_1 _4051_ (.A1(_2002_),
    .A2(_2017_),
    .B1(_2021_),
    .Y(_0563_));
 sky130_fd_sc_hd__nor3_4 _4052_ (.A(_0635_),
    .B(_0637_),
    .C(_0639_),
    .Y(_2022_));
 sky130_fd_sc_hd__nand2_2 _4053_ (.A(_1162_),
    .B(_2022_),
    .Y(_2023_));
 sky130_fd_sc_hd__mux2_1 _4054_ (.A0(_1797_),
    .A1(\tms1x00.RAM[13][0] ),
    .S(_2023_),
    .X(_2024_));
 sky130_fd_sc_hd__clkbuf_1 _4055_ (.A(_2024_),
    .X(_0564_));
 sky130_fd_sc_hd__mux2_1 _4056_ (.A0(_1800_),
    .A1(\tms1x00.RAM[13][1] ),
    .S(_2023_),
    .X(_2025_));
 sky130_fd_sc_hd__clkbuf_1 _4057_ (.A(_2025_),
    .X(_0565_));
 sky130_fd_sc_hd__mux2_1 _4058_ (.A0(_1802_),
    .A1(\tms1x00.RAM[13][2] ),
    .S(_2023_),
    .X(_2026_));
 sky130_fd_sc_hd__clkbuf_1 _4059_ (.A(_2026_),
    .X(_0566_));
 sky130_fd_sc_hd__mux2_1 _4060_ (.A0(_1804_),
    .A1(\tms1x00.RAM[13][3] ),
    .S(_2023_),
    .X(_2027_));
 sky130_fd_sc_hd__clkbuf_1 _4061_ (.A(_2027_),
    .X(_0567_));
 sky130_fd_sc_hd__or2_2 _4062_ (.A(_1460_),
    .B(_1320_),
    .X(_2028_));
 sky130_fd_sc_hd__mux2_1 _4063_ (.A0(_1797_),
    .A1(\tms1x00.RAM[18][0] ),
    .S(_2028_),
    .X(_2029_));
 sky130_fd_sc_hd__clkbuf_1 _4064_ (.A(_2029_),
    .X(_0568_));
 sky130_fd_sc_hd__mux2_1 _4065_ (.A0(_1800_),
    .A1(\tms1x00.RAM[18][1] ),
    .S(_2028_),
    .X(_2030_));
 sky130_fd_sc_hd__clkbuf_1 _4066_ (.A(_2030_),
    .X(_0569_));
 sky130_fd_sc_hd__mux2_1 _4067_ (.A0(_1802_),
    .A1(\tms1x00.RAM[18][2] ),
    .S(_2028_),
    .X(_2031_));
 sky130_fd_sc_hd__clkbuf_1 _4068_ (.A(_2031_),
    .X(_0570_));
 sky130_fd_sc_hd__mux2_1 _4069_ (.A0(_1804_),
    .A1(\tms1x00.RAM[18][3] ),
    .S(_2028_),
    .X(_2032_));
 sky130_fd_sc_hd__clkbuf_1 _4070_ (.A(_2032_),
    .X(_0571_));
 sky130_fd_sc_hd__nor2_2 _4071_ (.A(_1257_),
    .B(_1508_),
    .Y(_2033_));
 sky130_fd_sc_hd__mux2_1 _4072_ (.A0(\tms1x00.RAM[39][0] ),
    .A1(_1263_),
    .S(_2033_),
    .X(_2034_));
 sky130_fd_sc_hd__clkbuf_1 _4073_ (.A(_2034_),
    .X(_0572_));
 sky130_fd_sc_hd__mux2_1 _4074_ (.A0(\tms1x00.RAM[39][1] ),
    .A1(_1269_),
    .S(_2033_),
    .X(_2035_));
 sky130_fd_sc_hd__clkbuf_1 _4075_ (.A(_2035_),
    .X(_0573_));
 sky130_fd_sc_hd__mux2_1 _4076_ (.A0(\tms1x00.RAM[39][2] ),
    .A1(_1272_),
    .S(_2033_),
    .X(_2036_));
 sky130_fd_sc_hd__clkbuf_1 _4077_ (.A(_2036_),
    .X(_0574_));
 sky130_fd_sc_hd__mux2_1 _4078_ (.A0(\tms1x00.RAM[39][3] ),
    .A1(_1275_),
    .S(_2033_),
    .X(_2037_));
 sky130_fd_sc_hd__clkbuf_1 _4079_ (.A(_2037_),
    .X(_0575_));
 sky130_fd_sc_hd__nand2_2 _4080_ (.A(_1213_),
    .B(_2022_),
    .Y(_2038_));
 sky130_fd_sc_hd__mux2_1 _4081_ (.A0(_1797_),
    .A1(\tms1x00.RAM[14][0] ),
    .S(_2038_),
    .X(_2039_));
 sky130_fd_sc_hd__clkbuf_1 _4082_ (.A(_2039_),
    .X(_0576_));
 sky130_fd_sc_hd__mux2_1 _4083_ (.A0(_1800_),
    .A1(\tms1x00.RAM[14][1] ),
    .S(_2038_),
    .X(_2040_));
 sky130_fd_sc_hd__clkbuf_1 _4084_ (.A(_2040_),
    .X(_0577_));
 sky130_fd_sc_hd__mux2_1 _4085_ (.A0(_1802_),
    .A1(\tms1x00.RAM[14][2] ),
    .S(_2038_),
    .X(_2041_));
 sky130_fd_sc_hd__clkbuf_1 _4086_ (.A(_2041_),
    .X(_0578_));
 sky130_fd_sc_hd__mux2_1 _4087_ (.A0(_1804_),
    .A1(\tms1x00.RAM[14][3] ),
    .S(_2038_),
    .X(_2042_));
 sky130_fd_sc_hd__clkbuf_1 _4088_ (.A(_2042_),
    .X(_0579_));
 sky130_fd_sc_hd__or2_2 _4089_ (.A(_1194_),
    .B(_1200_),
    .X(_2043_));
 sky130_fd_sc_hd__mux2_1 _4090_ (.A0(_1797_),
    .A1(\tms1x00.RAM[17][0] ),
    .S(_2043_),
    .X(_2044_));
 sky130_fd_sc_hd__clkbuf_1 _4091_ (.A(_2044_),
    .X(_0580_));
 sky130_fd_sc_hd__mux2_1 _4092_ (.A0(_1800_),
    .A1(\tms1x00.RAM[17][1] ),
    .S(_2043_),
    .X(_2045_));
 sky130_fd_sc_hd__clkbuf_1 _4093_ (.A(_2045_),
    .X(_0581_));
 sky130_fd_sc_hd__mux2_1 _4094_ (.A0(_1802_),
    .A1(\tms1x00.RAM[17][2] ),
    .S(_2043_),
    .X(_2046_));
 sky130_fd_sc_hd__clkbuf_1 _4095_ (.A(_2046_),
    .X(_0582_));
 sky130_fd_sc_hd__mux2_1 _4096_ (.A0(_1804_),
    .A1(\tms1x00.RAM[17][3] ),
    .S(_2043_),
    .X(_2047_));
 sky130_fd_sc_hd__clkbuf_1 _4097_ (.A(_2047_),
    .X(_0583_));
 sky130_fd_sc_hd__nand2_2 _4098_ (.A(_1162_),
    .B(_1481_),
    .Y(_2048_));
 sky130_fd_sc_hd__mux2_1 _4099_ (.A0(_1797_),
    .A1(\tms1x00.RAM[29][0] ),
    .S(_2048_),
    .X(_2049_));
 sky130_fd_sc_hd__clkbuf_1 _4100_ (.A(_2049_),
    .X(_0584_));
 sky130_fd_sc_hd__mux2_1 _4101_ (.A0(_1800_),
    .A1(\tms1x00.RAM[29][1] ),
    .S(_2048_),
    .X(_2050_));
 sky130_fd_sc_hd__clkbuf_1 _4102_ (.A(_2050_),
    .X(_0585_));
 sky130_fd_sc_hd__mux2_1 _4103_ (.A0(_1802_),
    .A1(\tms1x00.RAM[29][2] ),
    .S(_2048_),
    .X(_2051_));
 sky130_fd_sc_hd__clkbuf_1 _4104_ (.A(_2051_),
    .X(_0586_));
 sky130_fd_sc_hd__mux2_1 _4105_ (.A0(_1804_),
    .A1(\tms1x00.RAM[29][3] ),
    .S(_2048_),
    .X(_2052_));
 sky130_fd_sc_hd__clkbuf_1 _4106_ (.A(_2052_),
    .X(_0587_));
 sky130_fd_sc_hd__or2_2 _4107_ (.A(_1460_),
    .B(_1311_),
    .X(_2053_));
 sky130_fd_sc_hd__mux2_1 _4108_ (.A0(_1797_),
    .A1(\tms1x00.RAM[16][0] ),
    .S(_2053_),
    .X(_2054_));
 sky130_fd_sc_hd__clkbuf_1 _4109_ (.A(_2054_),
    .X(_0588_));
 sky130_fd_sc_hd__mux2_1 _4110_ (.A0(_1800_),
    .A1(\tms1x00.RAM[16][1] ),
    .S(_2053_),
    .X(_2055_));
 sky130_fd_sc_hd__clkbuf_1 _4111_ (.A(_2055_),
    .X(_0589_));
 sky130_fd_sc_hd__mux2_1 _4112_ (.A0(_1802_),
    .A1(\tms1x00.RAM[16][2] ),
    .S(_2053_),
    .X(_2056_));
 sky130_fd_sc_hd__clkbuf_1 _4113_ (.A(_2056_),
    .X(_0590_));
 sky130_fd_sc_hd__mux2_1 _4114_ (.A0(_1804_),
    .A1(\tms1x00.RAM[16][3] ),
    .S(_2053_),
    .X(_2057_));
 sky130_fd_sc_hd__clkbuf_1 _4115_ (.A(_2057_),
    .X(_0591_));
 sky130_fd_sc_hd__or2_2 _4116_ (.A(_1337_),
    .B(_1257_),
    .X(_2058_));
 sky130_fd_sc_hd__mux2_1 _4117_ (.A0(_1797_),
    .A1(\tms1x00.RAM[119][0] ),
    .S(_2058_),
    .X(_2059_));
 sky130_fd_sc_hd__clkbuf_1 _4118_ (.A(_2059_),
    .X(_0592_));
 sky130_fd_sc_hd__mux2_1 _4119_ (.A0(_1800_),
    .A1(\tms1x00.RAM[119][1] ),
    .S(_2058_),
    .X(_2060_));
 sky130_fd_sc_hd__clkbuf_1 _4120_ (.A(_2060_),
    .X(_0593_));
 sky130_fd_sc_hd__mux2_1 _4121_ (.A0(_1802_),
    .A1(\tms1x00.RAM[119][2] ),
    .S(_2058_),
    .X(_2061_));
 sky130_fd_sc_hd__clkbuf_1 _4122_ (.A(_2061_),
    .X(_0594_));
 sky130_fd_sc_hd__mux2_1 _4123_ (.A0(_1804_),
    .A1(\tms1x00.RAM[119][3] ),
    .S(_2058_),
    .X(_2062_));
 sky130_fd_sc_hd__clkbuf_1 _4124_ (.A(_2062_),
    .X(_0595_));
 sky130_fd_sc_hd__nand2_2 _4125_ (.A(_1224_),
    .B(_2022_),
    .Y(_2063_));
 sky130_fd_sc_hd__mux2_1 _4126_ (.A0(_1135_),
    .A1(\tms1x00.RAM[12][0] ),
    .S(_2063_),
    .X(_2064_));
 sky130_fd_sc_hd__clkbuf_1 _4127_ (.A(_2064_),
    .X(_0596_));
 sky130_fd_sc_hd__mux2_1 _4128_ (.A0(_1143_),
    .A1(\tms1x00.RAM[12][1] ),
    .S(_2063_),
    .X(_2065_));
 sky130_fd_sc_hd__clkbuf_1 _4129_ (.A(_2065_),
    .X(_0597_));
 sky130_fd_sc_hd__mux2_1 _4130_ (.A0(_1145_),
    .A1(\tms1x00.RAM[12][2] ),
    .S(_2063_),
    .X(_2066_));
 sky130_fd_sc_hd__clkbuf_1 _4131_ (.A(_2066_),
    .X(_0598_));
 sky130_fd_sc_hd__mux2_1 _4132_ (.A0(_1147_),
    .A1(\tms1x00.RAM[12][3] ),
    .S(_2063_),
    .X(_2067_));
 sky130_fd_sc_hd__clkbuf_1 _4133_ (.A(_2067_),
    .X(_0599_));
 sky130_fd_sc_hd__nand2_2 _4134_ (.A(_1170_),
    .B(_2022_),
    .Y(_2068_));
 sky130_fd_sc_hd__mux2_1 _4135_ (.A0(_1135_),
    .A1(\tms1x00.RAM[15][0] ),
    .S(_2068_),
    .X(_2069_));
 sky130_fd_sc_hd__clkbuf_1 _4136_ (.A(_2069_),
    .X(_0600_));
 sky130_fd_sc_hd__mux2_1 _4137_ (.A0(_1143_),
    .A1(\tms1x00.RAM[15][1] ),
    .S(_2068_),
    .X(_2070_));
 sky130_fd_sc_hd__clkbuf_1 _4138_ (.A(_2070_),
    .X(_0601_));
 sky130_fd_sc_hd__mux2_1 _4139_ (.A0(_1145_),
    .A1(\tms1x00.RAM[15][2] ),
    .S(_2068_),
    .X(_2071_));
 sky130_fd_sc_hd__clkbuf_1 _4140_ (.A(_2071_),
    .X(_0602_));
 sky130_fd_sc_hd__mux2_1 _4141_ (.A0(_1147_),
    .A1(\tms1x00.RAM[15][3] ),
    .S(_2068_),
    .X(_2072_));
 sky130_fd_sc_hd__clkbuf_1 _4142_ (.A(_2072_),
    .X(_0603_));
 sky130_fd_sc_hd__buf_4 _4143_ (.A(_1962_),
    .X(_2073_));
 sky130_fd_sc_hd__mux2_1 _4144_ (.A0(\tms1x00.PC[0] ),
    .A1(\tms1x00.rom_addr[0] ),
    .S(_2073_),
    .X(_2074_));
 sky130_fd_sc_hd__clkbuf_1 _4145_ (.A(_2074_),
    .X(_0604_));
 sky130_fd_sc_hd__mux2_1 _4146_ (.A0(\tms1x00.PC[1] ),
    .A1(_1827_),
    .S(_2073_),
    .X(_2075_));
 sky130_fd_sc_hd__clkbuf_1 _4147_ (.A(_2075_),
    .X(_0605_));
 sky130_fd_sc_hd__mux2_1 _4148_ (.A0(\tms1x00.PC[2] ),
    .A1(net57),
    .S(_2073_),
    .X(_2076_));
 sky130_fd_sc_hd__clkbuf_1 _4149_ (.A(_2076_),
    .X(_0606_));
 sky130_fd_sc_hd__mux2_1 _4150_ (.A0(\tms1x00.PC[3] ),
    .A1(net58),
    .S(_2073_),
    .X(_2077_));
 sky130_fd_sc_hd__clkbuf_1 _4151_ (.A(_2077_),
    .X(_0607_));
 sky130_fd_sc_hd__mux2_1 _4152_ (.A0(\tms1x00.PC[4] ),
    .A1(net59),
    .S(_2073_),
    .X(_2078_));
 sky130_fd_sc_hd__clkbuf_1 _4153_ (.A(_2078_),
    .X(_0608_));
 sky130_fd_sc_hd__mux2_1 _4154_ (.A0(\tms1x00.PC[5] ),
    .A1(net60),
    .S(_2073_),
    .X(_2079_));
 sky130_fd_sc_hd__clkbuf_1 _4155_ (.A(_2079_),
    .X(_0609_));
 sky130_fd_sc_hd__mux2_1 _4156_ (.A0(\tms1x00.PA[0] ),
    .A1(net61),
    .S(_2073_),
    .X(_2080_));
 sky130_fd_sc_hd__clkbuf_1 _4157_ (.A(_2080_),
    .X(_0610_));
 sky130_fd_sc_hd__mux2_1 _4158_ (.A0(\tms1x00.PA[1] ),
    .A1(net62),
    .S(_2073_),
    .X(_2081_));
 sky130_fd_sc_hd__clkbuf_1 _4159_ (.A(_2081_),
    .X(_0611_));
 sky130_fd_sc_hd__mux2_1 _4160_ (.A0(\tms1x00.PA[2] ),
    .A1(net63),
    .S(_2073_),
    .X(_2082_));
 sky130_fd_sc_hd__clkbuf_1 _4161_ (.A(_2082_),
    .X(_0612_));
 sky130_fd_sc_hd__mux2_1 _4162_ (.A0(\tms1x00.PA[3] ),
    .A1(net64),
    .S(_2073_),
    .X(_2083_));
 sky130_fd_sc_hd__clkbuf_1 _4163_ (.A(_2083_),
    .X(_0613_));
 sky130_fd_sc_hd__nor2_2 _4164_ (.A(_1140_),
    .B(_1243_),
    .Y(_2084_));
 sky130_fd_sc_hd__mux2_1 _4165_ (.A0(\tms1x00.RAM[9][0] ),
    .A1(_1263_),
    .S(_2084_),
    .X(_2085_));
 sky130_fd_sc_hd__clkbuf_1 _4166_ (.A(_2085_),
    .X(_0614_));
 sky130_fd_sc_hd__mux2_1 _4167_ (.A0(\tms1x00.RAM[9][1] ),
    .A1(_1269_),
    .S(_2084_),
    .X(_2086_));
 sky130_fd_sc_hd__clkbuf_1 _4168_ (.A(_2086_),
    .X(_0615_));
 sky130_fd_sc_hd__mux2_1 _4169_ (.A0(\tms1x00.RAM[9][2] ),
    .A1(_1272_),
    .S(_2084_),
    .X(_2087_));
 sky130_fd_sc_hd__clkbuf_1 _4170_ (.A(_2087_),
    .X(_0616_));
 sky130_fd_sc_hd__mux2_1 _4171_ (.A0(\tms1x00.RAM[9][3] ),
    .A1(_1275_),
    .S(_2084_),
    .X(_2088_));
 sky130_fd_sc_hd__clkbuf_1 _4172_ (.A(_2088_),
    .X(_0617_));
 sky130_fd_sc_hd__dfxtp_1 _4173_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0015_),
    .Q(net40));
 sky130_fd_sc_hd__dfxtp_1 _4174_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_0000_),
    .Q(net77));
 sky130_fd_sc_hd__dfxtp_1 _4175_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0016_),
    .Q(\tms1x00.RAM[99][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4176_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0017_),
    .Q(\tms1x00.RAM[99][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4177_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0018_),
    .Q(\tms1x00.RAM[99][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4178_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0019_),
    .Q(\tms1x00.RAM[99][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4179_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0020_),
    .Q(\tms1x00.RAM[89][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4180_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0021_),
    .Q(\tms1x00.RAM[89][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4181_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0022_),
    .Q(\tms1x00.RAM[89][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4182_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0023_),
    .Q(\tms1x00.RAM[89][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4183_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0024_),
    .Q(\tms1x00.RAM[59][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4184_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0025_),
    .Q(\tms1x00.RAM[59][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4185_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0026_),
    .Q(\tms1x00.RAM[59][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4186_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0027_),
    .Q(\tms1x00.RAM[59][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4187_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0028_),
    .Q(\tms1x00.RAM[109][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4188_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0029_),
    .Q(\tms1x00.RAM[109][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4189_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0030_),
    .Q(\tms1x00.RAM[109][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4190_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0031_),
    .Q(\tms1x00.RAM[109][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4191_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0032_),
    .Q(\tms1x00.RAM[79][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4192_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0033_),
    .Q(\tms1x00.RAM[79][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4193_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0034_),
    .Q(\tms1x00.RAM[79][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4194_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0035_),
    .Q(\tms1x00.RAM[79][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4195_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0036_),
    .Q(\tms1x00.RAM[69][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4196_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0037_),
    .Q(\tms1x00.RAM[69][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4197_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0038_),
    .Q(\tms1x00.RAM[69][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4198_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0039_),
    .Q(\tms1x00.RAM[69][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4199_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0040_),
    .Q(\tms1x00.RAM[127][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4200_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0041_),
    .Q(\tms1x00.RAM[127][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4201_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0042_),
    .Q(\tms1x00.RAM[127][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4202_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0043_),
    .Q(\tms1x00.RAM[127][3] ));
 sky130_fd_sc_hd__dfxtp_4 _4203_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_0044_),
    .Q(net56));
 sky130_fd_sc_hd__dfxtp_1 _4204_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0045_),
    .Q(\tms1x00.RAM[49][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4205_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0046_),
    .Q(\tms1x00.RAM[49][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4206_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0047_),
    .Q(\tms1x00.RAM[49][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4207_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0048_),
    .Q(\tms1x00.RAM[49][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4208_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0049_),
    .Q(\tms1x00.RAM[19][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4209_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0050_),
    .Q(\tms1x00.RAM[19][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4210_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0051_),
    .Q(\tms1x00.RAM[19][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4211_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0052_),
    .Q(\tms1x00.RAM[19][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4212_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0053_),
    .Q(\tms1x00.RAM[95][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4213_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0054_),
    .Q(\tms1x00.RAM[95][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4214_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0055_),
    .Q(\tms1x00.RAM[95][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4215_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0056_),
    .Q(\tms1x00.RAM[95][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4216_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0057_),
    .Q(\tms1x00.RAM[94][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4217_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0058_),
    .Q(\tms1x00.RAM[94][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4218_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0059_),
    .Q(\tms1x00.RAM[94][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4219_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0060_),
    .Q(\tms1x00.RAM[94][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4220_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0061_),
    .Q(\tms1x00.RAM[93][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4221_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0062_),
    .Q(\tms1x00.RAM[93][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4222_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0063_),
    .Q(\tms1x00.RAM[93][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4223_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0064_),
    .Q(\tms1x00.RAM[93][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4224_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0065_),
    .Q(\tms1x00.RAM[92][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4225_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0066_),
    .Q(\tms1x00.RAM[92][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4226_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0067_),
    .Q(\tms1x00.RAM[92][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4227_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0068_),
    .Q(\tms1x00.RAM[92][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4228_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0069_),
    .Q(\tms1x00.RAM[91][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4229_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0070_),
    .Q(\tms1x00.RAM[91][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4230_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0071_),
    .Q(\tms1x00.RAM[91][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4231_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0072_),
    .Q(\tms1x00.RAM[91][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4232_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0073_),
    .Q(\tms1x00.RAM[90][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4233_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0074_),
    .Q(\tms1x00.RAM[90][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4234_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0075_),
    .Q(\tms1x00.RAM[90][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4235_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0076_),
    .Q(\tms1x00.RAM[90][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4236_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0077_),
    .Q(\tms1x00.RAM[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4237_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0078_),
    .Q(\tms1x00.RAM[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4238_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0079_),
    .Q(\tms1x00.RAM[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4239_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0080_),
    .Q(\tms1x00.RAM[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4240_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0081_),
    .Q(\tms1x00.RAM[88][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4241_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0082_),
    .Q(\tms1x00.RAM[88][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4242_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0083_),
    .Q(\tms1x00.RAM[88][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4243_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0084_),
    .Q(\tms1x00.RAM[88][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4244_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0085_),
    .Q(\tms1x00.RAM[87][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4245_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0086_),
    .Q(\tms1x00.RAM[87][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4246_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0087_),
    .Q(\tms1x00.RAM[87][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4247_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0088_),
    .Q(\tms1x00.RAM[87][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4248_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_0089_),
    .Q(\tms1x00.RAM[86][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4249_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0090_),
    .Q(\tms1x00.RAM[86][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4250_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_0091_),
    .Q(\tms1x00.RAM[86][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4251_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_0092_),
    .Q(\tms1x00.RAM[86][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4252_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0093_),
    .Q(\tms1x00.RAM[105][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4253_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0094_),
    .Q(\tms1x00.RAM[105][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4254_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0095_),
    .Q(\tms1x00.RAM[105][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4255_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0096_),
    .Q(\tms1x00.RAM[105][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4256_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_0097_),
    .Q(\tms1x00.RAM[104][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4257_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0098_),
    .Q(\tms1x00.RAM[104][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4258_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0099_),
    .Q(\tms1x00.RAM[104][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4259_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0100_),
    .Q(\tms1x00.RAM[104][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4260_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_0101_),
    .Q(\tms1x00.RAM[103][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4261_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_0102_),
    .Q(\tms1x00.RAM[103][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4262_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_0103_),
    .Q(\tms1x00.RAM[103][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4263_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_0104_),
    .Q(\tms1x00.RAM[103][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4264_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_0105_),
    .Q(\tms1x00.RAM[102][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4265_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_0106_),
    .Q(\tms1x00.RAM[102][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4266_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_0107_),
    .Q(\tms1x00.RAM[102][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4267_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_0108_),
    .Q(\tms1x00.RAM[102][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4268_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_0109_),
    .Q(\tms1x00.RAM[101][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4269_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_0110_),
    .Q(\tms1x00.RAM[101][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4270_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_0111_),
    .Q(\tms1x00.RAM[101][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4271_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_0112_),
    .Q(\tms1x00.RAM[101][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4272_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_0113_),
    .Q(\tms1x00.RAM[100][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4273_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_0114_),
    .Q(\tms1x00.RAM[100][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4274_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_0115_),
    .Q(\tms1x00.RAM[100][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4275_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_0116_),
    .Q(\tms1x00.RAM[100][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4276_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0117_),
    .Q(\tms1x00.RAM[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4277_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0118_),
    .Q(\tms1x00.RAM[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4278_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0119_),
    .Q(\tms1x00.RAM[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4279_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0120_),
    .Q(\tms1x00.RAM[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4280_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0121_),
    .Q(\tms1x00.RAM[98][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4281_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0122_),
    .Q(\tms1x00.RAM[98][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4282_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0123_),
    .Q(\tms1x00.RAM[98][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4283_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0124_),
    .Q(\tms1x00.RAM[98][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4284_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0125_),
    .Q(\tms1x00.RAM[97][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4285_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0126_),
    .Q(\tms1x00.RAM[97][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4286_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0127_),
    .Q(\tms1x00.RAM[97][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4287_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0128_),
    .Q(\tms1x00.RAM[97][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4288_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0129_),
    .Q(\tms1x00.RAM[96][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4289_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0130_),
    .Q(\tms1x00.RAM[96][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4290_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0131_),
    .Q(\tms1x00.RAM[96][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4291_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0132_),
    .Q(\tms1x00.RAM[96][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4292_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0133_),
    .Q(\tms1x00.RAM[115][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4293_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0134_),
    .Q(\tms1x00.RAM[115][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4294_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0135_),
    .Q(\tms1x00.RAM[115][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4295_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0136_),
    .Q(\tms1x00.RAM[115][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4296_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0137_),
    .Q(\tms1x00.RAM[114][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4297_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0138_),
    .Q(\tms1x00.RAM[114][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4298_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0139_),
    .Q(\tms1x00.RAM[114][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4299_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0140_),
    .Q(\tms1x00.RAM[114][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4300_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0141_),
    .Q(\tms1x00.RAM[113][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4301_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0142_),
    .Q(\tms1x00.RAM[113][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4302_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0143_),
    .Q(\tms1x00.RAM[113][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4303_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0144_),
    .Q(\tms1x00.RAM[113][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4304_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0145_),
    .Q(\tms1x00.RAM[112][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4305_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0146_),
    .Q(\tms1x00.RAM[112][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4306_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0147_),
    .Q(\tms1x00.RAM[112][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4307_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0148_),
    .Q(\tms1x00.RAM[112][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4308_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0149_),
    .Q(\tms1x00.RAM[111][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4309_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0150_),
    .Q(\tms1x00.RAM[111][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4310_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0151_),
    .Q(\tms1x00.RAM[111][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4311_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0152_),
    .Q(\tms1x00.RAM[111][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4312_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0153_),
    .Q(\tms1x00.RAM[110][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4313_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0154_),
    .Q(\tms1x00.RAM[110][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4314_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0155_),
    .Q(\tms1x00.RAM[110][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4315_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0156_),
    .Q(\tms1x00.RAM[110][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4316_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0157_),
    .Q(\tms1x00.RAM[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4317_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0158_),
    .Q(\tms1x00.RAM[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4318_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0159_),
    .Q(\tms1x00.RAM[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4319_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0160_),
    .Q(\tms1x00.RAM[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4320_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0161_),
    .Q(\tms1x00.RAM[108][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4321_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0162_),
    .Q(\tms1x00.RAM[108][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4322_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0163_),
    .Q(\tms1x00.RAM[108][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4323_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0164_),
    .Q(\tms1x00.RAM[108][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4324_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_0165_),
    .Q(\tms1x00.RAM[107][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4325_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_0166_),
    .Q(\tms1x00.RAM[107][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4326_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0167_),
    .Q(\tms1x00.RAM[107][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4327_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_0168_),
    .Q(\tms1x00.RAM[107][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4328_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_0169_),
    .Q(\tms1x00.RAM[106][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4329_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0170_),
    .Q(\tms1x00.RAM[106][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4330_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_0171_),
    .Q(\tms1x00.RAM[106][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4331_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_0172_),
    .Q(\tms1x00.RAM[106][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4332_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0173_),
    .Q(\tms1x00.RAM[125][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4333_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0174_),
    .Q(\tms1x00.RAM[125][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4334_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0175_),
    .Q(\tms1x00.RAM[125][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4335_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0176_),
    .Q(\tms1x00.RAM[125][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4336_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0177_),
    .Q(\tms1x00.RAM[124][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4337_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0178_),
    .Q(\tms1x00.RAM[124][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4338_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0179_),
    .Q(\tms1x00.RAM[124][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4339_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0180_),
    .Q(\tms1x00.RAM[124][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4340_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0181_),
    .Q(\tms1x00.RAM[123][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4341_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0182_),
    .Q(\tms1x00.RAM[123][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4342_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0183_),
    .Q(\tms1x00.RAM[123][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4343_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0184_),
    .Q(\tms1x00.RAM[123][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4344_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0185_),
    .Q(\tms1x00.RAM[122][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4345_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0186_),
    .Q(\tms1x00.RAM[122][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4346_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0187_),
    .Q(\tms1x00.RAM[122][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4347_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0188_),
    .Q(\tms1x00.RAM[122][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4348_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0189_),
    .Q(\tms1x00.RAM[121][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4349_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0190_),
    .Q(\tms1x00.RAM[121][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4350_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0191_),
    .Q(\tms1x00.RAM[121][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4351_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0192_),
    .Q(\tms1x00.RAM[121][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4352_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0193_),
    .Q(\tms1x00.RAM[120][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4353_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0194_),
    .Q(\tms1x00.RAM[120][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4354_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0195_),
    .Q(\tms1x00.RAM[120][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4355_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0196_),
    .Q(\tms1x00.RAM[120][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4356_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0197_),
    .Q(\tms1x00.RAM[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4357_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0198_),
    .Q(\tms1x00.RAM[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4358_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0199_),
    .Q(\tms1x00.RAM[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4359_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0200_),
    .Q(\tms1x00.RAM[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4360_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0201_),
    .Q(\tms1x00.RAM[118][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4361_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0202_),
    .Q(\tms1x00.RAM[118][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4362_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0203_),
    .Q(\tms1x00.RAM[118][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4363_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0204_),
    .Q(\tms1x00.RAM[118][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4364_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0205_),
    .Q(\tms1x00.RAM[117][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4365_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0206_),
    .Q(\tms1x00.RAM[117][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4366_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0207_),
    .Q(\tms1x00.RAM[117][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4367_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0208_),
    .Q(\tms1x00.RAM[117][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4368_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0209_),
    .Q(\tms1x00.RAM[116][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4369_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0210_),
    .Q(\tms1x00.RAM[116][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4370_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0211_),
    .Q(\tms1x00.RAM[116][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4371_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0212_),
    .Q(\tms1x00.RAM[116][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4372_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0213_),
    .Q(\tms1x00.RAM[126][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4373_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0214_),
    .Q(\tms1x00.RAM[126][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4374_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0215_),
    .Q(\tms1x00.RAM[126][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4375_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0216_),
    .Q(\tms1x00.RAM[126][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4376_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0217_),
    .Q(\tms1x00.RAM[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4377_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0218_),
    .Q(\tms1x00.RAM[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4378_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0219_),
    .Q(\tms1x00.RAM[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4379_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0220_),
    .Q(\tms1x00.RAM[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4380_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0221_),
    .Q(\tms1x00.RAM[23][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4381_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0222_),
    .Q(\tms1x00.RAM[23][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4382_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0223_),
    .Q(\tms1x00.RAM[23][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4383_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0224_),
    .Q(\tms1x00.RAM[23][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4384_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0225_),
    .Q(\tms1x00.RAM[22][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4385_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0226_),
    .Q(\tms1x00.RAM[22][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4386_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0227_),
    .Q(\tms1x00.RAM[22][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4387_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0228_),
    .Q(\tms1x00.RAM[22][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4388_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0229_),
    .Q(\tms1x00.RAM[21][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4389_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0230_),
    .Q(\tms1x00.RAM[21][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4390_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0231_),
    .Q(\tms1x00.RAM[21][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4391_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0232_),
    .Q(\tms1x00.RAM[21][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4392_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0233_),
    .Q(\tms1x00.RAM[20][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4393_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0234_),
    .Q(\tms1x00.RAM[20][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4394_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0235_),
    .Q(\tms1x00.RAM[20][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4395_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0236_),
    .Q(\tms1x00.RAM[20][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4396_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0237_),
    .Q(\tms1x00.RAM[28][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4397_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0238_),
    .Q(\tms1x00.RAM[28][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4398_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0239_),
    .Q(\tms1x00.RAM[28][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4399_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0240_),
    .Q(\tms1x00.RAM[28][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4400_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0241_),
    .Q(\tms1x00.RAM[27][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4401_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0242_),
    .Q(\tms1x00.RAM[27][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4402_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0243_),
    .Q(\tms1x00.RAM[27][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4403_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0244_),
    .Q(\tms1x00.RAM[27][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4404_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0245_),
    .Q(\tms1x00.RAM[26][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4405_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0246_),
    .Q(\tms1x00.RAM[26][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4406_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0247_),
    .Q(\tms1x00.RAM[26][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4407_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0248_),
    .Q(\tms1x00.RAM[26][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4408_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0249_),
    .Q(\tms1x00.RAM[25][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4409_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0250_),
    .Q(\tms1x00.RAM[25][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4410_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0251_),
    .Q(\tms1x00.RAM[25][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4411_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0252_),
    .Q(\tms1x00.RAM[25][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4412_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0253_),
    .Q(\tms1x00.RAM[24][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4413_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0254_),
    .Q(\tms1x00.RAM[24][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4414_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0255_),
    .Q(\tms1x00.RAM[24][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4415_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0256_),
    .Q(\tms1x00.RAM[24][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4416_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0257_),
    .Q(\tms1x00.RAM[32][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4417_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0258_),
    .Q(\tms1x00.RAM[32][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4418_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0259_),
    .Q(\tms1x00.RAM[32][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4419_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0260_),
    .Q(\tms1x00.RAM[32][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4420_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0261_),
    .Q(\tms1x00.RAM[31][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4421_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0262_),
    .Q(\tms1x00.RAM[31][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4422_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0263_),
    .Q(\tms1x00.RAM[31][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4423_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0264_),
    .Q(\tms1x00.RAM[31][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4424_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0265_),
    .Q(\tms1x00.RAM[30][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4425_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0266_),
    .Q(\tms1x00.RAM[30][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4426_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0267_),
    .Q(\tms1x00.RAM[30][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4427_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0268_),
    .Q(\tms1x00.RAM[30][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4428_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0269_),
    .Q(\tms1x00.RAM[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4429_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0270_),
    .Q(\tms1x00.RAM[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4430_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0271_),
    .Q(\tms1x00.RAM[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4431_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0272_),
    .Q(\tms1x00.RAM[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4432_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0273_),
    .Q(\tms1x00.RAM[36][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4433_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0274_),
    .Q(\tms1x00.RAM[36][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4434_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_0275_),
    .Q(\tms1x00.RAM[36][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4435_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_0276_),
    .Q(\tms1x00.RAM[36][3] ));
 sky130_fd_sc_hd__dfxtp_2 _4436_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0008_),
    .Q(_0001_));
 sky130_fd_sc_hd__dfxtp_4 _4437_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0009_),
    .Q(_0002_));
 sky130_fd_sc_hd__dfxtp_2 _4438_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0010_),
    .Q(_0003_));
 sky130_fd_sc_hd__dfxtp_2 _4439_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0011_),
    .Q(_0004_));
 sky130_fd_sc_hd__dfxtp_2 _4440_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0012_),
    .Q(_0005_));
 sky130_fd_sc_hd__dfxtp_1 _4441_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0013_),
    .Q(_0006_));
 sky130_fd_sc_hd__dfxtp_2 _4442_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0014_),
    .Q(_0007_));
 sky130_fd_sc_hd__dfxtp_1 _4443_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0277_),
    .Q(\tms1x00.RAM[35][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4444_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0278_),
    .Q(\tms1x00.RAM[35][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4445_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0279_),
    .Q(\tms1x00.RAM[35][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4446_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0280_),
    .Q(\tms1x00.RAM[35][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4447_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0281_),
    .Q(\tms1x00.RAM[34][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4448_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0282_),
    .Q(\tms1x00.RAM[34][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4449_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0283_),
    .Q(\tms1x00.RAM[34][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4450_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0284_),
    .Q(\tms1x00.RAM[34][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4451_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0285_),
    .Q(\tms1x00.RAM[33][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4452_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0286_),
    .Q(\tms1x00.RAM[33][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4453_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0287_),
    .Q(\tms1x00.RAM[33][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4454_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0288_),
    .Q(\tms1x00.RAM[33][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4455_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0289_),
    .Q(\tms1x00.RAM[41][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4456_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0290_),
    .Q(\tms1x00.RAM[41][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4457_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0291_),
    .Q(\tms1x00.RAM[41][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4458_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0292_),
    .Q(\tms1x00.RAM[41][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4459_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0293_),
    .Q(\tms1x00.RAM[40][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4460_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0294_),
    .Q(\tms1x00.RAM[40][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4461_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0295_),
    .Q(\tms1x00.RAM[40][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4462_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0296_),
    .Q(\tms1x00.RAM[40][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4463_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0297_),
    .Q(\tms1x00.RAM[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4464_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0298_),
    .Q(\tms1x00.RAM[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4465_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0299_),
    .Q(\tms1x00.RAM[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4466_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0300_),
    .Q(\tms1x00.RAM[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4467_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0301_),
    .Q(\tms1x00.RAM[38][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4468_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0302_),
    .Q(\tms1x00.RAM[38][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4469_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0303_),
    .Q(\tms1x00.RAM[38][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4470_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0304_),
    .Q(\tms1x00.RAM[38][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4471_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0305_),
    .Q(\tms1x00.RAM[37][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4472_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0306_),
    .Q(\tms1x00.RAM[37][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4473_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0307_),
    .Q(\tms1x00.RAM[37][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4474_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0308_),
    .Q(\tms1x00.RAM[37][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4475_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0309_),
    .Q(\tms1x00.RAM[45][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4476_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0310_),
    .Q(\tms1x00.RAM[45][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4477_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0311_),
    .Q(\tms1x00.RAM[45][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4478_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0312_),
    .Q(\tms1x00.RAM[45][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4479_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0313_),
    .Q(\tms1x00.RAM[44][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4480_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0314_),
    .Q(\tms1x00.RAM[44][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4481_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0315_),
    .Q(\tms1x00.RAM[44][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4482_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0316_),
    .Q(\tms1x00.RAM[44][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4483_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0317_),
    .Q(\tms1x00.RAM[43][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4484_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0318_),
    .Q(\tms1x00.RAM[43][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4485_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0319_),
    .Q(\tms1x00.RAM[43][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4486_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0320_),
    .Q(\tms1x00.RAM[43][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4487_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0321_),
    .Q(\tms1x00.RAM[42][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4488_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0322_),
    .Q(\tms1x00.RAM[42][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4489_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0323_),
    .Q(\tms1x00.RAM[42][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4490_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0324_),
    .Q(\tms1x00.RAM[42][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4491_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0325_),
    .Q(\tms1x00.RAM[50][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4492_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0326_),
    .Q(\tms1x00.RAM[50][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4493_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0327_),
    .Q(\tms1x00.RAM[50][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4494_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0328_),
    .Q(\tms1x00.RAM[50][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4495_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0329_),
    .Q(\tms1x00.RAM[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4496_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0330_),
    .Q(\tms1x00.RAM[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4497_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0331_),
    .Q(\tms1x00.RAM[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4498_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0332_),
    .Q(\tms1x00.RAM[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4499_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0333_),
    .Q(\tms1x00.RAM[48][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4500_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0334_),
    .Q(\tms1x00.RAM[48][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4501_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0335_),
    .Q(\tms1x00.RAM[48][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4502_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0336_),
    .Q(\tms1x00.RAM[48][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4503_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0337_),
    .Q(\tms1x00.RAM[47][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4504_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0338_),
    .Q(\tms1x00.RAM[47][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4505_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0339_),
    .Q(\tms1x00.RAM[47][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4506_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0340_),
    .Q(\tms1x00.RAM[47][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4507_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0341_),
    .Q(\tms1x00.RAM[46][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4508_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0342_),
    .Q(\tms1x00.RAM[46][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4509_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0343_),
    .Q(\tms1x00.RAM[46][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4510_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0344_),
    .Q(\tms1x00.RAM[46][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4511_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0345_),
    .Q(\tms1x00.RAM[54][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4512_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0346_),
    .Q(\tms1x00.RAM[54][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4513_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0347_),
    .Q(\tms1x00.RAM[54][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4514_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0348_),
    .Q(\tms1x00.RAM[54][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4515_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0349_),
    .Q(\tms1x00.RAM[53][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4516_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0350_),
    .Q(\tms1x00.RAM[53][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4517_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0351_),
    .Q(\tms1x00.RAM[53][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4518_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0352_),
    .Q(\tms1x00.RAM[53][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4519_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0353_),
    .Q(\tms1x00.RAM[52][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4520_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0354_),
    .Q(\tms1x00.RAM[52][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4521_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0355_),
    .Q(\tms1x00.RAM[52][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4522_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0356_),
    .Q(\tms1x00.RAM[52][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4523_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0357_),
    .Q(\tms1x00.RAM[51][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4524_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0358_),
    .Q(\tms1x00.RAM[51][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4525_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0359_),
    .Q(\tms1x00.RAM[51][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4526_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0360_),
    .Q(\tms1x00.RAM[51][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4527_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0361_),
    .Q(\tms1x00.RAM[58][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4528_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0362_),
    .Q(\tms1x00.RAM[58][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4529_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0363_),
    .Q(\tms1x00.RAM[58][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4530_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0364_),
    .Q(\tms1x00.RAM[58][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4531_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0365_),
    .Q(\tms1x00.RAM[57][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4532_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0366_),
    .Q(\tms1x00.RAM[57][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4533_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0367_),
    .Q(\tms1x00.RAM[57][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4534_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0368_),
    .Q(\tms1x00.RAM[57][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4535_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0369_),
    .Q(\tms1x00.RAM[56][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4536_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0370_),
    .Q(\tms1x00.RAM[56][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4537_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0371_),
    .Q(\tms1x00.RAM[56][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4538_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0372_),
    .Q(\tms1x00.RAM[56][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4539_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0373_),
    .Q(\tms1x00.RAM[55][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4540_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0374_),
    .Q(\tms1x00.RAM[55][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4541_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0375_),
    .Q(\tms1x00.RAM[55][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4542_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0376_),
    .Q(\tms1x00.RAM[55][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4543_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0377_),
    .Q(\tms1x00.RAM[63][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4544_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0378_),
    .Q(\tms1x00.RAM[63][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4545_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0379_),
    .Q(\tms1x00.RAM[63][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4546_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0380_),
    .Q(\tms1x00.RAM[63][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4547_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0381_),
    .Q(\tms1x00.RAM[62][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4548_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0382_),
    .Q(\tms1x00.RAM[62][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4549_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0383_),
    .Q(\tms1x00.RAM[62][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4550_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0384_),
    .Q(\tms1x00.RAM[62][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4551_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0385_),
    .Q(\tms1x00.RAM[61][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4552_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0386_),
    .Q(\tms1x00.RAM[61][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4553_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0387_),
    .Q(\tms1x00.RAM[61][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4554_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0388_),
    .Q(\tms1x00.RAM[61][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4555_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0389_),
    .Q(\tms1x00.RAM[60][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4556_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0390_),
    .Q(\tms1x00.RAM[60][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4557_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0391_),
    .Q(\tms1x00.RAM[60][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4558_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0392_),
    .Q(\tms1x00.RAM[60][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4559_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0393_),
    .Q(\tms1x00.RAM[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4560_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0394_),
    .Q(\tms1x00.RAM[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4561_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0395_),
    .Q(\tms1x00.RAM[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4562_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0396_),
    .Q(\tms1x00.RAM[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4563_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0397_),
    .Q(\tms1x00.RAM[67][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4564_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0398_),
    .Q(\tms1x00.RAM[67][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4565_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0399_),
    .Q(\tms1x00.RAM[67][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4566_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0400_),
    .Q(\tms1x00.RAM[67][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4567_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0401_),
    .Q(\tms1x00.RAM[66][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4568_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0402_),
    .Q(\tms1x00.RAM[66][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4569_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0403_),
    .Q(\tms1x00.RAM[66][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4570_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0404_),
    .Q(\tms1x00.RAM[66][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4571_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0405_),
    .Q(\tms1x00.RAM[65][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4572_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0406_),
    .Q(\tms1x00.RAM[65][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4573_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0407_),
    .Q(\tms1x00.RAM[65][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4574_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0408_),
    .Q(\tms1x00.RAM[65][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4575_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0409_),
    .Q(\tms1x00.RAM[64][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4576_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0410_),
    .Q(\tms1x00.RAM[64][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4577_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0411_),
    .Q(\tms1x00.RAM[64][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4578_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0412_),
    .Q(\tms1x00.RAM[64][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4579_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0413_),
    .Q(\tms1x00.RAM[71][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4580_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0414_),
    .Q(\tms1x00.RAM[71][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4581_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0415_),
    .Q(\tms1x00.RAM[71][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4582_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0416_),
    .Q(\tms1x00.RAM[71][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4583_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0417_),
    .Q(\tms1x00.RAM[70][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4584_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0418_),
    .Q(\tms1x00.RAM[70][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4585_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0419_),
    .Q(\tms1x00.RAM[70][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4586_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0420_),
    .Q(\tms1x00.RAM[70][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4587_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0421_),
    .Q(\tms1x00.RAM[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4588_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0422_),
    .Q(\tms1x00.RAM[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4589_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0423_),
    .Q(\tms1x00.RAM[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4590_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0424_),
    .Q(\tms1x00.RAM[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4591_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0425_),
    .Q(\tms1x00.RAM[68][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4592_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0426_),
    .Q(\tms1x00.RAM[68][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4593_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0427_),
    .Q(\tms1x00.RAM[68][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4594_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0428_),
    .Q(\tms1x00.RAM[68][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4595_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0429_),
    .Q(\tms1x00.RAM[76][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4596_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0430_),
    .Q(\tms1x00.RAM[76][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4597_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0431_),
    .Q(\tms1x00.RAM[76][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4598_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0432_),
    .Q(\tms1x00.RAM[76][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4599_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0433_),
    .Q(\tms1x00.RAM[75][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4600_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_0434_),
    .Q(\tms1x00.RAM[75][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4601_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0435_),
    .Q(\tms1x00.RAM[75][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4602_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_0436_),
    .Q(\tms1x00.RAM[75][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4603_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0437_),
    .Q(\tms1x00.RAM[74][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4604_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_0438_),
    .Q(\tms1x00.RAM[74][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4605_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0439_),
    .Q(\tms1x00.RAM[74][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4606_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_0440_),
    .Q(\tms1x00.RAM[74][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4607_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0441_),
    .Q(\tms1x00.RAM[73][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4608_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0442_),
    .Q(\tms1x00.RAM[73][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4609_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_0443_),
    .Q(\tms1x00.RAM[73][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4610_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_0444_),
    .Q(\tms1x00.RAM[73][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4611_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_0445_),
    .Q(\tms1x00.RAM[72][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4612_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_0446_),
    .Q(\tms1x00.RAM[72][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4613_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_0447_),
    .Q(\tms1x00.RAM[72][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4614_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_0448_),
    .Q(\tms1x00.RAM[72][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4615_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0449_),
    .Q(\tms1x00.RAM[77][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4616_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0450_),
    .Q(\tms1x00.RAM[77][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4617_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0451_),
    .Q(\tms1x00.RAM[77][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4618_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0452_),
    .Q(\tms1x00.RAM[77][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4619_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0453_),
    .Q(\tms1x00.RAM[80][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4620_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0454_),
    .Q(\tms1x00.RAM[80][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4621_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0455_),
    .Q(\tms1x00.RAM[80][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4622_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0456_),
    .Q(\tms1x00.RAM[80][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4623_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0457_),
    .Q(\tms1x00.RAM[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4624_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0458_),
    .Q(\tms1x00.RAM[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4625_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0459_),
    .Q(\tms1x00.RAM[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4626_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0460_),
    .Q(\tms1x00.RAM[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4627_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0461_),
    .Q(\tms1x00.RAM[78][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4628_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0462_),
    .Q(\tms1x00.RAM[78][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4629_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0463_),
    .Q(\tms1x00.RAM[78][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4630_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0464_),
    .Q(\tms1x00.RAM[78][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4631_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_0465_),
    .Q(\tms1x00.RAM[85][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4632_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0466_),
    .Q(\tms1x00.RAM[85][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4633_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0467_),
    .Q(\tms1x00.RAM[85][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4634_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0468_),
    .Q(\tms1x00.RAM[85][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4635_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0469_),
    .Q(\tms1x00.RAM[84][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4636_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0470_),
    .Q(\tms1x00.RAM[84][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4637_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0471_),
    .Q(\tms1x00.RAM[84][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4638_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_0472_),
    .Q(\tms1x00.RAM[84][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4639_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0473_),
    .Q(\tms1x00.RAM[83][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4640_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0474_),
    .Q(\tms1x00.RAM[83][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4641_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0475_),
    .Q(\tms1x00.RAM[83][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4642_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0476_),
    .Q(\tms1x00.RAM[83][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4643_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0477_),
    .Q(\tms1x00.RAM[82][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4644_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0478_),
    .Q(\tms1x00.RAM[82][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4645_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0479_),
    .Q(\tms1x00.RAM[82][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4646_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0480_),
    .Q(\tms1x00.RAM[82][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4647_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0481_),
    .Q(\tms1x00.RAM[81][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4648_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0482_),
    .Q(\tms1x00.RAM[81][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4649_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0483_),
    .Q(\tms1x00.RAM[81][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4650_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0484_),
    .Q(\tms1x00.RAM[81][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4651_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0485_),
    .Q(\tms1x00.ram_addr_buff[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4652_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0486_),
    .Q(\tms1x00.ram_addr_buff[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4653_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0487_),
    .Q(\tms1x00.ram_addr_buff[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4654_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0488_),
    .Q(\tms1x00.ram_addr_buff[3] ));
 sky130_fd_sc_hd__dfxtp_2 _4655_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0489_),
    .Q(\tms1x00.ram_addr_buff[4] ));
 sky130_fd_sc_hd__dfxtp_2 _4656_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0490_),
    .Q(\tms1x00.ram_addr_buff[5] ));
 sky130_fd_sc_hd__dfxtp_2 _4657_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0491_),
    .Q(\tms1x00.ram_addr_buff[6] ));
 sky130_fd_sc_hd__dfxtp_4 _4658_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0492_),
    .Q(net37));
 sky130_fd_sc_hd__dfxtp_4 _4659_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0493_),
    .Q(net38));
 sky130_fd_sc_hd__dfxtp_2 _4660_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0494_),
    .Q(net39));
 sky130_fd_sc_hd__dfxtp_1 _4661_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0495_),
    .Q(\tms1x00.ins_in[0] ));
 sky130_fd_sc_hd__dfxtp_2 _4662_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0496_),
    .Q(\tms1x00.ins_in[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4663_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0497_),
    .Q(\tms1x00.ins_in[2] ));
 sky130_fd_sc_hd__dfxtp_2 _4664_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0498_),
    .Q(\tms1x00.ins_in[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4665_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0499_),
    .Q(\tms1x00.ins_in[4] ));
 sky130_fd_sc_hd__dfxtp_2 _4666_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0500_),
    .Q(\tms1x00.ins_in[5] ));
 sky130_fd_sc_hd__dfxtp_1 _4667_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0501_),
    .Q(\tms1x00.ins_in[6] ));
 sky130_fd_sc_hd__dfxtp_2 _4668_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0502_),
    .Q(\tms1x00.ins_in[7] ));
 sky130_fd_sc_hd__dfxtp_1 _4669_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net1),
    .Q(\tms1x00.K_latch[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4670_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net2),
    .Q(\tms1x00.K_latch[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4671_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net3),
    .Q(\tms1x00.K_latch[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4672_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net4),
    .Q(\tms1x00.K_latch[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4673_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0503_),
    .Q(net41));
 sky130_fd_sc_hd__dfxtp_1 _4674_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0504_),
    .Q(net42));
 sky130_fd_sc_hd__dfxtp_1 _4675_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0505_),
    .Q(net43));
 sky130_fd_sc_hd__dfxtp_1 _4676_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0506_),
    .Q(net44));
 sky130_fd_sc_hd__dfxtp_1 _4677_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0507_),
    .Q(net45));
 sky130_fd_sc_hd__dfxtp_1 _4678_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0508_),
    .Q(net46));
 sky130_fd_sc_hd__dfxtp_1 _4679_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0509_),
    .Q(net47));
 sky130_fd_sc_hd__dfxtp_1 _4680_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0510_),
    .Q(net48));
 sky130_fd_sc_hd__dfxtp_1 _4681_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0511_),
    .Q(net49));
 sky130_fd_sc_hd__dfxtp_1 _4682_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0512_),
    .Q(net50));
 sky130_fd_sc_hd__dfxtp_1 _4683_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0513_),
    .Q(net51));
 sky130_fd_sc_hd__dfxtp_1 _4684_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0514_),
    .Q(net52));
 sky130_fd_sc_hd__dfxtp_1 _4685_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0515_),
    .Q(net53));
 sky130_fd_sc_hd__dfxtp_1 _4686_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0516_),
    .Q(net54));
 sky130_fd_sc_hd__dfxtp_1 _4687_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0517_),
    .Q(net55));
 sky130_fd_sc_hd__dfxtp_1 _4688_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0518_),
    .Q(net32));
 sky130_fd_sc_hd__dfxtp_1 _4689_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0519_),
    .Q(net33));
 sky130_fd_sc_hd__dfxtp_1 _4690_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0520_),
    .Q(net34));
 sky130_fd_sc_hd__dfxtp_1 _4691_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0521_),
    .Q(net35));
 sky130_fd_sc_hd__dfxtp_1 _4692_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0522_),
    .Q(net36));
 sky130_fd_sc_hd__dfxtp_1 _4693_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0523_),
    .Q(\tms1x00.CL ));
 sky130_fd_sc_hd__dfxtp_1 _4694_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0524_),
    .Q(\tms1x00.status ));
 sky130_fd_sc_hd__dfxtp_1 _4695_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0525_),
    .Q(\tms1x00.PB[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4696_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0526_),
    .Q(\tms1x00.PB[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4697_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0527_),
    .Q(\tms1x00.PB[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4698_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0528_),
    .Q(\tms1x00.PB[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4699_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0529_),
    .Q(\tms1x00.SR[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4700_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0530_),
    .Q(\tms1x00.SR[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4701_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_0531_),
    .Q(\tms1x00.SR[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4702_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_0532_),
    .Q(\tms1x00.SR[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4703_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_0533_),
    .Q(\tms1x00.SR[4] ));
 sky130_fd_sc_hd__dfxtp_1 _4704_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_0534_),
    .Q(\tms1x00.SR[5] ));
 sky130_fd_sc_hd__dfxtp_1 _4705_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_0535_),
    .Q(\tms1x00.PA[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4706_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0536_),
    .Q(\tms1x00.PA[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4707_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0537_),
    .Q(\tms1x00.PA[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4708_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0538_),
    .Q(\tms1x00.PA[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4709_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0539_),
    .Q(\tms1x00.PC[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4710_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0540_),
    .Q(\tms1x00.PC[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4711_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_0541_),
    .Q(\tms1x00.PC[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4712_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_0542_),
    .Q(\tms1x00.PC[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4713_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_0543_),
    .Q(\tms1x00.PC[4] ));
 sky130_fd_sc_hd__dfxtp_1 _4714_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_0544_),
    .Q(\tms1x00.PC[5] ));
 sky130_fd_sc_hd__dfxtp_1 _4715_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0545_),
    .Q(\tms1x00.P[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4716_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0546_),
    .Q(\tms1x00.P[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4717_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0547_),
    .Q(\tms1x00.P[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4718_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0548_),
    .Q(\tms1x00.P[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4719_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0549_),
    .Q(\tms1x00.Y[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4720_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0550_),
    .Q(\tms1x00.Y[1] ));
 sky130_fd_sc_hd__dfxtp_2 _4721_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0551_),
    .Q(\tms1x00.Y[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4722_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0552_),
    .Q(\tms1x00.Y[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4723_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0553_),
    .Q(\tms1x00.X[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4724_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0554_),
    .Q(\tms1x00.X[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4725_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0555_),
    .Q(\tms1x00.X[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4726_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0556_),
    .Q(\tms1x00.N[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4727_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0557_),
    .Q(\tms1x00.N[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4728_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0558_),
    .Q(\tms1x00.N[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4729_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0559_),
    .Q(\tms1x00.N[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4730_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0560_),
    .Q(\tms1x00.A[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4731_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0561_),
    .Q(\tms1x00.A[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4732_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0562_),
    .Q(\tms1x00.A[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4733_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0563_),
    .Q(\tms1x00.A[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4734_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0564_),
    .Q(\tms1x00.RAM[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4735_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0565_),
    .Q(\tms1x00.RAM[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4736_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0566_),
    .Q(\tms1x00.RAM[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4737_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0567_),
    .Q(\tms1x00.RAM[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4738_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0568_),
    .Q(\tms1x00.RAM[18][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4739_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0569_),
    .Q(\tms1x00.RAM[18][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4740_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0570_),
    .Q(\tms1x00.RAM[18][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4741_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0571_),
    .Q(\tms1x00.RAM[18][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4742_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0572_),
    .Q(\tms1x00.RAM[39][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4743_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0573_),
    .Q(\tms1x00.RAM[39][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4744_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0574_),
    .Q(\tms1x00.RAM[39][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4745_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0575_),
    .Q(\tms1x00.RAM[39][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4746_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0576_),
    .Q(\tms1x00.RAM[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4747_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0577_),
    .Q(\tms1x00.RAM[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4748_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0578_),
    .Q(\tms1x00.RAM[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4749_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0579_),
    .Q(\tms1x00.RAM[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4750_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0580_),
    .Q(\tms1x00.RAM[17][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4751_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0581_),
    .Q(\tms1x00.RAM[17][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4752_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0582_),
    .Q(\tms1x00.RAM[17][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4753_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0583_),
    .Q(\tms1x00.RAM[17][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4754_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0584_),
    .Q(\tms1x00.RAM[29][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4755_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0585_),
    .Q(\tms1x00.RAM[29][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4756_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0586_),
    .Q(\tms1x00.RAM[29][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4757_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0587_),
    .Q(\tms1x00.RAM[29][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4758_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0588_),
    .Q(\tms1x00.RAM[16][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4759_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0589_),
    .Q(\tms1x00.RAM[16][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4760_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0590_),
    .Q(\tms1x00.RAM[16][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4761_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0591_),
    .Q(\tms1x00.RAM[16][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4762_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0592_),
    .Q(\tms1x00.RAM[119][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4763_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0593_),
    .Q(\tms1x00.RAM[119][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4764_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0594_),
    .Q(\tms1x00.RAM[119][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4765_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0595_),
    .Q(\tms1x00.RAM[119][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4766_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0596_),
    .Q(\tms1x00.RAM[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4767_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0597_),
    .Q(\tms1x00.RAM[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4768_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0598_),
    .Q(\tms1x00.RAM[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4769_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0599_),
    .Q(\tms1x00.RAM[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4770_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0600_),
    .Q(\tms1x00.RAM[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4771_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0601_),
    .Q(\tms1x00.RAM[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4772_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0602_),
    .Q(\tms1x00.RAM[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4773_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0603_),
    .Q(\tms1x00.RAM[15][3] ));
 sky130_fd_sc_hd__dfxtp_4 _4774_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0604_),
    .Q(\tms1x00.rom_addr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4775_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0605_),
    .Q(\tms1x00.rom_addr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4776_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(_0606_),
    .Q(net57));
 sky130_fd_sc_hd__dfxtp_1 _4777_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(_0607_),
    .Q(net58));
 sky130_fd_sc_hd__dfxtp_1 _4778_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(_0608_),
    .Q(net59));
 sky130_fd_sc_hd__dfxtp_1 _4779_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(_0609_),
    .Q(net60));
 sky130_fd_sc_hd__dfxtp_1 _4780_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_0610_),
    .Q(net61));
 sky130_fd_sc_hd__dfxtp_1 _4781_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_0611_),
    .Q(net62));
 sky130_fd_sc_hd__dfxtp_1 _4782_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0612_),
    .Q(net63));
 sky130_fd_sc_hd__dfxtp_1 _4783_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0613_),
    .Q(net64));
 sky130_fd_sc_hd__dfxtp_1 _4784_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0614_),
    .Q(\tms1x00.RAM[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4785_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0615_),
    .Q(\tms1x00.RAM[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4786_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0616_),
    .Q(\tms1x00.RAM[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4787_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0617_),
    .Q(\tms1x00.RAM[9][3] ));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_126 (.HI(net126));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_127 (.HI(net127));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_128 (.HI(net128));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_129 (.HI(net129));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_130 (.HI(net130));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_131 (.HI(net131));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_132 (.HI(net132));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_133 (.HI(net133));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_79 (.LO(net79));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_80 (.LO(net80));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_81 (.LO(net81));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_82 (.LO(net82));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_83 (.LO(net83));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_84 (.LO(net84));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_85 (.LO(net85));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_86 (.LO(net86));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_87 (.LO(net87));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_88 (.LO(net88));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_89 (.LO(net89));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_90 (.LO(net90));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_91 (.LO(net91));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_92 (.LO(net92));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_93 (.LO(net93));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_94 (.LO(net94));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_95 (.LO(net95));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_96 (.LO(net96));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_97 (.LO(net97));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_98 (.LO(net98));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_99 (.LO(net99));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_100 (.LO(net100));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_101 (.LO(net101));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_102 (.LO(net102));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_103 (.LO(net103));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_104 (.LO(net104));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_105 (.LO(net105));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_106 (.LO(net106));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_107 (.LO(net107));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_108 (.LO(net108));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_109 (.LO(net109));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_110 (.LO(net110));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_111 (.LO(net111));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_112 (.LO(net112));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_113 (.LO(net113));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_114 (.LO(net114));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_115 (.LO(net115));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_116 (.LO(net116));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_117 (.LO(net117));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_118 (.LO(net118));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_119 (.LO(net119));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_120 (.LO(net120));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_121 (.LO(net121));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_122 (.LO(net122));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_123 (.LO(net123));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_124 (.LO(net124));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_125 (.HI(net125));
 sky130_fd_sc_hd__clkbuf_1 _4844_ (.A(net16),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_2 _4845_ (.A(net17),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_2 _4846_ (.A(net19),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 _4847_ (.A(net21),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_2 _4848_ (.A(net22),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_2 _4849_ (.A(net23),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_2 _4850_ (.A(net24),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_2 _4851_ (.A(net25),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_2 _4852_ (.A(net26),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_1 _4853_ (.A(net27),
    .X(net74));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(io_in[6]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(io_in[7]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(io_in[8]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(io_in[9]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(oram_value[0]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(oram_value[10]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(oram_value[1]),
    .X(net7));
 sky130_fd_sc_hd__dlymetal6s2s_1 input8 (.A(oram_value[2]),
    .X(net8));
 sky130_fd_sc_hd__dlymetal6s2s_1 input9 (.A(oram_value[3]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(oram_value[4]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(oram_value[5]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(oram_value[6]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(oram_value[7]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(oram_value[8]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(oram_value[9]),
    .X(net15));
 sky130_fd_sc_hd__buf_2 input16 (.A(wb_rst_i),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(wbs_adr_i[0]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(wbs_adr_i[16]),
    .X(net18));
 sky130_fd_sc_hd__dlymetal6s2s_1 input19 (.A(wbs_adr_i[1]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(wbs_adr_i[23]),
    .X(net20));
 sky130_fd_sc_hd__dlymetal6s2s_1 input21 (.A(wbs_adr_i[2]),
    .X(net21));
 sky130_fd_sc_hd__dlymetal6s2s_1 input22 (.A(wbs_adr_i[3]),
    .X(net22));
 sky130_fd_sc_hd__dlymetal6s2s_1 input23 (.A(wbs_adr_i[4]),
    .X(net23));
 sky130_fd_sc_hd__dlymetal6s2s_1 input24 (.A(wbs_adr_i[5]),
    .X(net24));
 sky130_fd_sc_hd__dlymetal6s2s_1 input25 (.A(wbs_adr_i[6]),
    .X(net25));
 sky130_fd_sc_hd__dlymetal6s2s_1 input26 (.A(wbs_adr_i[7]),
    .X(net26));
 sky130_fd_sc_hd__dlymetal6s2s_1 input27 (.A(wbs_adr_i[8]),
    .X(net27));
 sky130_fd_sc_hd__dlymetal6s2s_1 input28 (.A(wbs_cyc_i),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(wbs_dat_i),
    .X(net29));
 sky130_fd_sc_hd__dlymetal6s2s_1 input30 (.A(wbs_stb_i),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_2 input31 (.A(wbs_we_i),
    .X(net31));
 sky130_fd_sc_hd__buf_2 output32 (.A(net32),
    .X(io_out[10]));
 sky130_fd_sc_hd__buf_2 output33 (.A(net33),
    .X(io_out[11]));
 sky130_fd_sc_hd__buf_2 output34 (.A(net34),
    .X(io_out[12]));
 sky130_fd_sc_hd__buf_2 output35 (.A(net35),
    .X(io_out[13]));
 sky130_fd_sc_hd__buf_2 output36 (.A(net36),
    .X(io_out[14]));
 sky130_fd_sc_hd__buf_2 output37 (.A(net37),
    .X(io_out[15]));
 sky130_fd_sc_hd__buf_2 output38 (.A(net38),
    .X(io_out[16]));
 sky130_fd_sc_hd__buf_2 output39 (.A(net39),
    .X(io_out[17]));
 sky130_fd_sc_hd__buf_2 output40 (.A(net40),
    .X(io_out[18]));
 sky130_fd_sc_hd__buf_2 output41 (.A(net41),
    .X(io_out[19]));
 sky130_fd_sc_hd__buf_2 output42 (.A(net42),
    .X(io_out[20]));
 sky130_fd_sc_hd__buf_2 output43 (.A(net43),
    .X(io_out[21]));
 sky130_fd_sc_hd__buf_2 output44 (.A(net44),
    .X(io_out[22]));
 sky130_fd_sc_hd__buf_2 output45 (.A(net45),
    .X(io_out[23]));
 sky130_fd_sc_hd__buf_2 output46 (.A(net46),
    .X(io_out[24]));
 sky130_fd_sc_hd__buf_2 output47 (.A(net47),
    .X(io_out[25]));
 sky130_fd_sc_hd__buf_2 output48 (.A(net48),
    .X(io_out[26]));
 sky130_fd_sc_hd__buf_2 output49 (.A(net49),
    .X(io_out[27]));
 sky130_fd_sc_hd__buf_2 output50 (.A(net50),
    .X(io_out[28]));
 sky130_fd_sc_hd__buf_2 output51 (.A(net51),
    .X(io_out[29]));
 sky130_fd_sc_hd__buf_2 output52 (.A(net52),
    .X(io_out[30]));
 sky130_fd_sc_hd__buf_2 output53 (.A(net53),
    .X(io_out[31]));
 sky130_fd_sc_hd__buf_2 output54 (.A(net54),
    .X(io_out[32]));
 sky130_fd_sc_hd__buf_2 output55 (.A(net55),
    .X(io_out[33]));
 sky130_fd_sc_hd__buf_2 output56 (.A(net56),
    .X(io_out[37]));
 sky130_fd_sc_hd__buf_2 output57 (.A(net57),
    .X(oram_addr[0]));
 sky130_fd_sc_hd__buf_2 output58 (.A(net58),
    .X(oram_addr[1]));
 sky130_fd_sc_hd__buf_2 output59 (.A(net59),
    .X(oram_addr[2]));
 sky130_fd_sc_hd__buf_2 output60 (.A(net60),
    .X(oram_addr[3]));
 sky130_fd_sc_hd__buf_2 output61 (.A(net61),
    .X(oram_addr[4]));
 sky130_fd_sc_hd__buf_2 output62 (.A(net62),
    .X(oram_addr[5]));
 sky130_fd_sc_hd__buf_2 output63 (.A(net63),
    .X(oram_addr[6]));
 sky130_fd_sc_hd__buf_2 output64 (.A(net64),
    .X(oram_addr[7]));
 sky130_fd_sc_hd__buf_2 output65 (.A(net65),
    .X(oram_csb));
 sky130_fd_sc_hd__buf_2 output66 (.A(net66),
    .X(ram_adrb[0]));
 sky130_fd_sc_hd__buf_2 output67 (.A(net67),
    .X(ram_adrb[1]));
 sky130_fd_sc_hd__buf_2 output68 (.A(net68),
    .X(ram_adrb[2]));
 sky130_fd_sc_hd__buf_2 output69 (.A(net69),
    .X(ram_adrb[3]));
 sky130_fd_sc_hd__buf_2 output70 (.A(net70),
    .X(ram_adrb[4]));
 sky130_fd_sc_hd__buf_2 output71 (.A(net71),
    .X(ram_adrb[5]));
 sky130_fd_sc_hd__buf_2 output72 (.A(net72),
    .X(ram_adrb[6]));
 sky130_fd_sc_hd__buf_2 output73 (.A(net73),
    .X(ram_adrb[7]));
 sky130_fd_sc_hd__buf_2 output74 (.A(net74),
    .X(ram_adrb[8]));
 sky130_fd_sc_hd__buf_2 output75 (.A(net75),
    .X(ram_csb));
 sky130_fd_sc_hd__buf_2 output76 (.A(net76),
    .X(ram_web));
 sky130_fd_sc_hd__buf_2 output77 (.A(net77),
    .X(wbs_ack_o));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_78 (.LO(net78));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_21_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_23_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_25_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_26_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_28_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_29_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_32_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_33_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_34_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_36_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_37_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_38_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_39_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_40_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_41_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_42_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__2529__S1 (.DIODE(_0002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2226__A (.DIODE(_0002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2218__A (.DIODE(_0002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2189__A (.DIODE(_0002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2184__A (.DIODE(_0002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2169__A (.DIODE(_0002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2146__A (.DIODE(_0002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2547__B1 (.DIODE(_0004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2507__B1 (.DIODE(_0004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2228__A (.DIODE(_0004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2197__A (.DIODE(_0004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2178__A (.DIODE(_0004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2164__A (.DIODE(_0004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2610__C1 (.DIODE(_0005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2553__A1 (.DIODE(_0005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2541__B1 (.DIODE(_0005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2330__C1 (.DIODE(_0005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2243__A (.DIODE(_0005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2183__A (.DIODE(_0005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2181__A (.DIODE(_0005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2613__A1 (.DIODE(_0007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2612__A (.DIODE(_0007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2467__C1 (.DIODE(_0007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2365__B1 (.DIODE(_0007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2298__A (.DIODE(_0007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2246__C1 (.DIODE(_0007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4003__A1 (.DIODE(_0619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3983__A1 (.DIODE(_0619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3839__B (.DIODE(_0619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3830__B (.DIODE(_0619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3829__B (.DIODE(_0619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3825__C_N (.DIODE(_0619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3767__A0 (.DIODE(_0619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2133__C (.DIODE(_0619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2122__C (.DIODE(_0619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2098__A0 (.DIODE(_0619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3924__C (.DIODE(_0621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3866__A (.DIODE(_0621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3832__A (.DIODE(_0621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3807__A (.DIODE(_0621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2139__A (.DIODE(_0621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2096__A (.DIODE(_0621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3956__A1 (.DIODE(_0623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3955__A1 (.DIODE(_0623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3824__A2 (.DIODE(_0623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3821__A2 (.DIODE(_0623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3816__S (.DIODE(_0623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3808__A2 (.DIODE(_0623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3803__B (.DIODE(_0623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3794__S (.DIODE(_0623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3790__S (.DIODE(_0623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2096__B (.DIODE(_0623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4010__A1 (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3987__A1 (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3839__A (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3829__C_N (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3826__B (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3825__B (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3769__A0 (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2133__B (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2122__B (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2102__A0 (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4017__A1 (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3839__C_N (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3830__A (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3829__A (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3826__A (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3825__A (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3771__A0 (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2133__A (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2122__A (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2105__A0 (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3995__A1 (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3877__A1 (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3874__A1 (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3871__A1 (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3868__A1 (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3864__A1 (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3862__A1 (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3860__A1 (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3858__A1 (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2108__A (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4022__A1 (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3876__A (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3873__A (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3870__A (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3842__A1 (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3833__A1 (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3828__A1 (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3773__A0 (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2140__A1 (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2109__A0 (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4052__A (.DIODE(_0635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3775__A1 (.DIODE(_0635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3357__A (.DIODE(_0635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3184__C_N (.DIODE(_0635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2935__A (.DIODE(_0635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2725__C (.DIODE(_0635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2692__A (.DIODE(_0635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2666__A (.DIODE(_0635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2653__A_N (.DIODE(_0635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2112__A1 (.DIODE(_0635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4052__B (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3777__A1 (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3357__C_N (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3184__A (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2935__B (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2725__A_N (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2692__B (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2666__B (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2653__B (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2115__A1 (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4052__C (.DIODE(_0639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3779__A1 (.DIODE(_0639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3515__A (.DIODE(_0639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3357__B (.DIODE(_0639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3184__B (.DIODE(_0639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2725__B (.DIODE(_0639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2692__C (.DIODE(_0639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2666__C_N (.DIODE(_0639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2653__C (.DIODE(_0639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2118__A1 (.DIODE(_0639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4029__A (.DIODE(_0642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3971__A1 (.DIODE(_0642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3921__A0 (.DIODE(_0642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3895__A2 (.DIODE(_0642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3892__A1 (.DIODE(_0642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3889__A1 (.DIODE(_0642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3886__A1 (.DIODE(_0642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3883__A1 (.DIODE(_0642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3824__A1 (.DIODE(_0642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2129__A (.DIODE(_0642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4026__A (.DIODE(_0643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3979__B (.DIODE(_0643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3968__A1 (.DIODE(_0643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3917__A0 (.DIODE(_0643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3880__D (.DIODE(_0643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3821__A1 (.DIODE(_0643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2615__B (.DIODE(_0643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2516__A (.DIODE(_0643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2300__A2 (.DIODE(_0643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2129__B (.DIODE(_0643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3869__A2 (.DIODE(_0648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3865__B (.DIODE(_0648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3855__B (.DIODE(_0648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3850__B (.DIODE(_0648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3845__B (.DIODE(_0648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3836__B (.DIODE(_0648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2130__A (.DIODE(_0648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3878__A1 (.DIODE(_0649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3875__A1 (.DIODE(_0649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3872__A1 (.DIODE(_0649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3863__A2 (.DIODE(_0649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3861__A2 (.DIODE(_0649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3859__A3 (.DIODE(_0649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3842__A2 (.DIODE(_0649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3833__A2 (.DIODE(_0649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3828__A2 (.DIODE(_0649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2140__A3 (.DIODE(_0649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3864__A2 (.DIODE(_0655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3858__A3 (.DIODE(_0655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3854__A2 (.DIODE(_0655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3849__A2 (.DIODE(_0655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3844__A2 (.DIODE(_0655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3835__A2 (.DIODE(_0655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2137__A (.DIODE(_0655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4033__C1 (.DIODE(_0658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4031__C1 (.DIODE(_0658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4028__C1 (.DIODE(_0658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4022__C1 (.DIODE(_0658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4017__C1 (.DIODE(_0658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4010__C1 (.DIODE(_0658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4003__C1 (.DIODE(_0658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3896__C1 (.DIODE(_0658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3828__C1 (.DIODE(_0658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2140__C1 (.DIODE(_0658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2546__S1 (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2538__S1 (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2506__S1 (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2459__S1 (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2404__S1 (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2357__S1 (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2235__S1 (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2176__A (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2162__A (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2147__A (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2543__A (.DIODE(_0665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2537__S1 (.DIODE(_0665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2528__S1 (.DIODE(_0665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2525__A1 (.DIODE(_0665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2523__A_N (.DIODE(_0665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2324__S1 (.DIODE(_0665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2273__S1 (.DIODE(_0665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2247__A (.DIODE(_0665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2152__A (.DIODE(_0665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2148__A (.DIODE(_0665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2587__A1 (.DIODE(_0666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2545__A (.DIODE(_0666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2494__A (.DIODE(_0666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2447__A (.DIODE(_0666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2425__A1 (.DIODE(_0666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2392__A (.DIODE(_0666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2345__A (.DIODE(_0666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2323__A1 (.DIODE(_0666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2215__A (.DIODE(_0666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2158__A1 (.DIODE(_0666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2546__S0 (.DIODE(_0667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2542__S (.DIODE(_0667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2524__S (.DIODE(_0667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2506__S0 (.DIODE(_0667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2459__S0 (.DIODE(_0667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2421__S (.DIODE(_0667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2404__S0 (.DIODE(_0667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2357__S0 (.DIODE(_0667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2175__A (.DIODE(_0667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2150__S (.DIODE(_0667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2581__A1 (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2477__A1 (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2442__A1 (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2424__A (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2375__A1 (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2340__A1 (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2322__A (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2259__A1 (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2204__A1 (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2156__A (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2538__S0 (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2529__S0 (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2522__S (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2319__S (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2264__A (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2201__A (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2191__A (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2186__A (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2161__A (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2154__A (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2594__S (.DIODE(_0672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2584__S (.DIODE(_0672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2580__S (.DIODE(_0672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2562__S (.DIODE(_0672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2537__S0 (.DIODE(_0672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2476__S (.DIODE(_0672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2439__S (.DIODE(_0672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2423__S (.DIODE(_0672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2199__S (.DIODE(_0672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2155__S (.DIODE(_0672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2547__A1 (.DIODE(_0677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2507__A1 (.DIODE(_0677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2460__A1 (.DIODE(_0677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2405__A1 (.DIODE(_0677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2358__A1 (.DIODE(_0677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2291__A1 (.DIODE(_0677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2236__A1 (.DIODE(_0677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2196__A (.DIODE(_0677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2166__A (.DIODE(_0677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2160__A (.DIODE(_0677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2548__A1 (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2499__A1 (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2452__A1 (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2427__A1 (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2397__A1 (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2350__A1 (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2325__A1 (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2283__A1 (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2221__A1 (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2165__A1 (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2558__S0 (.DIODE(_0679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2483__S (.DIODE(_0679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2426__S0 (.DIODE(_0679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2391__S (.DIODE(_0679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2381__S (.DIODE(_0679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2344__S (.DIODE(_0679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2324__S0 (.DIODE(_0679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2277__S (.DIODE(_0679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2267__S (.DIODE(_0679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2163__S0 (.DIODE(_0679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2558__S1 (.DIODE(_0680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2496__A (.DIODE(_0680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2472__S1 (.DIODE(_0680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2449__A (.DIODE(_0680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2426__S1 (.DIODE(_0680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2370__S1 (.DIODE(_0680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2347__A (.DIODE(_0680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2328__S1 (.DIODE(_0680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2217__A (.DIODE(_0680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2163__S1 (.DIODE(_0680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2165__A2 (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2510__S0 (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2463__S0 (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2450__S0 (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2408__S0 (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2361__S0 (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2294__S0 (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2290__S0 (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2241__S0 (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2235__S0 (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2168__A (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2582__S0 (.DIODE(_0686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2564__S0 (.DIODE(_0686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2549__S0 (.DIODE(_0686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2478__S0 (.DIODE(_0686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2428__S0 (.DIODE(_0686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2376__S0 (.DIODE(_0686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2341__S0 (.DIODE(_0686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2326__S0 (.DIODE(_0686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2260__S0 (.DIODE(_0686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2171__S0 (.DIODE(_0686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2606__S1 (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2602__S1 (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2599__S1 (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2550__S1 (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2504__S1 (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2497__S1 (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2395__S1 (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2355__S1 (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2348__S1 (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2170__A (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2598__S1 (.DIODE(_0688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2588__S1 (.DIODE(_0688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2555__A_N (.DIODE(_0688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2500__S1 (.DIODE(_0688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2453__S1 (.DIODE(_0688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2443__S1 (.DIODE(_0688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2260__S1 (.DIODE(_0688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2223__S1 (.DIODE(_0688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2207__S1 (.DIODE(_0688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2171__S1 (.DIODE(_0688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2609__A1 (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2540__A1 (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2534__A (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2490__A1 (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2471__C1 (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2431__A1 (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2388__A1 (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2329__A1 (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2274__A1 (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2180__A1 (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2596__S0 (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2472__S0 (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2437__S0 (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2430__S0 (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2370__S0 (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2335__S0 (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2328__S0 (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2253__S0 (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2195__S0 (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2177__S0 (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2596__S1 (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2549__S1 (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2437__S1 (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2430__S1 (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2394__A (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2335__S1 (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2280__A (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2253__S1 (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2195__S1 (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2177__S1 (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2597__C1 (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2527__C1 (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2490__B1 (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2431__B1 (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2396__B1 (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2388__B1 (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2329__B1 (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2282__B1 (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2274__B1 (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2180__B1 (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2513__A1 (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2492__A1 (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2466__A1 (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2432__C1 (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2411__A1 (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2390__A1 (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2364__A1 (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2297__A1 (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2245__A1 (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2182__C1 (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2604__S1 (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2508__S1 (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2457__S1 (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2406__S1 (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2402__S1 (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2359__S1 (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2288__S1 (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2281__S1 (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2233__S1 (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2185__A (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2593__A_N (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2470__A_N (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2434__A_N (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2398__S1 (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2368__A_N (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2351__S1 (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2332__A_N (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2284__S1 (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2251__A_N (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2188__A_N (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2592__S (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2578__S (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2560__S (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2556__S (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2489__S0 (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2474__S (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2372__S (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2285__S0 (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2250__S (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2187__S (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2535__S1 (.DIODE(_0707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2533__S1 (.DIODE(_0707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2526__S1 (.DIODE(_0707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2501__S1 (.DIODE(_0707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2489__S1 (.DIODE(_0707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2399__S1 (.DIODE(_0707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2387__S1 (.DIODE(_0707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2352__S1 (.DIODE(_0707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2285__S1 (.DIODE(_0707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2190__A (.DIODE(_0707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2595__A1 (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2585__A_N (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2575__S1 (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2563__A1 (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2440__A_N (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2436__A1 (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2334__A1 (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2272__S1 (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2200__A_N (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2194__A1 (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2570__S (.DIODE(_0709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2528__S0 (.DIODE(_0709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2435__S (.DIODE(_0709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2387__S0 (.DIODE(_0709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2337__S (.DIODE(_0709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2333__S (.DIODE(_0709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2321__S (.DIODE(_0709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2273__S0 (.DIODE(_0709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2256__S (.DIODE(_0709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2192__S (.DIODE(_0709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2595__B1 (.DIODE(_0711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2563__B1 (.DIODE(_0711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2557__B1 (.DIODE(_0711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2511__A1 (.DIODE(_0711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2436__B1 (.DIODE(_0711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2409__A1 (.DIODE(_0711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2362__A1 (.DIODE(_0711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2334__B1 (.DIODE(_0711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2222__A (.DIODE(_0711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2194__B1 (.DIODE(_0711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2198__B1 (.DIODE(_0713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2586__S (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2544__S (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2493__S (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2446__S (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2441__S (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2374__S (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2339__S (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2258__S (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2214__S (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2202__S (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2587__B1 (.DIODE(_0721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2551__A1 (.DIODE(_0721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2505__A (.DIODE(_0721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2458__A (.DIODE(_0721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2442__B1 (.DIODE(_0721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2403__A (.DIODE(_0721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2356__A (.DIODE(_0721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2289__A (.DIODE(_0721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2234__A (.DIODE(_0721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2204__B1 (.DIODE(_0721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2602__S0 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2599__S0 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2550__S0 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2497__S0 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2448__S (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2395__S0 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2348__S0 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2219__S0 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2216__S (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2206__A (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2598__S0 (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2588__S0 (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2500__S0 (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2453__S0 (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2443__S0 (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2398__S0 (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2351__S0 (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2284__S0 (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2223__S0 (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2207__S0 (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2212__B1 (.DIODE(_0725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2607__A (.DIODE(_0726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2509__A (.DIODE(_0726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2498__A1 (.DIODE(_0726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2451__A1 (.DIODE(_0726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2396__A1 (.DIODE(_0726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2360__A (.DIODE(_0726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2349__A1 (.DIODE(_0726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2282__A1 (.DIODE(_0726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2220__A1 (.DIODE(_0726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2209__A (.DIODE(_0726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2601__A1 (.DIODE(_0727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2589__B2 (.DIODE(_0727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2577__A1 (.DIODE(_0727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2573__A1 (.DIODE(_0727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2491__A1 (.DIODE(_0727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2444__B2 (.DIODE(_0727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2389__A1 (.DIODE(_0727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2275__A1 (.DIODE(_0727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2261__B2 (.DIODE(_0727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2212__B2 (.DIODE(_0727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2609__B1 (.DIODE(_0728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2551__B1 (.DIODE(_0728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2498__B1 (.DIODE(_0728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2464__B1 (.DIODE(_0728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2451__B1 (.DIODE(_0728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2349__B1 (.DIODE(_0728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2295__B1 (.DIODE(_0728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2242__B1 (.DIODE(_0728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2220__B1 (.DIODE(_0728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2211__A (.DIODE(_0728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2589__C1 (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2576__B1 (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2565__C1 (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2541__A1 (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2480__A1 (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2444__C1 (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2378__A1 (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2342__C1 (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2262__A1 (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2212__C1 (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2510__S1 (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2463__S1 (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2450__S1 (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2408__S1 (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2361__S1 (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2294__S1 (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2290__S1 (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2263__A (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2241__S1 (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2219__S1 (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2576__A1 (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2572__C1 (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2503__A1 (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2456__A1 (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2401__A1 (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2369__C1 (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2354__A1 (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2287__A1 (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2252__C1 (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2230__A1 (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2605__A1 (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2486__A1 (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2462__A (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2455__A1 (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2407__A (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2384__A1 (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2293__A (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2270__A1 (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2239__A (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2229__A1 (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2554__S (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2501__S0 (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2485__S0 (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2481__S (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2454__S0 (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2383__S0 (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2379__S (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2269__S0 (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2248__A (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2227__S0 (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2608__S1 (.DIODE(_0744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2485__S1 (.DIODE(_0744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2461__S1 (.DIODE(_0744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2454__S1 (.DIODE(_0744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2383__S1 (.DIODE(_0744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2292__S1 (.DIODE(_0744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2269__S1 (.DIODE(_0744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2255__A (.DIODE(_0744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2238__S1 (.DIODE(_0744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2227__S1 (.DIODE(_0744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2605__B1 (.DIODE(_0746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2502__B1 (.DIODE(_0746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2460__B1 (.DIODE(_0746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2455__B1 (.DIODE(_0746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2405__B1 (.DIODE(_0746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2358__B1 (.DIODE(_0746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2353__B1 (.DIODE(_0746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2291__B1 (.DIODE(_0746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2236__B1 (.DIODE(_0746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2229__B1 (.DIODE(_0746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2513__C1 (.DIODE(_0749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2466__B1 (.DIODE(_0749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2411__C1 (.DIODE(_0749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2364__C1 (.DIODE(_0749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2297__C1 (.DIODE(_0749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2245__B1 (.DIODE(_0749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2606__S0 (.DIODE(_0750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2504__S0 (.DIODE(_0750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2495__S (.DIODE(_0750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2457__S0 (.DIODE(_0750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2402__S0 (.DIODE(_0750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2393__S (.DIODE(_0750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2355__S0 (.DIODE(_0750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2346__S (.DIODE(_0750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2281__S0 (.DIODE(_0750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2233__S0 (.DIODE(_0750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2234__B (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2236__A2 (.DIODE(_0753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2244__A2 (.DIODE(_0754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2608__S0 (.DIODE(_0755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2604__S0 (.DIODE(_0755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2508__S0 (.DIODE(_0755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2461__S0 (.DIODE(_0755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2406__S0 (.DIODE(_0755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2359__S0 (.DIODE(_0755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2292__S0 (.DIODE(_0755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2288__S0 (.DIODE(_0755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2279__S (.DIODE(_0755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2238__S0 (.DIODE(_0755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2603__A (.DIODE(_0758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2600__A (.DIODE(_0758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2581__B1 (.DIODE(_0758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2477__B1 (.DIODE(_0758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2464__A1 (.DIODE(_0758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2375__B1 (.DIODE(_0758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2340__B1 (.DIODE(_0758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2295__A1 (.DIODE(_0758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2259__B1 (.DIODE(_0758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2242__A1 (.DIODE(_0758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2242__A2 (.DIODE(_0759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2244__B2 (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2611__A1 (.DIODE(_0761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2532__A1 (.DIODE(_0761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2512__C1 (.DIODE(_0761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2465__C1 (.DIODE(_0761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2410__C1 (.DIODE(_0761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2363__C1 (.DIODE(_0761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2296__C1 (.DIODE(_0761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2244__C1 (.DIODE(_0761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3976__A (.DIODE(_0764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2300__B1 (.DIODE(_0764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2574__S1 (.DIODE(_0765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2572__A1 (.DIODE(_0765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2568__S1 (.DIODE(_0765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2484__A (.DIODE(_0765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2471__A1 (.DIODE(_0765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2382__A (.DIODE(_0765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2369__A1 (.DIODE(_0765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2278__A (.DIODE(_0765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2268__A (.DIODE(_0765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2252__A1 (.DIODE(_0765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2575__S0 (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2574__S0 (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2569__S (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2568__S0 (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2488__S0 (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2468__S (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2386__S0 (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2366__S (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2272__S0 (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2249__S (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2254__B (.DIODE(_0771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2579__A_N (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2571__A_N (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2561__A_N (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2557__A1 (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2488__S1 (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2475__A_N (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2386__S1 (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2373__A_N (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2338__A_N (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2257__A_N (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2259__A2 (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2582__S1 (.DIODE(_0781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2564__S1 (.DIODE(_0781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2482__A (.DIODE(_0781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2478__S1 (.DIODE(_0781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2428__S1 (.DIODE(_0781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2380__A (.DIODE(_0781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2376__S1 (.DIODE(_0781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2341__S1 (.DIODE(_0781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2326__S1 (.DIODE(_0781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2266__A (.DIODE(_0781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2535__S0 (.DIODE(_0782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2533__S0 (.DIODE(_0782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2526__S0 (.DIODE(_0782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2469__S (.DIODE(_0782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2433__S (.DIODE(_0782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2399__S0 (.DIODE(_0782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2367__S (.DIODE(_0782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2352__S0 (.DIODE(_0782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2331__S (.DIODE(_0782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2265__S (.DIODE(_0782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2268__B (.DIODE(_0785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2287__B1 (.DIODE(_0804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2291__A2 (.DIODE(_0808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3976__B (.DIODE(_0817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2300__B2 (.DIODE(_0817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2818__A (.DIODE(_0825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2308__A (.DIODE(_0825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3736__A (.DIODE(_0826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3534__A (.DIODE(_0826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3475__A (.DIODE(_0826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3326__A (.DIODE(_0826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3304__A (.DIODE(_0826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3125__A (.DIODE(_0826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3000__A (.DIODE(_0826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2893__A (.DIODE(_0826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2621__A (.DIODE(_0826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2309__A (.DIODE(_0826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2757__A0 (.DIODE(_0827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2747__A0 (.DIODE(_0827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2738__A0 (.DIODE(_0827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2727__A0 (.DIODE(_0827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2717__A0 (.DIODE(_0827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2707__A0 (.DIODE(_0827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2694__A0 (.DIODE(_0827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2670__A0 (.DIODE(_0827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2658__A0 (.DIODE(_0827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2317__A0 (.DIODE(_0827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3022__A (.DIODE(_0829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3013__A (.DIODE(_0829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2908__A (.DIODE(_0829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2884__A (.DIODE(_0829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2873__A (.DIODE(_0829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2864__A (.DIODE(_0829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2855__A (.DIODE(_0829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2846__A (.DIODE(_0829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2837__A (.DIODE(_0829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2316__A (.DIODE(_0829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3737__A (.DIODE(_0833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3565__A (.DIODE(_0833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3466__A (.DIODE(_0833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3327__A (.DIODE(_0833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3277__A (.DIODE(_0833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2937__A (.DIODE(_0833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2716__A (.DIODE(_0833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2316__B (.DIODE(_0833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2336__B1 (.DIODE(_0852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2342__B1 (.DIODE(_0858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2358__A2 (.DIODE(_0874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2362__A2 (.DIODE(_0878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2363__B2 (.DIODE(_0879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3985__A (.DIODE(_0882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2414__A1 (.DIODE(_0882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2375__A2 (.DIODE(_0891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2382__B (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2384__A2 (.DIODE(_0900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2401__B1 (.DIODE(_0917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2407__B (.DIODE(_0923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2409__A2 (.DIODE(_0925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3985__B (.DIODE(_0929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2414__A2 (.DIODE(_0929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3740__A (.DIODE(_0934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3538__A (.DIODE(_0934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3479__A (.DIODE(_0934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3330__A (.DIODE(_0934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3308__A (.DIODE(_0934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3129__A (.DIODE(_0934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3004__A (.DIODE(_0934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2898__A (.DIODE(_0934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2630__A (.DIODE(_0934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2418__A (.DIODE(_0934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2759__A0 (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2749__A0 (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2740__A0 (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2729__A0 (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2719__A0 (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2709__A0 (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2696__A0 (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2672__A0 (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2660__A0 (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2419__A0 (.DIODE(_0935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2427__A2 (.DIODE(_0942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2431__A2 (.DIODE(_0946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2438__B1 (.DIODE(_0953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2444__B1 (.DIODE(_0959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2458__B (.DIODE(_0973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2460__A2 (.DIODE(_0975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2464__A2 (.DIODE(_0979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3989__A (.DIODE(_0983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2515__A1 (.DIODE(_0983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2477__A2 (.DIODE(_0992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2484__B (.DIODE(_0999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2486__A2 (.DIODE(_1001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2509__B (.DIODE(_1024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3989__B (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2515__A2 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2829__A (.DIODE(_1033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2518__A (.DIODE(_1033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3743__A (.DIODE(_1034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3541__A (.DIODE(_1034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3482__A (.DIODE(_1034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3333__A (.DIODE(_1034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3311__A (.DIODE(_1034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3132__A (.DIODE(_1034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3007__A (.DIODE(_1034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2901__A (.DIODE(_1034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2633__A (.DIODE(_1034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2519__A (.DIODE(_1034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2761__A0 (.DIODE(_1035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2751__A0 (.DIODE(_1035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2742__A0 (.DIODE(_1035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2731__A0 (.DIODE(_1035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2721__A0 (.DIODE(_1035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2711__A0 (.DIODE(_1035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2698__A0 (.DIODE(_1035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2674__A0 (.DIODE(_1035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2662__A0 (.DIODE(_1035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2520__A0 (.DIODE(_1035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2534__B (.DIODE(_1048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2540__A2 (.DIODE(_1052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2539__B (.DIODE(_1053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2547__A2 (.DIODE(_1061_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2559__B1 (.DIODE(_1073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2565__B1 (.DIODE(_1079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2572__A2 (.DIODE(_1084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2589__B1 (.DIODE(_1103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2605__A2 (.DIODE(_1119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3994__A (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2616__B1 (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2833__A (.DIODE(_1131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2617__A (.DIODE(_1131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3746__A (.DIODE(_1132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3544__A (.DIODE(_1132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3485__A (.DIODE(_1132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3336__A (.DIODE(_1132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3314__A (.DIODE(_1132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3135__A (.DIODE(_1132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3010__A (.DIODE(_1132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2904__A (.DIODE(_1132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2636__A (.DIODE(_1132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2618__A (.DIODE(_1132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2763__A0 (.DIODE(_1133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2753__A0 (.DIODE(_1133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2744__A0 (.DIODE(_1133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2733__A0 (.DIODE(_1133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2723__A0 (.DIODE(_1133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2713__A0 (.DIODE(_1133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2700__A0 (.DIODE(_1133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2676__A0 (.DIODE(_1133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2664__A0 (.DIODE(_1133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2619__A0 (.DIODE(_1133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4135__A0 (.DIODE(_1135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4126__A0 (.DIODE(_1135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2810__A1 (.DIODE(_1135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2799__A1 (.DIODE(_1135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2790__A1 (.DIODE(_1135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2777__A1 (.DIODE(_1135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2766__A1 (.DIODE(_1135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2684__A1 (.DIODE(_1135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2645__A1 (.DIODE(_1135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2628__A1 (.DIODE(_1135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3749__A (.DIODE(_1137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3727__A (.DIODE(_1137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3718__A (.DIODE(_1137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3691__A (.DIODE(_1137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2822__A (.DIODE(_1137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2809__A (.DIODE(_1137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2798__A (.DIODE(_1137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2776__A (.DIODE(_1137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2765__A (.DIODE(_1137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2627__A (.DIODE(_1137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4164__A (.DIODE(_1140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3664__A (.DIODE(_1140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3488__A (.DIODE(_1140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3305__A (.DIODE(_1140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3212__A (.DIODE(_1140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3067__A (.DIODE(_1140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2837__B (.DIODE(_1140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2627__B (.DIODE(_1140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4137__A0 (.DIODE(_1143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4128__A0 (.DIODE(_1143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2812__A1 (.DIODE(_1143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2801__A1 (.DIODE(_1143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2792__A1 (.DIODE(_1143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2779__A1 (.DIODE(_1143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2768__A1 (.DIODE(_1143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2686__A1 (.DIODE(_1143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2647__A1 (.DIODE(_1143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2631__A1 (.DIODE(_1143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4139__A0 (.DIODE(_1145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4130__A0 (.DIODE(_1145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2814__A1 (.DIODE(_1145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2803__A1 (.DIODE(_1145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2794__A1 (.DIODE(_1145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2781__A1 (.DIODE(_1145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2770__A1 (.DIODE(_1145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2688__A1 (.DIODE(_1145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2649__A1 (.DIODE(_1145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2634__A1 (.DIODE(_1145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4141__A0 (.DIODE(_1147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4132__A0 (.DIODE(_1147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2816__A1 (.DIODE(_1147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2805__A1 (.DIODE(_1147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2796__A1 (.DIODE(_1147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2783__A1 (.DIODE(_1147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2772__A1 (.DIODE(_1147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2690__A1 (.DIODE(_1147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2651__A1 (.DIODE(_1147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2637__A1 (.DIODE(_1147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3506__A (.DIODE(_1151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3497__A (.DIODE(_1151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3488__B (.DIODE(_1151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3476__A (.DIODE(_1151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3457__A (.DIODE(_1151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3448__A (.DIODE(_1151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3439__A (.DIODE(_1151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3394__A (.DIODE(_1151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2706__A (.DIODE(_1151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2644__A (.DIODE(_1151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3646__A (.DIODE(_1153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3376__A (.DIODE(_1153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3194__A (.DIODE(_1153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3086__A (.DIODE(_1153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3049__A (.DIODE(_1153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3013__B (.DIODE(_1153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2765__B (.DIODE(_1153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2644__B (.DIODE(_1153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4098__A (.DIODE(_1162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4053__A (.DIODE(_1162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3682__A (.DIODE(_1162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3535__B (.DIODE(_1162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3358__A (.DIODE(_1162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3031__A (.DIODE(_1162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2746__B (.DIODE(_1162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2657__B (.DIODE(_1162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4134__A (.DIODE(_1170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3516__B (.DIODE(_1170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3421__A (.DIODE(_1170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3241__A (.DIODE(_1170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2973__B (.DIODE(_1170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2726__B (.DIODE(_1170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2693__A (.DIODE(_1170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2669__B (.DIODE(_1170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3673__A (.DIODE(_1177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3664__B (.DIODE(_1177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3655__A (.DIODE(_1177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3646__B (.DIODE(_1177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3628__A (.DIODE(_1177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3610__A (.DIODE(_1177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3601__A (.DIODE(_1177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3583__A (.DIODE(_1177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3574__A (.DIODE(_1177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2683__A (.DIODE(_1177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3718__B (.DIODE(_1180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3556__A (.DIODE(_1180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3448__B (.DIODE(_1180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3348__A (.DIODE(_1180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3166__A (.DIODE(_1180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3107__A (.DIODE(_1180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2873__B (.DIODE(_1180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2683__B (.DIODE(_1180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4089__A (.DIODE(_1194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3758__B (.DIODE(_1194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3583__B (.DIODE(_1194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3295__A (.DIODE(_1194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3138__A (.DIODE(_1194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2955__B (.DIODE(_1194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2917__B (.DIODE(_1194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2706__B (.DIODE(_1194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4080__A (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3709__B (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3525__B (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3430__A (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3250__B (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3126__B (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2982__B (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2737__B (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4125__A (.DIODE(_1224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3637__B (.DIODE(_1224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3547__B (.DIODE(_1224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3367__A (.DIODE(_1224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3185__B (.DIODE(_1224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3040__B (.DIODE(_1224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3001__B (.DIODE(_1224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2756__B (.DIODE(_1224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3655__B (.DIODE(_1236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3476__B (.DIODE(_1236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3385__A (.DIODE(_1236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3203__B (.DIODE(_1236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3058__B (.DIODE(_1236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3022__B (.DIODE(_1236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2991__A (.DIODE(_1236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2776__B (.DIODE(_1236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4164__B (.DIODE(_1243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3700__A (.DIODE(_1243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3619__A (.DIODE(_1243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3556__B (.DIODE(_1243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3403__A (.DIODE(_1243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3259__A (.DIODE(_1243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3086__B (.DIODE(_1243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2991__B (.DIODE(_1243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2895__A (.DIODE(_1243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2789__A (.DIODE(_1243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3673__B (.DIODE(_1245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3497__B (.DIODE(_1245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3317__A (.DIODE(_1245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3221__B (.DIODE(_1245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3076__B (.DIODE(_1245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2846__B (.DIODE(_1245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2798__B (.DIODE(_1245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2789__B (.DIODE(_1245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4116__B (.DIODE(_1257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4071__A (.DIODE(_1257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3700__B (.DIODE(_1257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3601__B (.DIODE(_1257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3506__B (.DIODE(_1257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3148__B (.DIODE(_1257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2855__B (.DIODE(_1257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2809__B (.DIODE(_1257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4165__A1 (.DIODE(_1263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4072__A1 (.DIODE(_1263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3728__A1 (.DIODE(_1263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3719__A1 (.DIODE(_1263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3701__A1 (.DIODE(_1263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3674__A1 (.DIODE(_1263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3665__A1 (.DIODE(_1263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3656__A1 (.DIODE(_1263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3085__A (.DIODE(_1263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2819__A (.DIODE(_1263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3023__A1 (.DIODE(_1264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3014__A1 (.DIODE(_1264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2992__A1 (.DIODE(_1264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2885__A1 (.DIODE(_1264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2874__A1 (.DIODE(_1264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2865__A1 (.DIODE(_1264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2856__A1 (.DIODE(_1264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2847__A1 (.DIODE(_1264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2838__A1 (.DIODE(_1264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2823__A1 (.DIODE(_1264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3619__B (.DIODE(_1266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3610__B (.DIODE(_1266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3439__B (.DIODE(_1266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3339__A (.DIODE(_1266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3157__B (.DIODE(_1266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3098__B (.DIODE(_1266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2864__B (.DIODE(_1266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2822__B (.DIODE(_1266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4167__A1 (.DIODE(_1269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4074__A1 (.DIODE(_1269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3730__A1 (.DIODE(_1269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3721__A1 (.DIODE(_1269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3703__A1 (.DIODE(_1269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3676__A1 (.DIODE(_1269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3667__A1 (.DIODE(_1269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3658__A1 (.DIODE(_1269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3089__A (.DIODE(_1269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2826__A (.DIODE(_1269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3025__A1 (.DIODE(_1270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3016__A1 (.DIODE(_1270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2994__A1 (.DIODE(_1270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2887__A1 (.DIODE(_1270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2876__A1 (.DIODE(_1270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2867__A1 (.DIODE(_1270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2858__A1 (.DIODE(_1270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2849__A1 (.DIODE(_1270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2840__A1 (.DIODE(_1270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2827__A1 (.DIODE(_1270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4169__A1 (.DIODE(_1272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4076__A1 (.DIODE(_1272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3732__A1 (.DIODE(_1272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3723__A1 (.DIODE(_1272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3705__A1 (.DIODE(_1272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3678__A1 (.DIODE(_1272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3669__A1 (.DIODE(_1272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3660__A1 (.DIODE(_1272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3092__A (.DIODE(_1272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2830__A (.DIODE(_1272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3027__A1 (.DIODE(_1273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3018__A1 (.DIODE(_1273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2996__A1 (.DIODE(_1273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2889__A1 (.DIODE(_1273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2878__A1 (.DIODE(_1273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2869__A1 (.DIODE(_1273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2860__A1 (.DIODE(_1273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2851__A1 (.DIODE(_1273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2842__A1 (.DIODE(_1273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2831__A1 (.DIODE(_1273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4171__A1 (.DIODE(_1275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4078__A1 (.DIODE(_1275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3734__A1 (.DIODE(_1275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3725__A1 (.DIODE(_1275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3707__A1 (.DIODE(_1275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3680__A1 (.DIODE(_1275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3671__A1 (.DIODE(_1275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3662__A1 (.DIODE(_1275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3095__A (.DIODE(_1275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2834__A (.DIODE(_1275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3727__B (.DIODE(_1304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3628__B (.DIODE(_1304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3457__B (.DIODE(_1304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3403__B (.DIODE(_1304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3268__A (.DIODE(_1304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3175__B (.DIODE(_1304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3116__B (.DIODE(_1304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2884__B (.DIODE(_1304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2983__A0 (.DIODE(_1310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2974__A0 (.DIODE(_1310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2965__A0 (.DIODE(_1310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2956__A0 (.DIODE(_1310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2947__A0 (.DIODE(_1310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2938__A0 (.DIODE(_1310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2927__A0 (.DIODE(_1310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2918__A0 (.DIODE(_1310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2909__A0 (.DIODE(_1310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2896__A0 (.DIODE(_1310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4107__B (.DIODE(_1311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3691__B (.DIODE(_1311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3592__B (.DIODE(_1311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3412__B (.DIODE(_1311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3232__A (.DIODE(_1311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2964__B (.DIODE(_1311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2926__B (.DIODE(_1311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2895__B (.DIODE(_1311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2985__A0 (.DIODE(_1314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2976__A0 (.DIODE(_1314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2967__A0 (.DIODE(_1314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2958__A0 (.DIODE(_1314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2949__A0 (.DIODE(_1314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2940__A0 (.DIODE(_1314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2929__A0 (.DIODE(_1314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2920__A0 (.DIODE(_1314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2911__A0 (.DIODE(_1314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2899__A0 (.DIODE(_1314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2987__A0 (.DIODE(_1316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2978__A0 (.DIODE(_1316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2969__A0 (.DIODE(_1316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2960__A0 (.DIODE(_1316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2951__A0 (.DIODE(_1316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2942__A0 (.DIODE(_1316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2931__A0 (.DIODE(_1316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2922__A0 (.DIODE(_1316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2913__A0 (.DIODE(_1316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2902__A0 (.DIODE(_1316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2989__A0 (.DIODE(_1318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2980__A0 (.DIODE(_1318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2971__A0 (.DIODE(_1318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2962__A0 (.DIODE(_1318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2953__A0 (.DIODE(_1318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2944__A0 (.DIODE(_1318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2933__A0 (.DIODE(_1318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2924__A0 (.DIODE(_1318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2915__A0 (.DIODE(_1318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2905__A0 (.DIODE(_1318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4062__B (.DIODE(_1320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3749__B (.DIODE(_1320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3574__B (.DIODE(_1320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3394__B (.DIODE(_1320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3286__A (.DIODE(_1320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3259__B (.DIODE(_1320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2946__B (.DIODE(_1320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2908__B (.DIODE(_1320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4116__A (.DIODE(_1337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3116__A (.DIODE(_1337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3098__A (.DIODE(_1337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3076__A (.DIODE(_1337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3058__A (.DIODE(_1337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3049__B (.DIODE(_1337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2964__A (.DIODE(_1337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2955__A (.DIODE(_1337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2946__A (.DIODE(_1337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2937__B (.DIODE(_1337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3117__A0 (.DIODE(_1373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3108__A0 (.DIODE(_1373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3099__A0 (.DIODE(_1373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3077__A0 (.DIODE(_1373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3068__A0 (.DIODE(_1373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3059__A0 (.DIODE(_1373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3050__A0 (.DIODE(_1373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3041__A0 (.DIODE(_1373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3032__A0 (.DIODE(_1373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3002__A0 (.DIODE(_1373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3119__A0 (.DIODE(_1376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3110__A0 (.DIODE(_1376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3101__A0 (.DIODE(_1376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3079__A0 (.DIODE(_1376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3070__A0 (.DIODE(_1376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3061__A0 (.DIODE(_1376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3052__A0 (.DIODE(_1376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3043__A0 (.DIODE(_1376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3034__A0 (.DIODE(_1376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3005__A0 (.DIODE(_1376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3121__A0 (.DIODE(_1378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3112__A0 (.DIODE(_1378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3103__A0 (.DIODE(_1378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3081__A0 (.DIODE(_1378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3072__A0 (.DIODE(_1378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3063__A0 (.DIODE(_1378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3054__A0 (.DIODE(_1378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3045__A0 (.DIODE(_1378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3036__A0 (.DIODE(_1378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3008__A0 (.DIODE(_1378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3123__A0 (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3114__A0 (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3105__A0 (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3083__A0 (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3074__A0 (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3065__A0 (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3056__A0 (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3047__A0 (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3038__A0 (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3011__A0 (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3269__A1 (.DIODE(_1422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3222__A1 (.DIODE(_1422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3213__A1 (.DIODE(_1422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3204__A1 (.DIODE(_1422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3195__A1 (.DIODE(_1422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3176__A1 (.DIODE(_1422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3167__A1 (.DIODE(_1422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3158__A1 (.DIODE(_1422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3149__A1 (.DIODE(_1422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3087__A1 (.DIODE(_1422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3271__A1 (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3224__A1 (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3215__A1 (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3206__A1 (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3197__A1 (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3178__A1 (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3169__A1 (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3160__A1 (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3151__A1 (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3090__A1 (.DIODE(_1425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3273__A1 (.DIODE(_1427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3226__A1 (.DIODE(_1427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3217__A1 (.DIODE(_1427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3208__A1 (.DIODE(_1427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3199__A1 (.DIODE(_1427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3180__A1 (.DIODE(_1427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3171__A1 (.DIODE(_1427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3162__A1 (.DIODE(_1427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3153__A1 (.DIODE(_1427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3093__A1 (.DIODE(_1427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3275__A1 (.DIODE(_1429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3228__A1 (.DIODE(_1429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3219__A1 (.DIODE(_1429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3210__A1 (.DIODE(_1429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3201__A1 (.DIODE(_1429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3182__A1 (.DIODE(_1429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3173__A1 (.DIODE(_1429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3164__A1 (.DIODE(_1429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3155__A1 (.DIODE(_1429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3096__A1 (.DIODE(_1429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3114__S (.DIODE(_1436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3112__S (.DIODE(_1436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3110__S (.DIODE(_1436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3108__S (.DIODE(_1436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3296__A0 (.DIODE(_1446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3287__A0 (.DIODE(_1446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3278__A0 (.DIODE(_1446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3260__A0 (.DIODE(_1446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3251__A0 (.DIODE(_1446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3242__A0 (.DIODE(_1446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3233__A0 (.DIODE(_1446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3186__A0 (.DIODE(_1446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3139__A0 (.DIODE(_1446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3127__A0 (.DIODE(_1446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3298__A0 (.DIODE(_1449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3289__A0 (.DIODE(_1449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3280__A0 (.DIODE(_1449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3262__A0 (.DIODE(_1449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3253__A0 (.DIODE(_1449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3244__A0 (.DIODE(_1449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3235__A0 (.DIODE(_1449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3188__A0 (.DIODE(_1449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3141__A0 (.DIODE(_1449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3130__A0 (.DIODE(_1449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3300__A0 (.DIODE(_1451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3291__A0 (.DIODE(_1451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3282__A0 (.DIODE(_1451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3264__A0 (.DIODE(_1451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3255__A0 (.DIODE(_1451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3246__A0 (.DIODE(_1451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3237__A0 (.DIODE(_1451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3190__A0 (.DIODE(_1451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3143__A0 (.DIODE(_1451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3133__A0 (.DIODE(_1451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3302__A0 (.DIODE(_1453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3293__A0 (.DIODE(_1453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3284__A0 (.DIODE(_1453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3266__A0 (.DIODE(_1453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3257__A0 (.DIODE(_1453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3248__A0 (.DIODE(_1453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3239__A0 (.DIODE(_1453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3192__A0 (.DIODE(_1453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3145__A0 (.DIODE(_1453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3136__A0 (.DIODE(_1453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4107__A (.DIODE(_1460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4062__A (.DIODE(_1460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3221__A (.DIODE(_1460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3212__B (.DIODE(_1460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3203__A (.DIODE(_1460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3194__B (.DIODE(_1460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3175__A (.DIODE(_1460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3166__B (.DIODE(_1460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3157__A (.DIODE(_1460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3148__A (.DIODE(_1460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4071__B (.DIODE(_1508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3385__B (.DIODE(_1508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3376__B (.DIODE(_1508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3348__B (.DIODE(_1508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3339__B (.DIODE(_1508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3317__B (.DIODE(_1508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3305__B (.DIODE(_1508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3277__B (.DIODE(_1508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3268__B (.DIODE(_1508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3232__B (.DIODE(_1508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3458__A1 (.DIODE(_1549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3449__A1 (.DIODE(_1549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3440__A1 (.DIODE(_1549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3404__A1 (.DIODE(_1549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3386__A1 (.DIODE(_1549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3377__A1 (.DIODE(_1549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3349__A1 (.DIODE(_1549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3340__A1 (.DIODE(_1549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3318__A1 (.DIODE(_1549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3306__A1 (.DIODE(_1549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3460__A1 (.DIODE(_1552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3451__A1 (.DIODE(_1552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3442__A1 (.DIODE(_1552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3406__A1 (.DIODE(_1552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3388__A1 (.DIODE(_1552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3379__A1 (.DIODE(_1552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3351__A1 (.DIODE(_1552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3342__A1 (.DIODE(_1552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3320__A1 (.DIODE(_1552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3309__A1 (.DIODE(_1552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3462__A1 (.DIODE(_1554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3453__A1 (.DIODE(_1554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3444__A1 (.DIODE(_1554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3408__A1 (.DIODE(_1554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3390__A1 (.DIODE(_1554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3381__A1 (.DIODE(_1554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3353__A1 (.DIODE(_1554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3344__A1 (.DIODE(_1554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3322__A1 (.DIODE(_1554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3312__A1 (.DIODE(_1554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3464__A1 (.DIODE(_1556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3455__A1 (.DIODE(_1556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3446__A1 (.DIODE(_1556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3410__A1 (.DIODE(_1556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3392__A1 (.DIODE(_1556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3383__A1 (.DIODE(_1556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3355__A1 (.DIODE(_1556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3346__A1 (.DIODE(_1556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3324__A1 (.DIODE(_1556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3315__A1 (.DIODE(_1556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3526__A0 (.DIODE(_1563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3517__A0 (.DIODE(_1563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3467__A0 (.DIODE(_1563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3431__A0 (.DIODE(_1563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3422__A0 (.DIODE(_1563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3413__A0 (.DIODE(_1563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3395__A0 (.DIODE(_1563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3368__A0 (.DIODE(_1563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3359__A0 (.DIODE(_1563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3328__A0 (.DIODE(_1563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3528__A0 (.DIODE(_1566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3519__A0 (.DIODE(_1566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3469__A0 (.DIODE(_1566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3433__A0 (.DIODE(_1566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3424__A0 (.DIODE(_1566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3415__A0 (.DIODE(_1566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3397__A0 (.DIODE(_1566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3370__A0 (.DIODE(_1566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3361__A0 (.DIODE(_1566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3331__A0 (.DIODE(_1566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3530__A0 (.DIODE(_1568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3521__A0 (.DIODE(_1568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3471__A0 (.DIODE(_1568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3435__A0 (.DIODE(_1568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3426__A0 (.DIODE(_1568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3417__A0 (.DIODE(_1568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3399__A0 (.DIODE(_1568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3372__A0 (.DIODE(_1568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3363__A0 (.DIODE(_1568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3334__A0 (.DIODE(_1568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3532__A0 (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3523__A0 (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3473__A0 (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3437__A0 (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3428__A0 (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3419__A0 (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3401__A0 (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3374__A0 (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3365__A0 (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3337__A0 (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3647__A1 (.DIODE(_1648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3629__A1 (.DIODE(_1648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3620__A1 (.DIODE(_1648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3611__A1 (.DIODE(_1648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3602__A1 (.DIODE(_1648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3557__A1 (.DIODE(_1648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3507__A1 (.DIODE(_1648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3498__A1 (.DIODE(_1648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3489__A1 (.DIODE(_1648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3477__A1 (.DIODE(_1648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3649__A1 (.DIODE(_1651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3631__A1 (.DIODE(_1651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3622__A1 (.DIODE(_1651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3613__A1 (.DIODE(_1651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3604__A1 (.DIODE(_1651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3559__A1 (.DIODE(_1651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3509__A1 (.DIODE(_1651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3500__A1 (.DIODE(_1651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3491__A1 (.DIODE(_1651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3480__A1 (.DIODE(_1651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3651__A1 (.DIODE(_1653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3633__A1 (.DIODE(_1653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3624__A1 (.DIODE(_1653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3615__A1 (.DIODE(_1653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3606__A1 (.DIODE(_1653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3561__A1 (.DIODE(_1653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3511__A1 (.DIODE(_1653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3502__A1 (.DIODE(_1653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3493__A1 (.DIODE(_1653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3483__A1 (.DIODE(_1653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3653__A1 (.DIODE(_1655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3635__A1 (.DIODE(_1655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3626__A1 (.DIODE(_1655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3617__A1 (.DIODE(_1655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3608__A1 (.DIODE(_1655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3563__A1 (.DIODE(_1655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3513__A1 (.DIODE(_1655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3504__A1 (.DIODE(_1655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3495__A1 (.DIODE(_1655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3486__A1 (.DIODE(_1655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3710__A0 (.DIODE(_1683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3692__A0 (.DIODE(_1683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3683__A0 (.DIODE(_1683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3638__A0 (.DIODE(_1683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3593__A0 (.DIODE(_1683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3584__A0 (.DIODE(_1683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3575__A0 (.DIODE(_1683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3566__A0 (.DIODE(_1683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3548__A0 (.DIODE(_1683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3536__A0 (.DIODE(_1683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3712__A0 (.DIODE(_1686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3694__A0 (.DIODE(_1686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3685__A0 (.DIODE(_1686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3640__A0 (.DIODE(_1686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3595__A0 (.DIODE(_1686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3586__A0 (.DIODE(_1686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3577__A0 (.DIODE(_1686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3568__A0 (.DIODE(_1686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3550__A0 (.DIODE(_1686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3539__A0 (.DIODE(_1686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3714__A0 (.DIODE(_1688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3696__A0 (.DIODE(_1688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3687__A0 (.DIODE(_1688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3642__A0 (.DIODE(_1688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3597__A0 (.DIODE(_1688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3588__A0 (.DIODE(_1688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3579__A0 (.DIODE(_1688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3570__A0 (.DIODE(_1688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3552__A0 (.DIODE(_1688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3542__A0 (.DIODE(_1688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3716__A0 (.DIODE(_1690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3698__A0 (.DIODE(_1690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3689__A0 (.DIODE(_1690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3644__A0 (.DIODE(_1690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3599__A0 (.DIODE(_1690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3590__A0 (.DIODE(_1690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3581__A0 (.DIODE(_1690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3572__A0 (.DIODE(_1690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3554__A0 (.DIODE(_1690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3545__A0 (.DIODE(_1690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4117__A0 (.DIODE(_1797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4108__A0 (.DIODE(_1797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4099__A0 (.DIODE(_1797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4090__A0 (.DIODE(_1797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4081__A0 (.DIODE(_1797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4063__A0 (.DIODE(_1797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4054__A0 (.DIODE(_1797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3759__A0 (.DIODE(_1797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3750__A0 (.DIODE(_1797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3738__A0 (.DIODE(_1797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4119__A0 (.DIODE(_1800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4110__A0 (.DIODE(_1800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4101__A0 (.DIODE(_1800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4092__A0 (.DIODE(_1800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4083__A0 (.DIODE(_1800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4065__A0 (.DIODE(_1800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4056__A0 (.DIODE(_1800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3761__A0 (.DIODE(_1800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3752__A0 (.DIODE(_1800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3741__A0 (.DIODE(_1800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4121__A0 (.DIODE(_1802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4112__A0 (.DIODE(_1802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4103__A0 (.DIODE(_1802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4094__A0 (.DIODE(_1802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4085__A0 (.DIODE(_1802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4067__A0 (.DIODE(_1802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4058__A0 (.DIODE(_1802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3763__A0 (.DIODE(_1802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3754__A0 (.DIODE(_1802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3744__A0 (.DIODE(_1802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4123__A0 (.DIODE(_1804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4114__A0 (.DIODE(_1804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4105__A0 (.DIODE(_1804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4096__A0 (.DIODE(_1804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4087__A0 (.DIODE(_1804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4069__A0 (.DIODE(_1804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4060__A0 (.DIODE(_1804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3765__A0 (.DIODE(_1804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3756__A0 (.DIODE(_1804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3747__A0 (.DIODE(_1804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3955__B1 (.DIODE(_1824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3915__C1 (.DIODE(_1824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3912__C1 (.DIODE(_1824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3904__C1 (.DIODE(_1824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3817__A (.DIODE(_1824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3795__A (.DIODE(_1824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3791__A (.DIODE(_1824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3787__B1 (.DIODE(_1824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3786__A (.DIODE(_1824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3783__B (.DIODE(_1824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3893__C1 (.DIODE(_1843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3890__C1 (.DIODE(_1843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3887__C1 (.DIODE(_1843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3884__C1 (.DIODE(_1843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3878__C1 (.DIODE(_1843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3875__C1 (.DIODE(_1843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3872__C1 (.DIODE(_1843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3824__C1 (.DIODE(_1843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3821__C1 (.DIODE(_1843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3808__C1 (.DIODE(_1843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4042__D_N (.DIODE(_1847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4023__B (.DIODE(_1847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3998__A2 (.DIODE(_1847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3997__A (.DIODE(_1847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3982__A1 (.DIODE(_1847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3979__D (.DIODE(_1847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3962__A1 (.DIODE(_1847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3911__A (.DIODE(_1847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3880__B (.DIODE(_1847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3813__B2 (.DIODE(_1847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4042__A (.DIODE(_1848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4032__A2 (.DIODE(_1848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4023__A (.DIODE(_1848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3997__C_N (.DIODE(_1848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3986__A1 (.DIODE(_1848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3979__C (.DIODE(_1848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3965__A1 (.DIODE(_1848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3914__A (.DIODE(_1848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3880__A_N (.DIODE(_1848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3816__A0 (.DIODE(_1848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4096__S (.DIODE(_2043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4094__S (.DIODE(_2043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4092__S (.DIODE(_2043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4090__S (.DIODE(_2043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4123__S (.DIODE(_2058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4121__S (.DIODE(_2058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4119__S (.DIODE(_2058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4117__S (.DIODE(_2058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4141__S (.DIODE(_2068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4139__S (.DIODE(_2068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4137__S (.DIODE(_2068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4135__S (.DIODE(_2068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4162__S (.DIODE(_2073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4160__S (.DIODE(_2073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4158__S (.DIODE(_2073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4156__S (.DIODE(_2073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4154__S (.DIODE(_2073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4152__S (.DIODE(_2073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4150__S (.DIODE(_2073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4148__S (.DIODE(_2073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4146__S (.DIODE(_2073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4144__S (.DIODE(_2073_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(io_in[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(io_in[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(io_in[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(io_in[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(oram_value[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(oram_value[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(oram_value[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(oram_value[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(oram_value[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(oram_value[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(oram_value[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(oram_value[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(oram_value[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(oram_value[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(oram_value[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA__2896__A1 (.DIODE(\tms1x00.RAM[0][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2253__A0 (.DIODE(\tms1x00.RAM[0][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2902__A1 (.DIODE(\tms1x00.RAM[0][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2472__A0 (.DIODE(\tms1x00.RAM[0][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3991__A1 (.DIODE(\tms1x00.Y[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3853__A (.DIODE(\tms1x00.Y[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3848__C (.DIODE(\tms1x00.Y[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3843__C (.DIODE(\tms1x00.Y[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3840__C_N (.DIODE(\tms1x00.Y[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3834__A_N (.DIODE(\tms1x00.Y[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2104__A (.DIODE(\tms1x00.Y[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3980__A (.DIODE(\tms1x00.ins_in[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3959__A1 (.DIODE(\tms1x00.ins_in[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3908__C (.DIODE(\tms1x00.ins_in[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3808__A1 (.DIODE(\tms1x00.ins_in[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2302__A (.DIODE(\tms1x00.ins_in[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2142__A_N (.DIODE(\tms1x00.ins_in[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2125__A (.DIODE(\tms1x00.ins_in[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2882__B (.DIODE(\tms1x00.ram_addr_buff[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2820__C_N (.DIODE(\tms1x00.ram_addr_buff[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2787__B (.DIODE(\tms1x00.ram_addr_buff[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2681__A (.DIODE(\tms1x00.ram_addr_buff[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2625__A (.DIODE(\tms1x00.ram_addr_buff[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2314__B (.DIODE(\tms1x00.ram_addr_buff[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2101__A (.DIODE(\tms1x00.ram_addr_buff[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3230__A (.DIODE(\tms1x00.ram_addr_buff[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2785__A (.DIODE(\tms1x00.ram_addr_buff[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2715__C_N (.DIODE(\tms1x00.ram_addr_buff[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2678__A (.DIODE(\tms1x00.ram_addr_buff[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2639__A (.DIODE(\tms1x00.ram_addr_buff[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2622__C (.DIODE(\tms1x00.ram_addr_buff[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2310__A_N (.DIODE(\tms1x00.ram_addr_buff[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2111__A (.DIODE(\tms1x00.ram_addr_buff[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3230__C_N (.DIODE(\tms1x00.ram_addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2785__B (.DIODE(\tms1x00.ram_addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2715__A (.DIODE(\tms1x00.ram_addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2678__B (.DIODE(\tms1x00.ram_addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2639__B (.DIODE(\tms1x00.ram_addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2622__A_N (.DIODE(\tms1x00.ram_addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2310__B (.DIODE(\tms1x00.ram_addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2114__A (.DIODE(\tms1x00.ram_addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3230__B (.DIODE(\tms1x00.ram_addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2935__C (.DIODE(\tms1x00.ram_addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2785__C (.DIODE(\tms1x00.ram_addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2715__B (.DIODE(\tms1x00.ram_addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2678__C_N (.DIODE(\tms1x00.ram_addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2640__A (.DIODE(\tms1x00.ram_addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2622__B (.DIODE(\tms1x00.ram_addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2310__C (.DIODE(\tms1x00.ram_addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2117__A (.DIODE(\tms1x00.ram_addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_wb_clk_i_A (.DIODE(wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(wb_rst_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(wbs_adr_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(wbs_adr_i[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(wbs_adr_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(wbs_adr_i[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(wbs_adr_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(wbs_adr_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(wbs_adr_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(wbs_adr_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(wbs_adr_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(wbs_adr_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(wbs_adr_i[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(wbs_cyc_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(wbs_dat_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(wbs_stb_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(wbs_we_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__3789__A0 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__4844__A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__4042__B (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__3973__C (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__3781__A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__2303__B (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__2144__B (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__2093__A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__4845__A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__4846__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__2702__A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__4847__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__4848__A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__4849__A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__4850__A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__4851__A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__4852__A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__4853__A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__2121__B (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__2089__B (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__2120__A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__2089__C (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_output32_A (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__3884__A1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_output34_A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__3890__A1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_output35_A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__3893__A1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_output36_A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__3896__A1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_output37_A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__3981__A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__3974__A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__3785__B (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__3784__A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__3783__A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__2143__B (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__2128__B (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__2094__A_N (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_output38_A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__3973__B (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__3797__A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__3785__A_N (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__3784__B (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__2143__C_N (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__2128__C (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__2095__A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_output39_A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__3973__A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__3785__C (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__2144__A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__2128__A_N (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__2094__B (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_output40_A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__2138__B1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_output41_A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__3827__B1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_output42_A (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__3831__B1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_output43_A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__3835__B1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_output44_A (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__3841__B1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_output45_A (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__3844__B1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_output46_A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__3849__B1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_output47_A (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__3854__B1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_output48_A (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__3858__B1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_output49_A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__3860__B1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_output50_A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__3862__B1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_output51_A (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__3864__B1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_output52_A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__3868__B1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_output53_A (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__3871__B1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_output54_A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__3874__B1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_output55_A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__3877__B1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_output56_A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__2703__A0 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_output66_A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_output67_A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_output68_A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_output69_A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_output70_A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_output71_A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_output72_A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_output73_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_output74_A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_output75_A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__4724__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4725__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4660__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4665__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4664__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4662__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4667__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4661__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4668__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4659__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4577__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4694__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4775__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4663__CLK (.DIODE(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4680__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4722__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4446__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4503__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4475__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4504__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4419__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4454__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4418__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4450__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4463__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4448__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4449__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4452__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4453__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4445__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4721__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4731__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4685__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4679__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4492__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4687__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4677__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4686__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4683__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4509__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4479__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4507__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4675__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4684__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4674__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4682__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4676__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4379__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4595__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4465__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4378__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4427__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4441__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4440__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4423__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4429__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4430__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4657__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4431__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4416__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4376__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4417__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4464__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4428__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4377__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4548__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4547__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4543__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4550__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4551__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4466__CLK (.DIODE(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4557__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4555__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4279__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4192__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4277__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4199__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4202__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4373__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4200__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4336__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4372__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4193__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4375__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4335__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4224__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4227__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4399__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4220__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4286__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4290__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4288__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4285__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4284__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4177__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4280__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4176__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4175__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4206__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4204__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4283__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4207__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4499__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4281__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4501__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4493__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4205__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4525__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4296__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4300__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4299__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4294__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4306__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4313__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4338__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4307__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4337__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4303__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4368__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4332__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4226__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4339__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4333__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4374__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4201__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4178__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4287__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4282__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4291__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4295__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4298__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4591__CLK (.DIODE(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4197__CLK (.DIODE(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4196__CLK (.DIODE(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4592__CLK (.DIODE(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4626__CLK (.DIODE(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4590__CLK (.DIODE(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4593__CLK (.DIODE(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4542__CLK (.DIODE(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4541__CLK (.DIODE(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4644__CLK (.DIODE(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4641__CLK (.DIODE(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4649__CLK (.DIODE(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4645__CLK (.DIODE(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4586__CLK (.DIODE(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4317__CLK (.DIODE(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4249__CLK (.DIODE(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4785__CLK (.DIODE(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4356__CLK (.DIODE(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4784__CLK (.DIODE(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4637__CLK (.DIODE(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4246__CLK (.DIODE(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4636__CLK (.DIODE(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4247__CLK (.DIODE(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4403__CLK (.DIODE(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4237__CLK (.DIODE(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4238__CLK (.DIODE(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4407__CLK (.DIODE(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4415__CLK (.DIODE(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4383__CLK (.DIODE(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4601__CLK (.DIODE(clknet_leaf_36_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4561__CLK (.DIODE(clknet_leaf_36_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4599__CLK (.DIODE(clknet_leaf_36_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4624__CLK (.DIODE(clknet_leaf_36_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4562__CLK (.DIODE(clknet_leaf_36_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4539__CLK (.DIODE(clknet_leaf_36_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4646__CLK (.DIODE(clknet_leaf_36_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4540__CLK (.DIODE(clknet_leaf_36_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4588__CLK (.DIODE(clknet_leaf_36_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4625__CLK (.DIODE(clknet_leaf_36_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4634__CLK (.DIODE(clknet_leaf_36_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4635__CLK (.DIODE(clknet_leaf_36_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4587__CLK (.DIODE(clknet_leaf_36_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4623__CLK (.DIODE(clknet_leaf_36_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4589__CLK (.DIODE(clknet_leaf_36_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4632__CLK (.DIODE(clknet_leaf_36_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4633__CLK (.DIODE(clknet_leaf_36_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4316__CLK (.DIODE(clknet_leaf_36_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4327__CLK (.DIODE(clknet_leaf_38_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4270__CLK (.DIODE(clknet_leaf_38_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4272__CLK (.DIODE(clknet_leaf_38_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4266__CLK (.DIODE(clknet_leaf_38_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4274__CLK (.DIODE(clknet_leaf_38_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4262__CLK (.DIODE(clknet_leaf_38_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4273__CLK (.DIODE(clknet_leaf_38_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4269__CLK (.DIODE(clknet_leaf_38_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4261__CLK (.DIODE(clknet_leaf_38_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4260__CLK (.DIODE(clknet_leaf_38_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4264__CLK (.DIODE(clknet_leaf_38_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4265__CLK (.DIODE(clknet_leaf_38_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4604__CLK (.DIODE(clknet_leaf_38_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4435__CLK (.DIODE(clknet_leaf_38_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4434__CLK (.DIODE(clknet_leaf_38_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4268__CLK (.DIODE(clknet_leaf_38_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_42_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_41_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_40_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_39_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_38_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_37_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__decap_4 FILLER_0_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_591 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_618 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_678 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_532 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_522 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_826 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_731 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_704 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_672 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_732 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_760 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_508 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_471 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_678 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_647 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_760 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_616 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_732 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_732 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_56 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_22 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_471 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_534 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_820 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_663 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_420 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_836 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_663 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_646 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_508 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_823 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_700 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_704 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_471 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_841 ();
 assign io_oeb[0] = net125;
 assign io_oeb[10] = net83;
 assign io_oeb[11] = net84;
 assign io_oeb[12] = net85;
 assign io_oeb[13] = net86;
 assign io_oeb[14] = net87;
 assign io_oeb[15] = net88;
 assign io_oeb[16] = net89;
 assign io_oeb[17] = net90;
 assign io_oeb[18] = net91;
 assign io_oeb[19] = net92;
 assign io_oeb[1] = net126;
 assign io_oeb[20] = net93;
 assign io_oeb[21] = net94;
 assign io_oeb[22] = net95;
 assign io_oeb[23] = net96;
 assign io_oeb[24] = net97;
 assign io_oeb[25] = net98;
 assign io_oeb[26] = net99;
 assign io_oeb[27] = net100;
 assign io_oeb[28] = net101;
 assign io_oeb[29] = net102;
 assign io_oeb[2] = net127;
 assign io_oeb[30] = net103;
 assign io_oeb[31] = net104;
 assign io_oeb[32] = net105;
 assign io_oeb[33] = net106;
 assign io_oeb[34] = net107;
 assign io_oeb[35] = net108;
 assign io_oeb[36] = net109;
 assign io_oeb[37] = net110;
 assign io_oeb[3] = net128;
 assign io_oeb[4] = net129;
 assign io_oeb[5] = net78;
 assign io_oeb[6] = net79;
 assign io_oeb[7] = net80;
 assign io_oeb[8] = net81;
 assign io_oeb[9] = net82;
 assign io_out[0] = net111;
 assign io_out[1] = net112;
 assign io_out[2] = net113;
 assign io_out[34] = net121;
 assign io_out[35] = net122;
 assign io_out[36] = net123;
 assign io_out[3] = net114;
 assign io_out[4] = net115;
 assign io_out[5] = net116;
 assign io_out[6] = net117;
 assign io_out[7] = net118;
 assign io_out[8] = net119;
 assign io_out[9] = net120;
 assign oram_addr[8] = net124;
 assign ram_wmask[0] = net130;
 assign ram_wmask[1] = net131;
 assign ram_wmask[2] = net132;
 assign ram_wmask[3] = net133;
endmodule

