magic
tech sky130B
magscale 1 2
timestamp 1671528632
<< obsli1 >>
rect 1104 2159 78844 47345
<< obsm1 >>
rect 934 1504 79014 47728
<< metal2 >>
rect 3514 49200 3570 50000
rect 4158 49200 4214 50000
rect 4802 49200 4858 50000
rect 5446 49200 5502 50000
rect 6090 49200 6146 50000
rect 6734 49200 6790 50000
rect 7378 49200 7434 50000
rect 8022 49200 8078 50000
rect 8666 49200 8722 50000
rect 9310 49200 9366 50000
rect 9954 49200 10010 50000
rect 10598 49200 10654 50000
rect 11242 49200 11298 50000
rect 11886 49200 11942 50000
rect 12530 49200 12586 50000
rect 13174 49200 13230 50000
rect 13818 49200 13874 50000
rect 14462 49200 14518 50000
rect 15106 49200 15162 50000
rect 15750 49200 15806 50000
rect 16394 49200 16450 50000
rect 17038 49200 17094 50000
rect 17682 49200 17738 50000
rect 18326 49200 18382 50000
rect 18970 49200 19026 50000
rect 19614 49200 19670 50000
rect 20258 49200 20314 50000
rect 20902 49200 20958 50000
rect 21546 49200 21602 50000
rect 22190 49200 22246 50000
rect 22834 49200 22890 50000
rect 23478 49200 23534 50000
rect 24122 49200 24178 50000
rect 24766 49200 24822 50000
rect 25410 49200 25466 50000
rect 26054 49200 26110 50000
rect 26698 49200 26754 50000
rect 27342 49200 27398 50000
rect 27986 49200 28042 50000
rect 28630 49200 28686 50000
rect 29274 49200 29330 50000
rect 29918 49200 29974 50000
rect 30562 49200 30618 50000
rect 31206 49200 31262 50000
rect 31850 49200 31906 50000
rect 32494 49200 32550 50000
rect 33138 49200 33194 50000
rect 33782 49200 33838 50000
rect 34426 49200 34482 50000
rect 35070 49200 35126 50000
rect 35714 49200 35770 50000
rect 36358 49200 36414 50000
rect 37002 49200 37058 50000
rect 37646 49200 37702 50000
rect 38290 49200 38346 50000
rect 38934 49200 38990 50000
rect 39578 49200 39634 50000
rect 40222 49200 40278 50000
rect 40866 49200 40922 50000
rect 41510 49200 41566 50000
rect 42154 49200 42210 50000
rect 42798 49200 42854 50000
rect 43442 49200 43498 50000
rect 44086 49200 44142 50000
rect 44730 49200 44786 50000
rect 45374 49200 45430 50000
rect 46018 49200 46074 50000
rect 46662 49200 46718 50000
rect 47306 49200 47362 50000
rect 47950 49200 48006 50000
rect 48594 49200 48650 50000
rect 49238 49200 49294 50000
rect 49882 49200 49938 50000
rect 50526 49200 50582 50000
rect 51170 49200 51226 50000
rect 51814 49200 51870 50000
rect 52458 49200 52514 50000
rect 53102 49200 53158 50000
rect 53746 49200 53802 50000
rect 54390 49200 54446 50000
rect 55034 49200 55090 50000
rect 55678 49200 55734 50000
rect 56322 49200 56378 50000
rect 56966 49200 57022 50000
rect 57610 49200 57666 50000
rect 58254 49200 58310 50000
rect 58898 49200 58954 50000
rect 59542 49200 59598 50000
rect 60186 49200 60242 50000
rect 60830 49200 60886 50000
rect 61474 49200 61530 50000
rect 62118 49200 62174 50000
rect 62762 49200 62818 50000
rect 63406 49200 63462 50000
rect 64050 49200 64106 50000
rect 64694 49200 64750 50000
rect 65338 49200 65394 50000
rect 65982 49200 66038 50000
rect 66626 49200 66682 50000
rect 67270 49200 67326 50000
rect 67914 49200 67970 50000
rect 68558 49200 68614 50000
rect 69202 49200 69258 50000
rect 69846 49200 69902 50000
rect 70490 49200 70546 50000
rect 71134 49200 71190 50000
rect 71778 49200 71834 50000
rect 72422 49200 72478 50000
rect 73066 49200 73122 50000
rect 73710 49200 73766 50000
rect 74354 49200 74410 50000
rect 74998 49200 75054 50000
rect 75642 49200 75698 50000
rect 76286 49200 76342 50000
rect 938 0 994 800
rect 2410 0 2466 800
rect 3882 0 3938 800
rect 5354 0 5410 800
rect 6826 0 6882 800
rect 8298 0 8354 800
rect 9770 0 9826 800
rect 11242 0 11298 800
rect 12714 0 12770 800
rect 14186 0 14242 800
rect 15658 0 15714 800
rect 17130 0 17186 800
rect 18602 0 18658 800
rect 20074 0 20130 800
rect 21546 0 21602 800
rect 23018 0 23074 800
rect 24490 0 24546 800
rect 25962 0 26018 800
rect 27434 0 27490 800
rect 28906 0 28962 800
rect 30378 0 30434 800
rect 31850 0 31906 800
rect 33322 0 33378 800
rect 34794 0 34850 800
rect 36266 0 36322 800
rect 37738 0 37794 800
rect 39210 0 39266 800
rect 40682 0 40738 800
rect 42154 0 42210 800
rect 43626 0 43682 800
rect 45098 0 45154 800
rect 46570 0 46626 800
rect 48042 0 48098 800
rect 49514 0 49570 800
rect 50986 0 51042 800
rect 52458 0 52514 800
rect 53930 0 53986 800
rect 55402 0 55458 800
rect 56874 0 56930 800
rect 58346 0 58402 800
rect 59818 0 59874 800
rect 61290 0 61346 800
rect 62762 0 62818 800
rect 64234 0 64290 800
rect 65706 0 65762 800
rect 67178 0 67234 800
rect 68650 0 68706 800
rect 70122 0 70178 800
rect 71594 0 71650 800
rect 73066 0 73122 800
rect 74538 0 74594 800
rect 76010 0 76066 800
rect 77482 0 77538 800
rect 78954 0 79010 800
<< obsm2 >>
rect 940 49144 3458 49314
rect 3626 49144 4102 49314
rect 4270 49144 4746 49314
rect 4914 49144 5390 49314
rect 5558 49144 6034 49314
rect 6202 49144 6678 49314
rect 6846 49144 7322 49314
rect 7490 49144 7966 49314
rect 8134 49144 8610 49314
rect 8778 49144 9254 49314
rect 9422 49144 9898 49314
rect 10066 49144 10542 49314
rect 10710 49144 11186 49314
rect 11354 49144 11830 49314
rect 11998 49144 12474 49314
rect 12642 49144 13118 49314
rect 13286 49144 13762 49314
rect 13930 49144 14406 49314
rect 14574 49144 15050 49314
rect 15218 49144 15694 49314
rect 15862 49144 16338 49314
rect 16506 49144 16982 49314
rect 17150 49144 17626 49314
rect 17794 49144 18270 49314
rect 18438 49144 18914 49314
rect 19082 49144 19558 49314
rect 19726 49144 20202 49314
rect 20370 49144 20846 49314
rect 21014 49144 21490 49314
rect 21658 49144 22134 49314
rect 22302 49144 22778 49314
rect 22946 49144 23422 49314
rect 23590 49144 24066 49314
rect 24234 49144 24710 49314
rect 24878 49144 25354 49314
rect 25522 49144 25998 49314
rect 26166 49144 26642 49314
rect 26810 49144 27286 49314
rect 27454 49144 27930 49314
rect 28098 49144 28574 49314
rect 28742 49144 29218 49314
rect 29386 49144 29862 49314
rect 30030 49144 30506 49314
rect 30674 49144 31150 49314
rect 31318 49144 31794 49314
rect 31962 49144 32438 49314
rect 32606 49144 33082 49314
rect 33250 49144 33726 49314
rect 33894 49144 34370 49314
rect 34538 49144 35014 49314
rect 35182 49144 35658 49314
rect 35826 49144 36302 49314
rect 36470 49144 36946 49314
rect 37114 49144 37590 49314
rect 37758 49144 38234 49314
rect 38402 49144 38878 49314
rect 39046 49144 39522 49314
rect 39690 49144 40166 49314
rect 40334 49144 40810 49314
rect 40978 49144 41454 49314
rect 41622 49144 42098 49314
rect 42266 49144 42742 49314
rect 42910 49144 43386 49314
rect 43554 49144 44030 49314
rect 44198 49144 44674 49314
rect 44842 49144 45318 49314
rect 45486 49144 45962 49314
rect 46130 49144 46606 49314
rect 46774 49144 47250 49314
rect 47418 49144 47894 49314
rect 48062 49144 48538 49314
rect 48706 49144 49182 49314
rect 49350 49144 49826 49314
rect 49994 49144 50470 49314
rect 50638 49144 51114 49314
rect 51282 49144 51758 49314
rect 51926 49144 52402 49314
rect 52570 49144 53046 49314
rect 53214 49144 53690 49314
rect 53858 49144 54334 49314
rect 54502 49144 54978 49314
rect 55146 49144 55622 49314
rect 55790 49144 56266 49314
rect 56434 49144 56910 49314
rect 57078 49144 57554 49314
rect 57722 49144 58198 49314
rect 58366 49144 58842 49314
rect 59010 49144 59486 49314
rect 59654 49144 60130 49314
rect 60298 49144 60774 49314
rect 60942 49144 61418 49314
rect 61586 49144 62062 49314
rect 62230 49144 62706 49314
rect 62874 49144 63350 49314
rect 63518 49144 63994 49314
rect 64162 49144 64638 49314
rect 64806 49144 65282 49314
rect 65450 49144 65926 49314
rect 66094 49144 66570 49314
rect 66738 49144 67214 49314
rect 67382 49144 67858 49314
rect 68026 49144 68502 49314
rect 68670 49144 69146 49314
rect 69314 49144 69790 49314
rect 69958 49144 70434 49314
rect 70602 49144 71078 49314
rect 71246 49144 71722 49314
rect 71890 49144 72366 49314
rect 72534 49144 73010 49314
rect 73178 49144 73654 49314
rect 73822 49144 74298 49314
rect 74466 49144 74942 49314
rect 75110 49144 75586 49314
rect 75754 49144 76230 49314
rect 76398 49144 79008 49314
rect 940 856 79008 49144
rect 1050 800 2354 856
rect 2522 800 3826 856
rect 3994 800 5298 856
rect 5466 800 6770 856
rect 6938 800 8242 856
rect 8410 800 9714 856
rect 9882 800 11186 856
rect 11354 800 12658 856
rect 12826 800 14130 856
rect 14298 800 15602 856
rect 15770 800 17074 856
rect 17242 800 18546 856
rect 18714 800 20018 856
rect 20186 800 21490 856
rect 21658 800 22962 856
rect 23130 800 24434 856
rect 24602 800 25906 856
rect 26074 800 27378 856
rect 27546 800 28850 856
rect 29018 800 30322 856
rect 30490 800 31794 856
rect 31962 800 33266 856
rect 33434 800 34738 856
rect 34906 800 36210 856
rect 36378 800 37682 856
rect 37850 800 39154 856
rect 39322 800 40626 856
rect 40794 800 42098 856
rect 42266 800 43570 856
rect 43738 800 45042 856
rect 45210 800 46514 856
rect 46682 800 47986 856
rect 48154 800 49458 856
rect 49626 800 50930 856
rect 51098 800 52402 856
rect 52570 800 53874 856
rect 54042 800 55346 856
rect 55514 800 56818 856
rect 56986 800 58290 856
rect 58458 800 59762 856
rect 59930 800 61234 856
rect 61402 800 62706 856
rect 62874 800 64178 856
rect 64346 800 65650 856
rect 65818 800 67122 856
rect 67290 800 68594 856
rect 68762 800 70066 856
rect 70234 800 71538 856
rect 71706 800 73010 856
rect 73178 800 74482 856
rect 74650 800 75954 856
rect 76122 800 77426 856
rect 77594 800 78898 856
<< metal3 >>
rect 0 47200 800 47320
rect 0 46112 800 46232
rect 0 45024 800 45144
rect 0 43936 800 44056
rect 0 42848 800 42968
rect 0 41760 800 41880
rect 0 40672 800 40792
rect 0 39584 800 39704
rect 0 38496 800 38616
rect 0 37408 800 37528
rect 0 36320 800 36440
rect 0 35232 800 35352
rect 0 34144 800 34264
rect 0 33056 800 33176
rect 0 31968 800 32088
rect 0 30880 800 31000
rect 0 29792 800 29912
rect 0 28704 800 28824
rect 0 27616 800 27736
rect 0 26528 800 26648
rect 0 25440 800 25560
rect 0 24352 800 24472
rect 0 23264 800 23384
rect 0 22176 800 22296
rect 0 21088 800 21208
rect 0 20000 800 20120
rect 0 18912 800 19032
rect 0 17824 800 17944
rect 0 16736 800 16856
rect 0 15648 800 15768
rect 0 14560 800 14680
rect 0 13472 800 13592
rect 0 12384 800 12504
rect 0 11296 800 11416
rect 0 10208 800 10328
rect 0 9120 800 9240
rect 0 8032 800 8152
rect 0 6944 800 7064
rect 0 5856 800 5976
rect 0 4768 800 4888
rect 0 3680 800 3800
rect 0 2592 800 2712
<< obsm3 >>
rect 880 47120 78279 47361
rect 800 46312 78279 47120
rect 880 46032 78279 46312
rect 800 45224 78279 46032
rect 880 44944 78279 45224
rect 800 44136 78279 44944
rect 880 43856 78279 44136
rect 800 43048 78279 43856
rect 880 42768 78279 43048
rect 800 41960 78279 42768
rect 880 41680 78279 41960
rect 800 40872 78279 41680
rect 880 40592 78279 40872
rect 800 39784 78279 40592
rect 880 39504 78279 39784
rect 800 38696 78279 39504
rect 880 38416 78279 38696
rect 800 37608 78279 38416
rect 880 37328 78279 37608
rect 800 36520 78279 37328
rect 880 36240 78279 36520
rect 800 35432 78279 36240
rect 880 35152 78279 35432
rect 800 34344 78279 35152
rect 880 34064 78279 34344
rect 800 33256 78279 34064
rect 880 32976 78279 33256
rect 800 32168 78279 32976
rect 880 31888 78279 32168
rect 800 31080 78279 31888
rect 880 30800 78279 31080
rect 800 29992 78279 30800
rect 880 29712 78279 29992
rect 800 28904 78279 29712
rect 880 28624 78279 28904
rect 800 27816 78279 28624
rect 880 27536 78279 27816
rect 800 26728 78279 27536
rect 880 26448 78279 26728
rect 800 25640 78279 26448
rect 880 25360 78279 25640
rect 800 24552 78279 25360
rect 880 24272 78279 24552
rect 800 23464 78279 24272
rect 880 23184 78279 23464
rect 800 22376 78279 23184
rect 880 22096 78279 22376
rect 800 21288 78279 22096
rect 880 21008 78279 21288
rect 800 20200 78279 21008
rect 880 19920 78279 20200
rect 800 19112 78279 19920
rect 880 18832 78279 19112
rect 800 18024 78279 18832
rect 880 17744 78279 18024
rect 800 16936 78279 17744
rect 880 16656 78279 16936
rect 800 15848 78279 16656
rect 880 15568 78279 15848
rect 800 14760 78279 15568
rect 880 14480 78279 14760
rect 800 13672 78279 14480
rect 880 13392 78279 13672
rect 800 12584 78279 13392
rect 880 12304 78279 12584
rect 800 11496 78279 12304
rect 880 11216 78279 11496
rect 800 10408 78279 11216
rect 880 10128 78279 10408
rect 800 9320 78279 10128
rect 880 9040 78279 9320
rect 800 8232 78279 9040
rect 880 7952 78279 8232
rect 800 7144 78279 7952
rect 880 6864 78279 7144
rect 800 6056 78279 6864
rect 880 5776 78279 6056
rect 800 4968 78279 5776
rect 880 4688 78279 4968
rect 800 3880 78279 4688
rect 880 3600 78279 3880
rect 800 2792 78279 3600
rect 880 2512 78279 2792
rect 800 2143 78279 2512
<< metal4 >>
rect 4208 2128 4528 47376
rect 19568 2128 19888 47376
rect 34928 2128 35248 47376
rect 50288 2128 50608 47376
rect 65648 2128 65968 47376
<< obsm4 >>
rect 11099 5883 19488 45661
rect 19968 5883 34848 45661
rect 35328 5883 50208 45661
rect 50688 5883 65568 45661
rect 66048 5883 67469 45661
<< labels >>
rlabel metal2 s 3514 49200 3570 50000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 22834 49200 22890 50000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 24766 49200 24822 50000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 26698 49200 26754 50000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 28630 49200 28686 50000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 30562 49200 30618 50000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 32494 49200 32550 50000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 34426 49200 34482 50000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 36358 49200 36414 50000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 38290 49200 38346 50000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 40222 49200 40278 50000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 5446 49200 5502 50000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 42154 49200 42210 50000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 44086 49200 44142 50000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 46018 49200 46074 50000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 47950 49200 48006 50000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 49882 49200 49938 50000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 51814 49200 51870 50000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 53746 49200 53802 50000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 55678 49200 55734 50000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 57610 49200 57666 50000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 59542 49200 59598 50000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 7378 49200 7434 50000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 61474 49200 61530 50000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 63406 49200 63462 50000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 65338 49200 65394 50000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 67270 49200 67326 50000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 69202 49200 69258 50000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 71134 49200 71190 50000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 73066 49200 73122 50000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 74998 49200 75054 50000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 9310 49200 9366 50000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 11242 49200 11298 50000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 13174 49200 13230 50000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 15106 49200 15162 50000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 17038 49200 17094 50000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 18970 49200 19026 50000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 20902 49200 20958 50000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 4158 49200 4214 50000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 23478 49200 23534 50000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 25410 49200 25466 50000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 27342 49200 27398 50000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 29274 49200 29330 50000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 31206 49200 31262 50000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 33138 49200 33194 50000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 35070 49200 35126 50000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 37002 49200 37058 50000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 38934 49200 38990 50000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 40866 49200 40922 50000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 6090 49200 6146 50000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 42798 49200 42854 50000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 44730 49200 44786 50000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 46662 49200 46718 50000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 48594 49200 48650 50000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 50526 49200 50582 50000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 52458 49200 52514 50000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 54390 49200 54446 50000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 56322 49200 56378 50000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 58254 49200 58310 50000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 60186 49200 60242 50000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 8022 49200 8078 50000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 62118 49200 62174 50000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 64050 49200 64106 50000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 65982 49200 66038 50000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 67914 49200 67970 50000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 69846 49200 69902 50000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 71778 49200 71834 50000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 73710 49200 73766 50000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 75642 49200 75698 50000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 9954 49200 10010 50000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 11886 49200 11942 50000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 13818 49200 13874 50000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 15750 49200 15806 50000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 17682 49200 17738 50000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 19614 49200 19670 50000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 21546 49200 21602 50000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 4802 49200 4858 50000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 24122 49200 24178 50000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 26054 49200 26110 50000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 27986 49200 28042 50000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 29918 49200 29974 50000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 31850 49200 31906 50000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 33782 49200 33838 50000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 35714 49200 35770 50000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 37646 49200 37702 50000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 39578 49200 39634 50000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 41510 49200 41566 50000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 6734 49200 6790 50000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 43442 49200 43498 50000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 45374 49200 45430 50000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 47306 49200 47362 50000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 49238 49200 49294 50000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 51170 49200 51226 50000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 53102 49200 53158 50000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 55034 49200 55090 50000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 56966 49200 57022 50000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 58898 49200 58954 50000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 60830 49200 60886 50000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 8666 49200 8722 50000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 62762 49200 62818 50000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 64694 49200 64750 50000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 66626 49200 66682 50000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 68558 49200 68614 50000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 70490 49200 70546 50000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 72422 49200 72478 50000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 74354 49200 74410 50000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 76286 49200 76342 50000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 10598 49200 10654 50000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 12530 49200 12586 50000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 14462 49200 14518 50000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 16394 49200 16450 50000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 18326 49200 18382 50000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 20258 49200 20314 50000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 22190 49200 22246 50000 6 io_out[9]
port 114 nsew signal output
rlabel metal3 s 0 3680 800 3800 6 oram_addr[0]
port 115 nsew signal output
rlabel metal3 s 0 5856 800 5976 6 oram_addr[1]
port 116 nsew signal output
rlabel metal3 s 0 8032 800 8152 6 oram_addr[2]
port 117 nsew signal output
rlabel metal3 s 0 10208 800 10328 6 oram_addr[3]
port 118 nsew signal output
rlabel metal3 s 0 12384 800 12504 6 oram_addr[4]
port 119 nsew signal output
rlabel metal3 s 0 14560 800 14680 6 oram_addr[5]
port 120 nsew signal output
rlabel metal3 s 0 16736 800 16856 6 oram_addr[6]
port 121 nsew signal output
rlabel metal3 s 0 18912 800 19032 6 oram_addr[7]
port 122 nsew signal output
rlabel metal3 s 0 21088 800 21208 6 oram_addr[8]
port 123 nsew signal output
rlabel metal3 s 0 2592 800 2712 6 oram_csb
port 124 nsew signal output
rlabel metal3 s 0 4768 800 4888 6 oram_value[0]
port 125 nsew signal input
rlabel metal3 s 0 24352 800 24472 6 oram_value[10]
port 126 nsew signal input
rlabel metal3 s 0 25440 800 25560 6 oram_value[11]
port 127 nsew signal input
rlabel metal3 s 0 26528 800 26648 6 oram_value[12]
port 128 nsew signal input
rlabel metal3 s 0 27616 800 27736 6 oram_value[13]
port 129 nsew signal input
rlabel metal3 s 0 28704 800 28824 6 oram_value[14]
port 130 nsew signal input
rlabel metal3 s 0 29792 800 29912 6 oram_value[15]
port 131 nsew signal input
rlabel metal3 s 0 30880 800 31000 6 oram_value[16]
port 132 nsew signal input
rlabel metal3 s 0 31968 800 32088 6 oram_value[17]
port 133 nsew signal input
rlabel metal3 s 0 33056 800 33176 6 oram_value[18]
port 134 nsew signal input
rlabel metal3 s 0 34144 800 34264 6 oram_value[19]
port 135 nsew signal input
rlabel metal3 s 0 6944 800 7064 6 oram_value[1]
port 136 nsew signal input
rlabel metal3 s 0 35232 800 35352 6 oram_value[20]
port 137 nsew signal input
rlabel metal3 s 0 36320 800 36440 6 oram_value[21]
port 138 nsew signal input
rlabel metal3 s 0 37408 800 37528 6 oram_value[22]
port 139 nsew signal input
rlabel metal3 s 0 38496 800 38616 6 oram_value[23]
port 140 nsew signal input
rlabel metal3 s 0 39584 800 39704 6 oram_value[24]
port 141 nsew signal input
rlabel metal3 s 0 40672 800 40792 6 oram_value[25]
port 142 nsew signal input
rlabel metal3 s 0 41760 800 41880 6 oram_value[26]
port 143 nsew signal input
rlabel metal3 s 0 42848 800 42968 6 oram_value[27]
port 144 nsew signal input
rlabel metal3 s 0 43936 800 44056 6 oram_value[28]
port 145 nsew signal input
rlabel metal3 s 0 45024 800 45144 6 oram_value[29]
port 146 nsew signal input
rlabel metal3 s 0 9120 800 9240 6 oram_value[2]
port 147 nsew signal input
rlabel metal3 s 0 46112 800 46232 6 oram_value[30]
port 148 nsew signal input
rlabel metal3 s 0 47200 800 47320 6 oram_value[31]
port 149 nsew signal input
rlabel metal3 s 0 11296 800 11416 6 oram_value[3]
port 150 nsew signal input
rlabel metal3 s 0 13472 800 13592 6 oram_value[4]
port 151 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 oram_value[5]
port 152 nsew signal input
rlabel metal3 s 0 17824 800 17944 6 oram_value[6]
port 153 nsew signal input
rlabel metal3 s 0 20000 800 20120 6 oram_value[7]
port 154 nsew signal input
rlabel metal3 s 0 22176 800 22296 6 oram_value[8]
port 155 nsew signal input
rlabel metal3 s 0 23264 800 23384 6 oram_value[9]
port 156 nsew signal input
rlabel metal2 s 61290 0 61346 800 6 ram_adrb[0]
port 157 nsew signal output
rlabel metal2 s 64234 0 64290 800 6 ram_adrb[1]
port 158 nsew signal output
rlabel metal2 s 67178 0 67234 800 6 ram_adrb[2]
port 159 nsew signal output
rlabel metal2 s 70122 0 70178 800 6 ram_adrb[3]
port 160 nsew signal output
rlabel metal2 s 73066 0 73122 800 6 ram_adrb[4]
port 161 nsew signal output
rlabel metal2 s 74538 0 74594 800 6 ram_adrb[5]
port 162 nsew signal output
rlabel metal2 s 76010 0 76066 800 6 ram_adrb[6]
port 163 nsew signal output
rlabel metal2 s 77482 0 77538 800 6 ram_adrb[7]
port 164 nsew signal output
rlabel metal2 s 78954 0 79010 800 6 ram_adrb[8]
port 165 nsew signal output
rlabel metal2 s 58346 0 58402 800 6 ram_csb
port 166 nsew signal output
rlabel metal2 s 59818 0 59874 800 6 ram_web
port 167 nsew signal output
rlabel metal2 s 62762 0 62818 800 6 ram_wmask[0]
port 168 nsew signal output
rlabel metal2 s 65706 0 65762 800 6 ram_wmask[1]
port 169 nsew signal output
rlabel metal2 s 68650 0 68706 800 6 ram_wmask[2]
port 170 nsew signal output
rlabel metal2 s 71594 0 71650 800 6 ram_wmask[3]
port 171 nsew signal output
rlabel metal4 s 4208 2128 4528 47376 6 vccd1
port 172 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 47376 6 vccd1
port 172 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 47376 6 vccd1
port 172 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 47376 6 vssd1
port 173 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 47376 6 vssd1
port 173 nsew ground bidirectional
rlabel metal2 s 938 0 994 800 6 wb_clk_i
port 174 nsew signal input
rlabel metal2 s 2410 0 2466 800 6 wb_rst_i
port 175 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 wbs_ack_o
port 176 nsew signal output
rlabel metal2 s 11242 0 11298 800 6 wbs_adr_i[0]
port 177 nsew signal input
rlabel metal2 s 25962 0 26018 800 6 wbs_adr_i[10]
port 178 nsew signal input
rlabel metal2 s 27434 0 27490 800 6 wbs_adr_i[11]
port 179 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 wbs_adr_i[12]
port 180 nsew signal input
rlabel metal2 s 30378 0 30434 800 6 wbs_adr_i[13]
port 181 nsew signal input
rlabel metal2 s 31850 0 31906 800 6 wbs_adr_i[14]
port 182 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 wbs_adr_i[15]
port 183 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 wbs_adr_i[16]
port 184 nsew signal input
rlabel metal2 s 36266 0 36322 800 6 wbs_adr_i[17]
port 185 nsew signal input
rlabel metal2 s 37738 0 37794 800 6 wbs_adr_i[18]
port 186 nsew signal input
rlabel metal2 s 39210 0 39266 800 6 wbs_adr_i[19]
port 187 nsew signal input
rlabel metal2 s 12714 0 12770 800 6 wbs_adr_i[1]
port 188 nsew signal input
rlabel metal2 s 40682 0 40738 800 6 wbs_adr_i[20]
port 189 nsew signal input
rlabel metal2 s 42154 0 42210 800 6 wbs_adr_i[21]
port 190 nsew signal input
rlabel metal2 s 43626 0 43682 800 6 wbs_adr_i[22]
port 191 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 wbs_adr_i[23]
port 192 nsew signal input
rlabel metal2 s 46570 0 46626 800 6 wbs_adr_i[24]
port 193 nsew signal input
rlabel metal2 s 48042 0 48098 800 6 wbs_adr_i[25]
port 194 nsew signal input
rlabel metal2 s 49514 0 49570 800 6 wbs_adr_i[26]
port 195 nsew signal input
rlabel metal2 s 50986 0 51042 800 6 wbs_adr_i[27]
port 196 nsew signal input
rlabel metal2 s 52458 0 52514 800 6 wbs_adr_i[28]
port 197 nsew signal input
rlabel metal2 s 53930 0 53986 800 6 wbs_adr_i[29]
port 198 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 wbs_adr_i[2]
port 199 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 wbs_adr_i[30]
port 200 nsew signal input
rlabel metal2 s 56874 0 56930 800 6 wbs_adr_i[31]
port 201 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 wbs_adr_i[3]
port 202 nsew signal input
rlabel metal2 s 17130 0 17186 800 6 wbs_adr_i[4]
port 203 nsew signal input
rlabel metal2 s 18602 0 18658 800 6 wbs_adr_i[5]
port 204 nsew signal input
rlabel metal2 s 20074 0 20130 800 6 wbs_adr_i[6]
port 205 nsew signal input
rlabel metal2 s 21546 0 21602 800 6 wbs_adr_i[7]
port 206 nsew signal input
rlabel metal2 s 23018 0 23074 800 6 wbs_adr_i[8]
port 207 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 wbs_adr_i[9]
port 208 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 wbs_cyc_i
port 209 nsew signal input
rlabel metal2 s 6826 0 6882 800 6 wbs_dat_i
port 210 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 wbs_stb_i
port 211 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 wbs_we_i
port 212 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 80000 50000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 10410696
string GDS_FILE /home/optimal/mpw_builds/mpw-8-as1x00/openlane/wrapped_tms1x00/runs/22_12_20_09_23/results/signoff/wrapped_tms1x00.magic.gds
string GDS_START 573076
<< end >>

