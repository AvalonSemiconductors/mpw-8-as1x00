magic
tech sky130B
magscale 1 2
timestamp 1671191882
<< obsli1 >>
rect 1104 2159 158884 97393
<< obsm1 >>
rect 1104 2128 158884 97424
<< metal2 >>
rect 1950 99200 2006 100000
rect 3330 99200 3386 100000
rect 4710 99200 4766 100000
rect 6090 99200 6146 100000
rect 7470 99200 7526 100000
rect 8850 99200 8906 100000
rect 10230 99200 10286 100000
rect 11610 99200 11666 100000
rect 12990 99200 13046 100000
rect 14370 99200 14426 100000
rect 15750 99200 15806 100000
rect 17130 99200 17186 100000
rect 18510 99200 18566 100000
rect 19890 99200 19946 100000
rect 21270 99200 21326 100000
rect 22650 99200 22706 100000
rect 24030 99200 24086 100000
rect 25410 99200 25466 100000
rect 26790 99200 26846 100000
rect 28170 99200 28226 100000
rect 29550 99200 29606 100000
rect 30930 99200 30986 100000
rect 32310 99200 32366 100000
rect 33690 99200 33746 100000
rect 35070 99200 35126 100000
rect 36450 99200 36506 100000
rect 37830 99200 37886 100000
rect 39210 99200 39266 100000
rect 40590 99200 40646 100000
rect 41970 99200 42026 100000
rect 43350 99200 43406 100000
rect 44730 99200 44786 100000
rect 46110 99200 46166 100000
rect 47490 99200 47546 100000
rect 48870 99200 48926 100000
rect 50250 99200 50306 100000
rect 51630 99200 51686 100000
rect 53010 99200 53066 100000
rect 54390 99200 54446 100000
rect 55770 99200 55826 100000
rect 57150 99200 57206 100000
rect 58530 99200 58586 100000
rect 59910 99200 59966 100000
rect 61290 99200 61346 100000
rect 62670 99200 62726 100000
rect 64050 99200 64106 100000
rect 65430 99200 65486 100000
rect 66810 99200 66866 100000
rect 68190 99200 68246 100000
rect 69570 99200 69626 100000
rect 70950 99200 71006 100000
rect 72330 99200 72386 100000
rect 73710 99200 73766 100000
rect 75090 99200 75146 100000
rect 76470 99200 76526 100000
rect 77850 99200 77906 100000
rect 79230 99200 79286 100000
rect 80610 99200 80666 100000
rect 81990 99200 82046 100000
rect 83370 99200 83426 100000
rect 84750 99200 84806 100000
rect 86130 99200 86186 100000
rect 87510 99200 87566 100000
rect 88890 99200 88946 100000
rect 90270 99200 90326 100000
rect 91650 99200 91706 100000
rect 93030 99200 93086 100000
rect 94410 99200 94466 100000
rect 95790 99200 95846 100000
rect 97170 99200 97226 100000
rect 98550 99200 98606 100000
rect 99930 99200 99986 100000
rect 101310 99200 101366 100000
rect 102690 99200 102746 100000
rect 104070 99200 104126 100000
rect 105450 99200 105506 100000
rect 106830 99200 106886 100000
rect 108210 99200 108266 100000
rect 109590 99200 109646 100000
rect 110970 99200 111026 100000
rect 112350 99200 112406 100000
rect 113730 99200 113786 100000
rect 115110 99200 115166 100000
rect 116490 99200 116546 100000
rect 117870 99200 117926 100000
rect 119250 99200 119306 100000
rect 120630 99200 120686 100000
rect 122010 99200 122066 100000
rect 123390 99200 123446 100000
rect 124770 99200 124826 100000
rect 126150 99200 126206 100000
rect 127530 99200 127586 100000
rect 128910 99200 128966 100000
rect 130290 99200 130346 100000
rect 131670 99200 131726 100000
rect 133050 99200 133106 100000
rect 134430 99200 134486 100000
rect 135810 99200 135866 100000
rect 137190 99200 137246 100000
rect 138570 99200 138626 100000
rect 139950 99200 140006 100000
rect 141330 99200 141386 100000
rect 142710 99200 142766 100000
rect 144090 99200 144146 100000
rect 145470 99200 145526 100000
rect 146850 99200 146906 100000
rect 148230 99200 148286 100000
rect 149610 99200 149666 100000
rect 150990 99200 151046 100000
rect 152370 99200 152426 100000
rect 153750 99200 153806 100000
rect 155130 99200 155186 100000
rect 156510 99200 156566 100000
rect 157890 99200 157946 100000
rect 39946 0 40002 800
rect 119894 0 119950 800
<< obsm2 >>
rect 1582 99144 1894 99362
rect 2062 99144 3274 99362
rect 3442 99144 4654 99362
rect 4822 99144 6034 99362
rect 6202 99144 7414 99362
rect 7582 99144 8794 99362
rect 8962 99144 10174 99362
rect 10342 99144 11554 99362
rect 11722 99144 12934 99362
rect 13102 99144 14314 99362
rect 14482 99144 15694 99362
rect 15862 99144 17074 99362
rect 17242 99144 18454 99362
rect 18622 99144 19834 99362
rect 20002 99144 21214 99362
rect 21382 99144 22594 99362
rect 22762 99144 23974 99362
rect 24142 99144 25354 99362
rect 25522 99144 26734 99362
rect 26902 99144 28114 99362
rect 28282 99144 29494 99362
rect 29662 99144 30874 99362
rect 31042 99144 32254 99362
rect 32422 99144 33634 99362
rect 33802 99144 35014 99362
rect 35182 99144 36394 99362
rect 36562 99144 37774 99362
rect 37942 99144 39154 99362
rect 39322 99144 40534 99362
rect 40702 99144 41914 99362
rect 42082 99144 43294 99362
rect 43462 99144 44674 99362
rect 44842 99144 46054 99362
rect 46222 99144 47434 99362
rect 47602 99144 48814 99362
rect 48982 99144 50194 99362
rect 50362 99144 51574 99362
rect 51742 99144 52954 99362
rect 53122 99144 54334 99362
rect 54502 99144 55714 99362
rect 55882 99144 57094 99362
rect 57262 99144 58474 99362
rect 58642 99144 59854 99362
rect 60022 99144 61234 99362
rect 61402 99144 62614 99362
rect 62782 99144 63994 99362
rect 64162 99144 65374 99362
rect 65542 99144 66754 99362
rect 66922 99144 68134 99362
rect 68302 99144 69514 99362
rect 69682 99144 70894 99362
rect 71062 99144 72274 99362
rect 72442 99144 73654 99362
rect 73822 99144 75034 99362
rect 75202 99144 76414 99362
rect 76582 99144 77794 99362
rect 77962 99144 79174 99362
rect 79342 99144 80554 99362
rect 80722 99144 81934 99362
rect 82102 99144 83314 99362
rect 83482 99144 84694 99362
rect 84862 99144 86074 99362
rect 86242 99144 87454 99362
rect 87622 99144 88834 99362
rect 89002 99144 90214 99362
rect 90382 99144 91594 99362
rect 91762 99144 92974 99362
rect 93142 99144 94354 99362
rect 94522 99144 95734 99362
rect 95902 99144 97114 99362
rect 97282 99144 98494 99362
rect 98662 99144 99874 99362
rect 100042 99144 101254 99362
rect 101422 99144 102634 99362
rect 102802 99144 104014 99362
rect 104182 99144 105394 99362
rect 105562 99144 106774 99362
rect 106942 99144 108154 99362
rect 108322 99144 109534 99362
rect 109702 99144 110914 99362
rect 111082 99144 112294 99362
rect 112462 99144 113674 99362
rect 113842 99144 115054 99362
rect 115222 99144 116434 99362
rect 116602 99144 117814 99362
rect 117982 99144 119194 99362
rect 119362 99144 120574 99362
rect 120742 99144 121954 99362
rect 122122 99144 123334 99362
rect 123502 99144 124714 99362
rect 124882 99144 126094 99362
rect 126262 99144 127474 99362
rect 127642 99144 128854 99362
rect 129022 99144 130234 99362
rect 130402 99144 131614 99362
rect 131782 99144 132994 99362
rect 133162 99144 134374 99362
rect 134542 99144 135754 99362
rect 135922 99144 137134 99362
rect 137302 99144 138514 99362
rect 138682 99144 139894 99362
rect 140062 99144 141274 99362
rect 141442 99144 142654 99362
rect 142822 99144 144034 99362
rect 144202 99144 145414 99362
rect 145582 99144 146794 99362
rect 146962 99144 148174 99362
rect 148342 99144 149554 99362
rect 149722 99144 150934 99362
rect 151102 99144 152314 99362
rect 152482 99144 153694 99362
rect 153862 99144 155074 99362
rect 155242 99144 156454 99362
rect 156622 99144 157834 99362
rect 158002 99144 158122 99362
rect 1582 856 158122 99144
rect 1582 800 39890 856
rect 40058 800 119838 856
rect 120006 800 158122 856
<< metal3 >>
rect 0 96160 800 96280
rect 0 93848 800 93968
rect 0 91536 800 91656
rect 0 89224 800 89344
rect 0 86912 800 87032
rect 0 84600 800 84720
rect 0 82288 800 82408
rect 0 79976 800 80096
rect 0 77664 800 77784
rect 0 75352 800 75472
rect 0 73040 800 73160
rect 0 70728 800 70848
rect 0 68416 800 68536
rect 0 66104 800 66224
rect 0 63792 800 63912
rect 0 61480 800 61600
rect 0 59168 800 59288
rect 0 56856 800 56976
rect 0 54544 800 54664
rect 0 52232 800 52352
rect 0 49920 800 50040
rect 0 47608 800 47728
rect 0 45296 800 45416
rect 0 42984 800 43104
rect 0 40672 800 40792
rect 0 38360 800 38480
rect 0 36048 800 36168
rect 0 33736 800 33856
rect 0 31424 800 31544
rect 0 29112 800 29232
rect 0 26800 800 26920
rect 0 24488 800 24608
rect 0 22176 800 22296
rect 0 19864 800 19984
rect 0 17552 800 17672
rect 0 15240 800 15360
rect 0 12928 800 13048
rect 0 10616 800 10736
rect 0 8304 800 8424
rect 0 5992 800 6112
rect 0 3680 800 3800
<< obsm3 >>
rect 800 96360 158126 97409
rect 880 96080 158126 96360
rect 800 94048 158126 96080
rect 880 93768 158126 94048
rect 800 91736 158126 93768
rect 880 91456 158126 91736
rect 800 89424 158126 91456
rect 880 89144 158126 89424
rect 800 87112 158126 89144
rect 880 86832 158126 87112
rect 800 84800 158126 86832
rect 880 84520 158126 84800
rect 800 82488 158126 84520
rect 880 82208 158126 82488
rect 800 80176 158126 82208
rect 880 79896 158126 80176
rect 800 77864 158126 79896
rect 880 77584 158126 77864
rect 800 75552 158126 77584
rect 880 75272 158126 75552
rect 800 73240 158126 75272
rect 880 72960 158126 73240
rect 800 70928 158126 72960
rect 880 70648 158126 70928
rect 800 68616 158126 70648
rect 880 68336 158126 68616
rect 800 66304 158126 68336
rect 880 66024 158126 66304
rect 800 63992 158126 66024
rect 880 63712 158126 63992
rect 800 61680 158126 63712
rect 880 61400 158126 61680
rect 800 59368 158126 61400
rect 880 59088 158126 59368
rect 800 57056 158126 59088
rect 880 56776 158126 57056
rect 800 54744 158126 56776
rect 880 54464 158126 54744
rect 800 52432 158126 54464
rect 880 52152 158126 52432
rect 800 50120 158126 52152
rect 880 49840 158126 50120
rect 800 47808 158126 49840
rect 880 47528 158126 47808
rect 800 45496 158126 47528
rect 880 45216 158126 45496
rect 800 43184 158126 45216
rect 880 42904 158126 43184
rect 800 40872 158126 42904
rect 880 40592 158126 40872
rect 800 38560 158126 40592
rect 880 38280 158126 38560
rect 800 36248 158126 38280
rect 880 35968 158126 36248
rect 800 33936 158126 35968
rect 880 33656 158126 33936
rect 800 31624 158126 33656
rect 880 31344 158126 31624
rect 800 29312 158126 31344
rect 880 29032 158126 29312
rect 800 27000 158126 29032
rect 880 26720 158126 27000
rect 800 24688 158126 26720
rect 880 24408 158126 24688
rect 800 22376 158126 24408
rect 880 22096 158126 22376
rect 800 20064 158126 22096
rect 880 19784 158126 20064
rect 800 17752 158126 19784
rect 880 17472 158126 17752
rect 800 15440 158126 17472
rect 880 15160 158126 15440
rect 800 13128 158126 15160
rect 880 12848 158126 13128
rect 800 10816 158126 12848
rect 880 10536 158126 10816
rect 800 8504 158126 10536
rect 880 8224 158126 8504
rect 800 6192 158126 8224
rect 880 5912 158126 6192
rect 800 3880 158126 5912
rect 880 3600 158126 3880
rect 800 2143 158126 3600
<< metal4 >>
rect 4208 2128 4528 97424
rect 19568 2128 19888 97424
rect 34928 2128 35248 97424
rect 50288 2128 50608 97424
rect 65648 2128 65968 97424
rect 81008 2128 81328 97424
rect 96368 2128 96688 97424
rect 111728 2128 112048 97424
rect 127088 2128 127408 97424
rect 142448 2128 142768 97424
rect 157808 2128 158128 97424
<< obsm4 >>
rect 42931 5883 42997 9757
<< labels >>
rlabel metal2 s 1950 99200 2006 100000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 43350 99200 43406 100000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 47490 99200 47546 100000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 51630 99200 51686 100000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 55770 99200 55826 100000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 59910 99200 59966 100000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 64050 99200 64106 100000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 68190 99200 68246 100000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 72330 99200 72386 100000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 76470 99200 76526 100000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 80610 99200 80666 100000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 6090 99200 6146 100000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 84750 99200 84806 100000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 88890 99200 88946 100000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 93030 99200 93086 100000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 97170 99200 97226 100000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 101310 99200 101366 100000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 105450 99200 105506 100000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 109590 99200 109646 100000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 113730 99200 113786 100000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 117870 99200 117926 100000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 122010 99200 122066 100000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 10230 99200 10286 100000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 126150 99200 126206 100000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 130290 99200 130346 100000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 134430 99200 134486 100000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 138570 99200 138626 100000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 142710 99200 142766 100000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 146850 99200 146906 100000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 150990 99200 151046 100000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 155130 99200 155186 100000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 14370 99200 14426 100000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 18510 99200 18566 100000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 22650 99200 22706 100000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 26790 99200 26846 100000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 30930 99200 30986 100000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 35070 99200 35126 100000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 39210 99200 39266 100000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 3330 99200 3386 100000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 44730 99200 44786 100000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 48870 99200 48926 100000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 53010 99200 53066 100000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 57150 99200 57206 100000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 61290 99200 61346 100000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 65430 99200 65486 100000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 69570 99200 69626 100000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 73710 99200 73766 100000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 77850 99200 77906 100000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 81990 99200 82046 100000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 7470 99200 7526 100000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 86130 99200 86186 100000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 90270 99200 90326 100000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 94410 99200 94466 100000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 98550 99200 98606 100000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 102690 99200 102746 100000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 106830 99200 106886 100000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 110970 99200 111026 100000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 115110 99200 115166 100000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 119250 99200 119306 100000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 123390 99200 123446 100000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 11610 99200 11666 100000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 127530 99200 127586 100000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 131670 99200 131726 100000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 135810 99200 135866 100000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 139950 99200 140006 100000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 144090 99200 144146 100000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 148230 99200 148286 100000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 152370 99200 152426 100000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 156510 99200 156566 100000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 15750 99200 15806 100000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 19890 99200 19946 100000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 24030 99200 24086 100000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 28170 99200 28226 100000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 32310 99200 32366 100000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 36450 99200 36506 100000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 40590 99200 40646 100000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 4710 99200 4766 100000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 46110 99200 46166 100000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 50250 99200 50306 100000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 54390 99200 54446 100000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 58530 99200 58586 100000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 62670 99200 62726 100000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 66810 99200 66866 100000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 70950 99200 71006 100000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 75090 99200 75146 100000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 79230 99200 79286 100000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 83370 99200 83426 100000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 8850 99200 8906 100000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 87510 99200 87566 100000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 91650 99200 91706 100000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 95790 99200 95846 100000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 99930 99200 99986 100000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 104070 99200 104126 100000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 108210 99200 108266 100000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 112350 99200 112406 100000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 116490 99200 116546 100000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 120630 99200 120686 100000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 124770 99200 124826 100000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 12990 99200 13046 100000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 128910 99200 128966 100000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 133050 99200 133106 100000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 137190 99200 137246 100000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 141330 99200 141386 100000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 145470 99200 145526 100000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 149610 99200 149666 100000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 153750 99200 153806 100000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 157890 99200 157946 100000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 17130 99200 17186 100000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 21270 99200 21326 100000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 25410 99200 25466 100000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 29550 99200 29606 100000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 33690 99200 33746 100000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 37830 99200 37886 100000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 41970 99200 42026 100000 6 io_out[9]
port 114 nsew signal output
rlabel metal3 s 0 3680 800 3800 6 oram_addr[0]
port 115 nsew signal output
rlabel metal3 s 0 8304 800 8424 6 oram_addr[1]
port 116 nsew signal output
rlabel metal3 s 0 12928 800 13048 6 oram_addr[2]
port 117 nsew signal output
rlabel metal3 s 0 17552 800 17672 6 oram_addr[3]
port 118 nsew signal output
rlabel metal3 s 0 22176 800 22296 6 oram_addr[4]
port 119 nsew signal output
rlabel metal3 s 0 26800 800 26920 6 oram_addr[5]
port 120 nsew signal output
rlabel metal3 s 0 31424 800 31544 6 oram_addr[6]
port 121 nsew signal output
rlabel metal3 s 0 36048 800 36168 6 oram_addr[7]
port 122 nsew signal output
rlabel metal3 s 0 40672 800 40792 6 oram_addr[8]
port 123 nsew signal output
rlabel metal3 s 0 5992 800 6112 6 oram_value[0]
port 124 nsew signal input
rlabel metal3 s 0 47608 800 47728 6 oram_value[10]
port 125 nsew signal input
rlabel metal3 s 0 49920 800 50040 6 oram_value[11]
port 126 nsew signal input
rlabel metal3 s 0 52232 800 52352 6 oram_value[12]
port 127 nsew signal input
rlabel metal3 s 0 54544 800 54664 6 oram_value[13]
port 128 nsew signal input
rlabel metal3 s 0 56856 800 56976 6 oram_value[14]
port 129 nsew signal input
rlabel metal3 s 0 59168 800 59288 6 oram_value[15]
port 130 nsew signal input
rlabel metal3 s 0 61480 800 61600 6 oram_value[16]
port 131 nsew signal input
rlabel metal3 s 0 63792 800 63912 6 oram_value[17]
port 132 nsew signal input
rlabel metal3 s 0 66104 800 66224 6 oram_value[18]
port 133 nsew signal input
rlabel metal3 s 0 68416 800 68536 6 oram_value[19]
port 134 nsew signal input
rlabel metal3 s 0 10616 800 10736 6 oram_value[1]
port 135 nsew signal input
rlabel metal3 s 0 70728 800 70848 6 oram_value[20]
port 136 nsew signal input
rlabel metal3 s 0 73040 800 73160 6 oram_value[21]
port 137 nsew signal input
rlabel metal3 s 0 75352 800 75472 6 oram_value[22]
port 138 nsew signal input
rlabel metal3 s 0 77664 800 77784 6 oram_value[23]
port 139 nsew signal input
rlabel metal3 s 0 79976 800 80096 6 oram_value[24]
port 140 nsew signal input
rlabel metal3 s 0 82288 800 82408 6 oram_value[25]
port 141 nsew signal input
rlabel metal3 s 0 84600 800 84720 6 oram_value[26]
port 142 nsew signal input
rlabel metal3 s 0 86912 800 87032 6 oram_value[27]
port 143 nsew signal input
rlabel metal3 s 0 89224 800 89344 6 oram_value[28]
port 144 nsew signal input
rlabel metal3 s 0 91536 800 91656 6 oram_value[29]
port 145 nsew signal input
rlabel metal3 s 0 15240 800 15360 6 oram_value[2]
port 146 nsew signal input
rlabel metal3 s 0 93848 800 93968 6 oram_value[30]
port 147 nsew signal input
rlabel metal3 s 0 96160 800 96280 6 oram_value[31]
port 148 nsew signal input
rlabel metal3 s 0 19864 800 19984 6 oram_value[3]
port 149 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 oram_value[4]
port 150 nsew signal input
rlabel metal3 s 0 29112 800 29232 6 oram_value[5]
port 151 nsew signal input
rlabel metal3 s 0 33736 800 33856 6 oram_value[6]
port 152 nsew signal input
rlabel metal3 s 0 38360 800 38480 6 oram_value[7]
port 153 nsew signal input
rlabel metal3 s 0 42984 800 43104 6 oram_value[8]
port 154 nsew signal input
rlabel metal3 s 0 45296 800 45416 6 oram_value[9]
port 155 nsew signal input
rlabel metal4 s 4208 2128 4528 97424 6 vccd1
port 156 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 97424 6 vccd1
port 156 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 97424 6 vccd1
port 156 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 97424 6 vccd1
port 156 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 97424 6 vccd1
port 156 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 97424 6 vccd1
port 156 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 97424 6 vssd1
port 157 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 97424 6 vssd1
port 157 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 97424 6 vssd1
port 157 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 97424 6 vssd1
port 157 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 97424 6 vssd1
port 157 nsew ground bidirectional
rlabel metal2 s 39946 0 40002 800 6 wb_clk_i
port 158 nsew signal input
rlabel metal2 s 119894 0 119950 800 6 wb_rst_i
port 159 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 160000 100000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 4954566
string GDS_FILE /run/media/tholin/e6042058-84c8-448b-be8a-b40bc065b34b/caravel_user_project/openlane/wrapped_tms1x00/runs/22_12_16_12_52/results/signoff/wrapped_tms1x00.magic.gds
string GDS_START 287960
<< end >>

