VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_tms1x00
  CLASS BLOCK ;
  FOREIGN wrapped_tms1x00 ;
  ORIGIN 0.000 0.000 ;
  SIZE 650.000 BY 450.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 446.000 13.250 450.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.570 446.000 178.850 450.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.130 446.000 195.410 450.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.690 446.000 211.970 450.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.250 446.000 228.530 450.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 446.000 245.090 450.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.370 446.000 261.650 450.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.930 446.000 278.210 450.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.490 446.000 294.770 450.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.050 446.000 311.330 450.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.610 446.000 327.890 450.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 446.000 29.810 450.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.170 446.000 344.450 450.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 446.000 361.010 450.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.290 446.000 377.570 450.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.850 446.000 394.130 450.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.410 446.000 410.690 450.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.970 446.000 427.250 450.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.530 446.000 443.810 450.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.090 446.000 460.370 450.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.650 446.000 476.930 450.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.210 446.000 493.490 450.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 446.000 46.370 450.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.770 446.000 510.050 450.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.330 446.000 526.610 450.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.890 446.000 543.170 450.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.450 446.000 559.730 450.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.010 446.000 576.290 450.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.570 446.000 592.850 450.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.130 446.000 609.410 450.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 625.690 446.000 625.970 450.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 446.000 62.930 450.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 446.000 79.490 450.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 446.000 96.050 450.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 446.000 112.610 450.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 446.000 129.170 450.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.450 446.000 145.730 450.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 446.000 162.290 450.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 446.000 18.770 450.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 446.000 184.370 450.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.650 446.000 200.930 450.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.210 446.000 217.490 450.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 446.000 234.050 450.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.330 446.000 250.610 450.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 446.000 267.170 450.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 446.000 283.730 450.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.010 446.000 300.290 450.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.570 446.000 316.850 450.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.130 446.000 333.410 450.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 446.000 35.330 450.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.690 446.000 349.970 450.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.250 446.000 366.530 450.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.810 446.000 383.090 450.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 446.000 399.650 450.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.930 446.000 416.210 450.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.490 446.000 432.770 450.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.050 446.000 449.330 450.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.610 446.000 465.890 450.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.170 446.000 482.450 450.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.730 446.000 499.010 450.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 446.000 51.890 450.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.290 446.000 515.570 450.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.850 446.000 532.130 450.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 548.410 446.000 548.690 450.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.970 446.000 565.250 450.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.530 446.000 581.810 450.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.090 446.000 598.370 450.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.650 446.000 614.930 450.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.210 446.000 631.490 450.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 446.000 68.450 450.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 446.000 85.010 450.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 446.000 101.570 450.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 446.000 118.130 450.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.410 446.000 134.690 450.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 446.000 151.250 450.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 446.000 167.810 450.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 446.000 24.290 450.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.610 446.000 189.890 450.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 446.000 206.450 450.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.730 446.000 223.010 450.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.290 446.000 239.570 450.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.850 446.000 256.130 450.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.410 446.000 272.690 450.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.970 446.000 289.250 450.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.530 446.000 305.810 450.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 446.000 322.370 450.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.650 446.000 338.930 450.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 446.000 40.850 450.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.210 446.000 355.490 450.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.770 446.000 372.050 450.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.330 446.000 388.610 450.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.890 446.000 405.170 450.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.450 446.000 421.730 450.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 446.000 438.290 450.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.570 446.000 454.850 450.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.130 446.000 471.410 450.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.690 446.000 487.970 450.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.250 446.000 504.530 450.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 446.000 57.410 450.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.810 446.000 521.090 450.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.370 446.000 537.650 450.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 446.000 554.210 450.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.490 446.000 570.770 450.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.050 446.000 587.330 450.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.610 446.000 603.890 450.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.170 446.000 620.450 450.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 636.730 446.000 637.010 450.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 446.000 73.970 450.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 446.000 90.530 450.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 446.000 107.090 450.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 446.000 123.650 450.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.930 446.000 140.210 450.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.490 446.000 156.770 450.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.050 446.000 173.330 450.000 ;
    END
  END io_out[9]
  PIN ram_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 646.000 43.560 650.000 44.160 ;
    END
  END ram_addr[0]
  PIN ram_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 646.000 127.200 650.000 127.800 ;
    END
  END ram_addr[1]
  PIN ram_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 646.000 210.840 650.000 211.440 ;
    END
  END ram_addr[2]
  PIN ram_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 646.000 294.480 650.000 295.080 ;
    END
  END ram_addr[3]
  PIN ram_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 646.000 378.120 650.000 378.720 ;
    END
  END ram_addr[4]
  PIN ram_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 646.000 406.000 650.000 406.600 ;
    END
  END ram_addr[5]
  PIN ram_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 646.000 433.880 650.000 434.480 ;
    END
  END ram_addr[6]
  PIN ram_val_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 646.000 71.440 650.000 72.040 ;
    END
  END ram_val_in[0]
  PIN ram_val_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 646.000 155.080 650.000 155.680 ;
    END
  END ram_val_in[1]
  PIN ram_val_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 646.000 238.720 650.000 239.320 ;
    END
  END ram_val_in[2]
  PIN ram_val_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 646.000 322.360 650.000 322.960 ;
    END
  END ram_val_in[3]
  PIN ram_val_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 646.000 99.320 650.000 99.920 ;
    END
  END ram_val_out[0]
  PIN ram_val_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 646.000 182.960 650.000 183.560 ;
    END
  END ram_val_out[1]
  PIN ram_val_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 646.000 266.600 650.000 267.200 ;
    END
  END ram_val_out[2]
  PIN ram_val_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 646.000 350.240 650.000 350.840 ;
    END
  END ram_val_out[3]
  PIN ram_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 646.000 15.680 650.000 16.280 ;
    END
  END ram_we
  PIN rom_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END rom_addr[0]
  PIN rom_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END rom_addr[1]
  PIN rom_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 4.000 67.280 ;
    END
  END rom_addr[2]
  PIN rom_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END rom_addr[3]
  PIN rom_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 4.000 108.080 ;
    END
  END rom_addr[4]
  PIN rom_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END rom_addr[5]
  PIN rom_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 4.000 148.880 ;
    END
  END rom_addr[6]
  PIN rom_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 4.000 169.280 ;
    END
  END rom_addr[7]
  PIN rom_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 4.000 189.680 ;
    END
  END rom_addr[8]
  PIN rom_csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.680 4.000 16.280 ;
    END
  END rom_csb
  PIN rom_value[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.080 4.000 36.680 ;
    END
  END rom_value[0]
  PIN rom_value[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.680 4.000 220.280 ;
    END
  END rom_value[10]
  PIN rom_value[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.880 4.000 230.480 ;
    END
  END rom_value[11]
  PIN rom_value[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.080 4.000 240.680 ;
    END
  END rom_value[12]
  PIN rom_value[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.280 4.000 250.880 ;
    END
  END rom_value[13]
  PIN rom_value[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 260.480 4.000 261.080 ;
    END
  END rom_value[14]
  PIN rom_value[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.680 4.000 271.280 ;
    END
  END rom_value[15]
  PIN rom_value[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.880 4.000 281.480 ;
    END
  END rom_value[16]
  PIN rom_value[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.080 4.000 291.680 ;
    END
  END rom_value[17]
  PIN rom_value[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.280 4.000 301.880 ;
    END
  END rom_value[18]
  PIN rom_value[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 311.480 4.000 312.080 ;
    END
  END rom_value[19]
  PIN rom_value[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.480 4.000 57.080 ;
    END
  END rom_value[1]
  PIN rom_value[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.680 4.000 322.280 ;
    END
  END rom_value[20]
  PIN rom_value[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.880 4.000 332.480 ;
    END
  END rom_value[21]
  PIN rom_value[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.080 4.000 342.680 ;
    END
  END rom_value[22]
  PIN rom_value[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.280 4.000 352.880 ;
    END
  END rom_value[23]
  PIN rom_value[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 362.480 4.000 363.080 ;
    END
  END rom_value[24]
  PIN rom_value[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 372.680 4.000 373.280 ;
    END
  END rom_value[25]
  PIN rom_value[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 382.880 4.000 383.480 ;
    END
  END rom_value[26]
  PIN rom_value[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.080 4.000 393.680 ;
    END
  END rom_value[27]
  PIN rom_value[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 403.280 4.000 403.880 ;
    END
  END rom_value[28]
  PIN rom_value[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 413.480 4.000 414.080 ;
    END
  END rom_value[29]
  PIN rom_value[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.880 4.000 77.480 ;
    END
  END rom_value[2]
  PIN rom_value[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 423.680 4.000 424.280 ;
    END
  END rom_value[30]
  PIN rom_value[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 433.880 4.000 434.480 ;
    END
  END rom_value[31]
  PIN rom_value[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.280 4.000 97.880 ;
    END
  END rom_value[3]
  PIN rom_value[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.680 4.000 118.280 ;
    END
  END rom_value[4]
  PIN rom_value[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.080 4.000 138.680 ;
    END
  END rom_value[5]
  PIN rom_value[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 158.480 4.000 159.080 ;
    END
  END rom_value[6]
  PIN rom_value[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.880 4.000 179.480 ;
    END
  END rom_value[7]
  PIN rom_value[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.280 4.000 199.880 ;
    END
  END rom_value[8]
  PIN rom_value[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END rom_value[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 438.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 438.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 438.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 438.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 438.160 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 438.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 438.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 438.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 438.160 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 4.000 ;
    END
  END wb_clk_i
  PIN wb_rom_adrb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 4.000 ;
    END
  END wb_rom_adrb[0]
  PIN wb_rom_adrb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END wb_rom_adrb[1]
  PIN wb_rom_adrb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 4.000 ;
    END
  END wb_rom_adrb[2]
  PIN wb_rom_adrb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 4.000 ;
    END
  END wb_rom_adrb[3]
  PIN wb_rom_adrb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 0.000 76.730 4.000 ;
    END
  END wb_rom_adrb[4]
  PIN wb_rom_adrb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 0.000 85.010 4.000 ;
    END
  END wb_rom_adrb[5]
  PIN wb_rom_adrb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 4.000 ;
    END
  END wb_rom_adrb[6]
  PIN wb_rom_adrb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 0.000 101.570 4.000 ;
    END
  END wb_rom_adrb[7]
  PIN wb_rom_adrb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END wb_rom_adrb[8]
  PIN wb_rom_csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 0.000 31.190 4.000 ;
    END
  END wb_rom_csb
  PIN wb_rom_val[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 0.000 47.750 4.000 ;
    END
  END wb_rom_val[0]
  PIN wb_rom_val[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 0.000 122.270 4.000 ;
    END
  END wb_rom_val[10]
  PIN wb_rom_val[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 0.000 126.410 4.000 ;
    END
  END wb_rom_val[11]
  PIN wb_rom_val[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.270 0.000 130.550 4.000 ;
    END
  END wb_rom_val[12]
  PIN wb_rom_val[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.410 0.000 134.690 4.000 ;
    END
  END wb_rom_val[13]
  PIN wb_rom_val[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END wb_rom_val[14]
  PIN wb_rom_val[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END wb_rom_val[15]
  PIN wb_rom_val[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 0.000 147.110 4.000 ;
    END
  END wb_rom_val[16]
  PIN wb_rom_val[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 0.000 151.250 4.000 ;
    END
  END wb_rom_val[17]
  PIN wb_rom_val[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 0.000 155.390 4.000 ;
    END
  END wb_rom_val[18]
  PIN wb_rom_val[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.250 0.000 159.530 4.000 ;
    END
  END wb_rom_val[19]
  PIN wb_rom_val[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 4.000 ;
    END
  END wb_rom_val[1]
  PIN wb_rom_val[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 0.000 163.670 4.000 ;
    END
  END wb_rom_val[20]
  PIN wb_rom_val[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END wb_rom_val[21]
  PIN wb_rom_val[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.670 0.000 171.950 4.000 ;
    END
  END wb_rom_val[22]
  PIN wb_rom_val[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.810 0.000 176.090 4.000 ;
    END
  END wb_rom_val[23]
  PIN wb_rom_val[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.950 0.000 180.230 4.000 ;
    END
  END wb_rom_val[24]
  PIN wb_rom_val[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 0.000 184.370 4.000 ;
    END
  END wb_rom_val[25]
  PIN wb_rom_val[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.230 0.000 188.510 4.000 ;
    END
  END wb_rom_val[26]
  PIN wb_rom_val[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 0.000 192.650 4.000 ;
    END
  END wb_rom_val[27]
  PIN wb_rom_val[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 0.000 196.790 4.000 ;
    END
  END wb_rom_val[28]
  PIN wb_rom_val[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.650 0.000 200.930 4.000 ;
    END
  END wb_rom_val[29]
  PIN wb_rom_val[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 0.000 64.310 4.000 ;
    END
  END wb_rom_val[2]
  PIN wb_rom_val[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.790 0.000 205.070 4.000 ;
    END
  END wb_rom_val[30]
  PIN wb_rom_val[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.930 0.000 209.210 4.000 ;
    END
  END wb_rom_val[31]
  PIN wb_rom_val[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 4.000 ;
    END
  END wb_rom_val[3]
  PIN wb_rom_val[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END wb_rom_val[4]
  PIN wb_rom_val[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 0.000 89.150 4.000 ;
    END
  END wb_rom_val[5]
  PIN wb_rom_val[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.150 0.000 97.430 4.000 ;
    END
  END wb_rom_val[6]
  PIN wb_rom_val[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 0.000 105.710 4.000 ;
    END
  END wb_rom_val[7]
  PIN wb_rom_val[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.710 0.000 113.990 4.000 ;
    END
  END wb_rom_val[8]
  PIN wb_rom_val[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 0.000 118.130 4.000 ;
    END
  END wb_rom_val[9]
  PIN wb_rom_web
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 4.000 ;
    END
  END wb_rom_web
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 0.000 39.470 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.070 0.000 213.350 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 0.000 229.910 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.830 0.000 354.110 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.250 0.000 366.530 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.670 0.000 378.950 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.090 0.000 391.370 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.510 0.000 403.790 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.930 0.000 416.210 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 0.000 428.630 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.770 0.000 441.050 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.190 0.000 453.470 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.610 0.000 465.890 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.050 0.000 242.330 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.030 0.000 478.310 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.450 0.000 490.730 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.870 0.000 503.150 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.290 0.000 515.570 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.710 0.000 527.990 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.130 0.000 540.410 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.550 0.000 552.830 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.970 0.000 565.250 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.390 0.000 577.670 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.810 0.000 590.090 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 0.000 254.750 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.230 0.000 602.510 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.650 0.000 614.930 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 0.000 267.170 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.310 0.000 279.590 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.730 0.000 292.010 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.150 0.000 304.430 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.570 0.000 316.850 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.990 0.000 329.270 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 0.000 341.690 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.210 0.000 217.490 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 0.000 234.050 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.970 0.000 358.250 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.810 0.000 383.090 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.230 0.000 395.510 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.650 0.000 407.930 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.070 0.000 420.350 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.490 0.000 432.770 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.910 0.000 445.190 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 0.000 457.610 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.750 0.000 470.030 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.190 0.000 246.470 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.170 0.000 482.450 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 494.590 0.000 494.870 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.010 0.000 507.290 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.430 0.000 519.710 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.850 0.000 532.130 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 0.000 544.550 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.690 0.000 556.970 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.110 0.000 569.390 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.530 0.000 581.810 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.950 0.000 594.230 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 0.000 258.890 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.370 0.000 606.650 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.790 0.000 619.070 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.030 0.000 271.310 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.870 0.000 296.150 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.290 0.000 308.570 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.710 0.000 320.990 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.130 0.000 333.410 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.550 0.000 345.830 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.910 0.000 238.190 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.110 0.000 362.390 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.530 0.000 374.810 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.950 0.000 387.230 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 0.000 399.650 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.790 0.000 412.070 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.210 0.000 424.490 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.630 0.000 436.910 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.050 0.000 449.330 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.470 0.000 461.750 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.890 0.000 474.170 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.330 0.000 250.610 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.310 0.000 486.590 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.730 0.000 499.010 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.150 0.000 511.430 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.570 0.000 523.850 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.990 0.000 536.270 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 548.410 0.000 548.690 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.830 0.000 561.110 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 0.000 573.530 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.670 0.000 585.950 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.090 0.000 598.370 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.750 0.000 263.030 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.510 0.000 610.790 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.930 0.000 623.210 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.170 0.000 275.450 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.590 0.000 287.870 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.010 0.000 300.290 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 0.000 312.710 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.850 0.000 325.130 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.270 0.000 337.550 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.690 0.000 349.970 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.350 0.000 221.630 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 644.460 438.005 ;
      LAYER met1 ;
        RECT 4.670 2.420 645.310 438.160 ;
      LAYER met2 ;
        RECT 4.690 445.720 12.690 446.490 ;
        RECT 13.530 445.720 18.210 446.490 ;
        RECT 19.050 445.720 23.730 446.490 ;
        RECT 24.570 445.720 29.250 446.490 ;
        RECT 30.090 445.720 34.770 446.490 ;
        RECT 35.610 445.720 40.290 446.490 ;
        RECT 41.130 445.720 45.810 446.490 ;
        RECT 46.650 445.720 51.330 446.490 ;
        RECT 52.170 445.720 56.850 446.490 ;
        RECT 57.690 445.720 62.370 446.490 ;
        RECT 63.210 445.720 67.890 446.490 ;
        RECT 68.730 445.720 73.410 446.490 ;
        RECT 74.250 445.720 78.930 446.490 ;
        RECT 79.770 445.720 84.450 446.490 ;
        RECT 85.290 445.720 89.970 446.490 ;
        RECT 90.810 445.720 95.490 446.490 ;
        RECT 96.330 445.720 101.010 446.490 ;
        RECT 101.850 445.720 106.530 446.490 ;
        RECT 107.370 445.720 112.050 446.490 ;
        RECT 112.890 445.720 117.570 446.490 ;
        RECT 118.410 445.720 123.090 446.490 ;
        RECT 123.930 445.720 128.610 446.490 ;
        RECT 129.450 445.720 134.130 446.490 ;
        RECT 134.970 445.720 139.650 446.490 ;
        RECT 140.490 445.720 145.170 446.490 ;
        RECT 146.010 445.720 150.690 446.490 ;
        RECT 151.530 445.720 156.210 446.490 ;
        RECT 157.050 445.720 161.730 446.490 ;
        RECT 162.570 445.720 167.250 446.490 ;
        RECT 168.090 445.720 172.770 446.490 ;
        RECT 173.610 445.720 178.290 446.490 ;
        RECT 179.130 445.720 183.810 446.490 ;
        RECT 184.650 445.720 189.330 446.490 ;
        RECT 190.170 445.720 194.850 446.490 ;
        RECT 195.690 445.720 200.370 446.490 ;
        RECT 201.210 445.720 205.890 446.490 ;
        RECT 206.730 445.720 211.410 446.490 ;
        RECT 212.250 445.720 216.930 446.490 ;
        RECT 217.770 445.720 222.450 446.490 ;
        RECT 223.290 445.720 227.970 446.490 ;
        RECT 228.810 445.720 233.490 446.490 ;
        RECT 234.330 445.720 239.010 446.490 ;
        RECT 239.850 445.720 244.530 446.490 ;
        RECT 245.370 445.720 250.050 446.490 ;
        RECT 250.890 445.720 255.570 446.490 ;
        RECT 256.410 445.720 261.090 446.490 ;
        RECT 261.930 445.720 266.610 446.490 ;
        RECT 267.450 445.720 272.130 446.490 ;
        RECT 272.970 445.720 277.650 446.490 ;
        RECT 278.490 445.720 283.170 446.490 ;
        RECT 284.010 445.720 288.690 446.490 ;
        RECT 289.530 445.720 294.210 446.490 ;
        RECT 295.050 445.720 299.730 446.490 ;
        RECT 300.570 445.720 305.250 446.490 ;
        RECT 306.090 445.720 310.770 446.490 ;
        RECT 311.610 445.720 316.290 446.490 ;
        RECT 317.130 445.720 321.810 446.490 ;
        RECT 322.650 445.720 327.330 446.490 ;
        RECT 328.170 445.720 332.850 446.490 ;
        RECT 333.690 445.720 338.370 446.490 ;
        RECT 339.210 445.720 343.890 446.490 ;
        RECT 344.730 445.720 349.410 446.490 ;
        RECT 350.250 445.720 354.930 446.490 ;
        RECT 355.770 445.720 360.450 446.490 ;
        RECT 361.290 445.720 365.970 446.490 ;
        RECT 366.810 445.720 371.490 446.490 ;
        RECT 372.330 445.720 377.010 446.490 ;
        RECT 377.850 445.720 382.530 446.490 ;
        RECT 383.370 445.720 388.050 446.490 ;
        RECT 388.890 445.720 393.570 446.490 ;
        RECT 394.410 445.720 399.090 446.490 ;
        RECT 399.930 445.720 404.610 446.490 ;
        RECT 405.450 445.720 410.130 446.490 ;
        RECT 410.970 445.720 415.650 446.490 ;
        RECT 416.490 445.720 421.170 446.490 ;
        RECT 422.010 445.720 426.690 446.490 ;
        RECT 427.530 445.720 432.210 446.490 ;
        RECT 433.050 445.720 437.730 446.490 ;
        RECT 438.570 445.720 443.250 446.490 ;
        RECT 444.090 445.720 448.770 446.490 ;
        RECT 449.610 445.720 454.290 446.490 ;
        RECT 455.130 445.720 459.810 446.490 ;
        RECT 460.650 445.720 465.330 446.490 ;
        RECT 466.170 445.720 470.850 446.490 ;
        RECT 471.690 445.720 476.370 446.490 ;
        RECT 477.210 445.720 481.890 446.490 ;
        RECT 482.730 445.720 487.410 446.490 ;
        RECT 488.250 445.720 492.930 446.490 ;
        RECT 493.770 445.720 498.450 446.490 ;
        RECT 499.290 445.720 503.970 446.490 ;
        RECT 504.810 445.720 509.490 446.490 ;
        RECT 510.330 445.720 515.010 446.490 ;
        RECT 515.850 445.720 520.530 446.490 ;
        RECT 521.370 445.720 526.050 446.490 ;
        RECT 526.890 445.720 531.570 446.490 ;
        RECT 532.410 445.720 537.090 446.490 ;
        RECT 537.930 445.720 542.610 446.490 ;
        RECT 543.450 445.720 548.130 446.490 ;
        RECT 548.970 445.720 553.650 446.490 ;
        RECT 554.490 445.720 559.170 446.490 ;
        RECT 560.010 445.720 564.690 446.490 ;
        RECT 565.530 445.720 570.210 446.490 ;
        RECT 571.050 445.720 575.730 446.490 ;
        RECT 576.570 445.720 581.250 446.490 ;
        RECT 582.090 445.720 586.770 446.490 ;
        RECT 587.610 445.720 592.290 446.490 ;
        RECT 593.130 445.720 597.810 446.490 ;
        RECT 598.650 445.720 603.330 446.490 ;
        RECT 604.170 445.720 608.850 446.490 ;
        RECT 609.690 445.720 614.370 446.490 ;
        RECT 615.210 445.720 619.890 446.490 ;
        RECT 620.730 445.720 625.410 446.490 ;
        RECT 626.250 445.720 630.930 446.490 ;
        RECT 631.770 445.720 636.450 446.490 ;
        RECT 637.290 445.720 645.290 446.490 ;
        RECT 4.690 4.280 645.290 445.720 ;
        RECT 4.690 2.390 26.490 4.280 ;
        RECT 27.330 2.390 30.630 4.280 ;
        RECT 31.470 2.390 34.770 4.280 ;
        RECT 35.610 2.390 38.910 4.280 ;
        RECT 39.750 2.390 43.050 4.280 ;
        RECT 43.890 2.390 47.190 4.280 ;
        RECT 48.030 2.390 51.330 4.280 ;
        RECT 52.170 2.390 55.470 4.280 ;
        RECT 56.310 2.390 59.610 4.280 ;
        RECT 60.450 2.390 63.750 4.280 ;
        RECT 64.590 2.390 67.890 4.280 ;
        RECT 68.730 2.390 72.030 4.280 ;
        RECT 72.870 2.390 76.170 4.280 ;
        RECT 77.010 2.390 80.310 4.280 ;
        RECT 81.150 2.390 84.450 4.280 ;
        RECT 85.290 2.390 88.590 4.280 ;
        RECT 89.430 2.390 92.730 4.280 ;
        RECT 93.570 2.390 96.870 4.280 ;
        RECT 97.710 2.390 101.010 4.280 ;
        RECT 101.850 2.390 105.150 4.280 ;
        RECT 105.990 2.390 109.290 4.280 ;
        RECT 110.130 2.390 113.430 4.280 ;
        RECT 114.270 2.390 117.570 4.280 ;
        RECT 118.410 2.390 121.710 4.280 ;
        RECT 122.550 2.390 125.850 4.280 ;
        RECT 126.690 2.390 129.990 4.280 ;
        RECT 130.830 2.390 134.130 4.280 ;
        RECT 134.970 2.390 138.270 4.280 ;
        RECT 139.110 2.390 142.410 4.280 ;
        RECT 143.250 2.390 146.550 4.280 ;
        RECT 147.390 2.390 150.690 4.280 ;
        RECT 151.530 2.390 154.830 4.280 ;
        RECT 155.670 2.390 158.970 4.280 ;
        RECT 159.810 2.390 163.110 4.280 ;
        RECT 163.950 2.390 167.250 4.280 ;
        RECT 168.090 2.390 171.390 4.280 ;
        RECT 172.230 2.390 175.530 4.280 ;
        RECT 176.370 2.390 179.670 4.280 ;
        RECT 180.510 2.390 183.810 4.280 ;
        RECT 184.650 2.390 187.950 4.280 ;
        RECT 188.790 2.390 192.090 4.280 ;
        RECT 192.930 2.390 196.230 4.280 ;
        RECT 197.070 2.390 200.370 4.280 ;
        RECT 201.210 2.390 204.510 4.280 ;
        RECT 205.350 2.390 208.650 4.280 ;
        RECT 209.490 2.390 212.790 4.280 ;
        RECT 213.630 2.390 216.930 4.280 ;
        RECT 217.770 2.390 221.070 4.280 ;
        RECT 221.910 2.390 225.210 4.280 ;
        RECT 226.050 2.390 229.350 4.280 ;
        RECT 230.190 2.390 233.490 4.280 ;
        RECT 234.330 2.390 237.630 4.280 ;
        RECT 238.470 2.390 241.770 4.280 ;
        RECT 242.610 2.390 245.910 4.280 ;
        RECT 246.750 2.390 250.050 4.280 ;
        RECT 250.890 2.390 254.190 4.280 ;
        RECT 255.030 2.390 258.330 4.280 ;
        RECT 259.170 2.390 262.470 4.280 ;
        RECT 263.310 2.390 266.610 4.280 ;
        RECT 267.450 2.390 270.750 4.280 ;
        RECT 271.590 2.390 274.890 4.280 ;
        RECT 275.730 2.390 279.030 4.280 ;
        RECT 279.870 2.390 283.170 4.280 ;
        RECT 284.010 2.390 287.310 4.280 ;
        RECT 288.150 2.390 291.450 4.280 ;
        RECT 292.290 2.390 295.590 4.280 ;
        RECT 296.430 2.390 299.730 4.280 ;
        RECT 300.570 2.390 303.870 4.280 ;
        RECT 304.710 2.390 308.010 4.280 ;
        RECT 308.850 2.390 312.150 4.280 ;
        RECT 312.990 2.390 316.290 4.280 ;
        RECT 317.130 2.390 320.430 4.280 ;
        RECT 321.270 2.390 324.570 4.280 ;
        RECT 325.410 2.390 328.710 4.280 ;
        RECT 329.550 2.390 332.850 4.280 ;
        RECT 333.690 2.390 336.990 4.280 ;
        RECT 337.830 2.390 341.130 4.280 ;
        RECT 341.970 2.390 345.270 4.280 ;
        RECT 346.110 2.390 349.410 4.280 ;
        RECT 350.250 2.390 353.550 4.280 ;
        RECT 354.390 2.390 357.690 4.280 ;
        RECT 358.530 2.390 361.830 4.280 ;
        RECT 362.670 2.390 365.970 4.280 ;
        RECT 366.810 2.390 370.110 4.280 ;
        RECT 370.950 2.390 374.250 4.280 ;
        RECT 375.090 2.390 378.390 4.280 ;
        RECT 379.230 2.390 382.530 4.280 ;
        RECT 383.370 2.390 386.670 4.280 ;
        RECT 387.510 2.390 390.810 4.280 ;
        RECT 391.650 2.390 394.950 4.280 ;
        RECT 395.790 2.390 399.090 4.280 ;
        RECT 399.930 2.390 403.230 4.280 ;
        RECT 404.070 2.390 407.370 4.280 ;
        RECT 408.210 2.390 411.510 4.280 ;
        RECT 412.350 2.390 415.650 4.280 ;
        RECT 416.490 2.390 419.790 4.280 ;
        RECT 420.630 2.390 423.930 4.280 ;
        RECT 424.770 2.390 428.070 4.280 ;
        RECT 428.910 2.390 432.210 4.280 ;
        RECT 433.050 2.390 436.350 4.280 ;
        RECT 437.190 2.390 440.490 4.280 ;
        RECT 441.330 2.390 444.630 4.280 ;
        RECT 445.470 2.390 448.770 4.280 ;
        RECT 449.610 2.390 452.910 4.280 ;
        RECT 453.750 2.390 457.050 4.280 ;
        RECT 457.890 2.390 461.190 4.280 ;
        RECT 462.030 2.390 465.330 4.280 ;
        RECT 466.170 2.390 469.470 4.280 ;
        RECT 470.310 2.390 473.610 4.280 ;
        RECT 474.450 2.390 477.750 4.280 ;
        RECT 478.590 2.390 481.890 4.280 ;
        RECT 482.730 2.390 486.030 4.280 ;
        RECT 486.870 2.390 490.170 4.280 ;
        RECT 491.010 2.390 494.310 4.280 ;
        RECT 495.150 2.390 498.450 4.280 ;
        RECT 499.290 2.390 502.590 4.280 ;
        RECT 503.430 2.390 506.730 4.280 ;
        RECT 507.570 2.390 510.870 4.280 ;
        RECT 511.710 2.390 515.010 4.280 ;
        RECT 515.850 2.390 519.150 4.280 ;
        RECT 519.990 2.390 523.290 4.280 ;
        RECT 524.130 2.390 527.430 4.280 ;
        RECT 528.270 2.390 531.570 4.280 ;
        RECT 532.410 2.390 535.710 4.280 ;
        RECT 536.550 2.390 539.850 4.280 ;
        RECT 540.690 2.390 543.990 4.280 ;
        RECT 544.830 2.390 548.130 4.280 ;
        RECT 548.970 2.390 552.270 4.280 ;
        RECT 553.110 2.390 556.410 4.280 ;
        RECT 557.250 2.390 560.550 4.280 ;
        RECT 561.390 2.390 564.690 4.280 ;
        RECT 565.530 2.390 568.830 4.280 ;
        RECT 569.670 2.390 572.970 4.280 ;
        RECT 573.810 2.390 577.110 4.280 ;
        RECT 577.950 2.390 581.250 4.280 ;
        RECT 582.090 2.390 585.390 4.280 ;
        RECT 586.230 2.390 589.530 4.280 ;
        RECT 590.370 2.390 593.670 4.280 ;
        RECT 594.510 2.390 597.810 4.280 ;
        RECT 598.650 2.390 601.950 4.280 ;
        RECT 602.790 2.390 606.090 4.280 ;
        RECT 606.930 2.390 610.230 4.280 ;
        RECT 611.070 2.390 614.370 4.280 ;
        RECT 615.210 2.390 618.510 4.280 ;
        RECT 619.350 2.390 622.650 4.280 ;
        RECT 623.490 2.390 645.290 4.280 ;
      LAYER met3 ;
        RECT 4.000 434.880 646.000 438.085 ;
        RECT 4.400 433.480 645.600 434.880 ;
        RECT 4.000 424.680 646.000 433.480 ;
        RECT 4.400 423.280 646.000 424.680 ;
        RECT 4.000 414.480 646.000 423.280 ;
        RECT 4.400 413.080 646.000 414.480 ;
        RECT 4.000 407.000 646.000 413.080 ;
        RECT 4.000 405.600 645.600 407.000 ;
        RECT 4.000 404.280 646.000 405.600 ;
        RECT 4.400 402.880 646.000 404.280 ;
        RECT 4.000 394.080 646.000 402.880 ;
        RECT 4.400 392.680 646.000 394.080 ;
        RECT 4.000 383.880 646.000 392.680 ;
        RECT 4.400 382.480 646.000 383.880 ;
        RECT 4.000 379.120 646.000 382.480 ;
        RECT 4.000 377.720 645.600 379.120 ;
        RECT 4.000 373.680 646.000 377.720 ;
        RECT 4.400 372.280 646.000 373.680 ;
        RECT 4.000 363.480 646.000 372.280 ;
        RECT 4.400 362.080 646.000 363.480 ;
        RECT 4.000 353.280 646.000 362.080 ;
        RECT 4.400 351.880 646.000 353.280 ;
        RECT 4.000 351.240 646.000 351.880 ;
        RECT 4.000 349.840 645.600 351.240 ;
        RECT 4.000 343.080 646.000 349.840 ;
        RECT 4.400 341.680 646.000 343.080 ;
        RECT 4.000 332.880 646.000 341.680 ;
        RECT 4.400 331.480 646.000 332.880 ;
        RECT 4.000 323.360 646.000 331.480 ;
        RECT 4.000 322.680 645.600 323.360 ;
        RECT 4.400 321.960 645.600 322.680 ;
        RECT 4.400 321.280 646.000 321.960 ;
        RECT 4.000 312.480 646.000 321.280 ;
        RECT 4.400 311.080 646.000 312.480 ;
        RECT 4.000 302.280 646.000 311.080 ;
        RECT 4.400 300.880 646.000 302.280 ;
        RECT 4.000 295.480 646.000 300.880 ;
        RECT 4.000 294.080 645.600 295.480 ;
        RECT 4.000 292.080 646.000 294.080 ;
        RECT 4.400 290.680 646.000 292.080 ;
        RECT 4.000 281.880 646.000 290.680 ;
        RECT 4.400 280.480 646.000 281.880 ;
        RECT 4.000 271.680 646.000 280.480 ;
        RECT 4.400 270.280 646.000 271.680 ;
        RECT 4.000 267.600 646.000 270.280 ;
        RECT 4.000 266.200 645.600 267.600 ;
        RECT 4.000 261.480 646.000 266.200 ;
        RECT 4.400 260.080 646.000 261.480 ;
        RECT 4.000 251.280 646.000 260.080 ;
        RECT 4.400 249.880 646.000 251.280 ;
        RECT 4.000 241.080 646.000 249.880 ;
        RECT 4.400 239.720 646.000 241.080 ;
        RECT 4.400 239.680 645.600 239.720 ;
        RECT 4.000 238.320 645.600 239.680 ;
        RECT 4.000 230.880 646.000 238.320 ;
        RECT 4.400 229.480 646.000 230.880 ;
        RECT 4.000 220.680 646.000 229.480 ;
        RECT 4.400 219.280 646.000 220.680 ;
        RECT 4.000 211.840 646.000 219.280 ;
        RECT 4.000 210.480 645.600 211.840 ;
        RECT 4.400 210.440 645.600 210.480 ;
        RECT 4.400 209.080 646.000 210.440 ;
        RECT 4.000 200.280 646.000 209.080 ;
        RECT 4.400 198.880 646.000 200.280 ;
        RECT 4.000 190.080 646.000 198.880 ;
        RECT 4.400 188.680 646.000 190.080 ;
        RECT 4.000 183.960 646.000 188.680 ;
        RECT 4.000 182.560 645.600 183.960 ;
        RECT 4.000 179.880 646.000 182.560 ;
        RECT 4.400 178.480 646.000 179.880 ;
        RECT 4.000 169.680 646.000 178.480 ;
        RECT 4.400 168.280 646.000 169.680 ;
        RECT 4.000 159.480 646.000 168.280 ;
        RECT 4.400 158.080 646.000 159.480 ;
        RECT 4.000 156.080 646.000 158.080 ;
        RECT 4.000 154.680 645.600 156.080 ;
        RECT 4.000 149.280 646.000 154.680 ;
        RECT 4.400 147.880 646.000 149.280 ;
        RECT 4.000 139.080 646.000 147.880 ;
        RECT 4.400 137.680 646.000 139.080 ;
        RECT 4.000 128.880 646.000 137.680 ;
        RECT 4.400 128.200 646.000 128.880 ;
        RECT 4.400 127.480 645.600 128.200 ;
        RECT 4.000 126.800 645.600 127.480 ;
        RECT 4.000 118.680 646.000 126.800 ;
        RECT 4.400 117.280 646.000 118.680 ;
        RECT 4.000 108.480 646.000 117.280 ;
        RECT 4.400 107.080 646.000 108.480 ;
        RECT 4.000 100.320 646.000 107.080 ;
        RECT 4.000 98.920 645.600 100.320 ;
        RECT 4.000 98.280 646.000 98.920 ;
        RECT 4.400 96.880 646.000 98.280 ;
        RECT 4.000 88.080 646.000 96.880 ;
        RECT 4.400 86.680 646.000 88.080 ;
        RECT 4.000 77.880 646.000 86.680 ;
        RECT 4.400 76.480 646.000 77.880 ;
        RECT 4.000 72.440 646.000 76.480 ;
        RECT 4.000 71.040 645.600 72.440 ;
        RECT 4.000 67.680 646.000 71.040 ;
        RECT 4.400 66.280 646.000 67.680 ;
        RECT 4.000 57.480 646.000 66.280 ;
        RECT 4.400 56.080 646.000 57.480 ;
        RECT 4.000 47.280 646.000 56.080 ;
        RECT 4.400 45.880 646.000 47.280 ;
        RECT 4.000 44.560 646.000 45.880 ;
        RECT 4.000 43.160 645.600 44.560 ;
        RECT 4.000 37.080 646.000 43.160 ;
        RECT 4.400 35.680 646.000 37.080 ;
        RECT 4.000 26.880 646.000 35.680 ;
        RECT 4.400 25.480 646.000 26.880 ;
        RECT 4.000 16.680 646.000 25.480 ;
        RECT 4.400 15.280 645.600 16.680 ;
        RECT 4.000 9.015 646.000 15.280 ;
      LAYER met4 ;
        RECT 8.575 12.415 20.640 436.385 ;
        RECT 23.040 12.415 97.440 436.385 ;
        RECT 99.840 12.415 174.240 436.385 ;
        RECT 176.640 12.415 251.040 436.385 ;
        RECT 253.440 12.415 327.840 436.385 ;
        RECT 330.240 12.415 404.640 436.385 ;
        RECT 407.040 12.415 481.440 436.385 ;
        RECT 483.840 12.415 558.240 436.385 ;
        RECT 560.640 12.415 593.105 436.385 ;
  END
END wrapped_tms1x00
END LIBRARY

