VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tms1x00_ram
  CLASS BLOCK ;
  FOREIGN tms1x00_ram ;
  ORIGIN 0.000 0.000 ;
  SIZE 256.000 BY 256.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 252.000 191.730 256.000 ;
    END
  END clk
  PIN r_val[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.200 4.000 195.800 ;
    END
  END r_val[0]
  PIN r_val[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.200 4.000 212.800 ;
    END
  END r_val[1]
  PIN r_val[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.200 4.000 229.800 ;
    END
  END r_val[2]
  PIN r_val[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.200 4.000 246.800 ;
    END
  END r_val[3]
  PIN ram_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 4.000 8.800 ;
    END
  END ram_addr[0]
  PIN ram_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 4.000 25.800 ;
    END
  END ram_addr[1]
  PIN ram_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END ram_addr[2]
  PIN ram_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 4.000 59.800 ;
    END
  END ram_addr[3]
  PIN ram_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 4.000 76.800 ;
    END
  END ram_addr[4]
  PIN ram_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.200 4.000 93.800 ;
    END
  END ram_addr[5]
  PIN ram_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 4.000 110.800 ;
    END
  END ram_addr[6]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 245.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 245.040 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 245.040 ;
    END
  END vssd1
  PIN w_val[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.200 4.000 127.800 ;
    END
  END w_val[0]
  PIN w_val[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.200 4.000 144.800 ;
    END
  END w_val[1]
  PIN w_val[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.200 4.000 161.800 ;
    END
  END w_val[2]
  PIN w_val[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 4.000 178.800 ;
    END
  END w_val[3]
  PIN wen
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 252.000 63.850 256.000 ;
    END
  END wen
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 250.240 244.885 ;
      LAYER met1 ;
        RECT 4.670 10.640 250.240 245.040 ;
      LAYER met2 ;
        RECT 4.690 251.720 63.290 252.000 ;
        RECT 64.130 251.720 191.170 252.000 ;
        RECT 192.010 251.720 222.080 252.000 ;
        RECT 4.690 8.315 222.080 251.720 ;
      LAYER met3 ;
        RECT 4.400 245.800 203.255 246.665 ;
        RECT 4.000 230.200 203.255 245.800 ;
        RECT 4.400 228.800 203.255 230.200 ;
        RECT 4.000 213.200 203.255 228.800 ;
        RECT 4.400 211.800 203.255 213.200 ;
        RECT 4.000 196.200 203.255 211.800 ;
        RECT 4.400 194.800 203.255 196.200 ;
        RECT 4.000 179.200 203.255 194.800 ;
        RECT 4.400 177.800 203.255 179.200 ;
        RECT 4.000 162.200 203.255 177.800 ;
        RECT 4.400 160.800 203.255 162.200 ;
        RECT 4.000 145.200 203.255 160.800 ;
        RECT 4.400 143.800 203.255 145.200 ;
        RECT 4.000 128.200 203.255 143.800 ;
        RECT 4.400 126.800 203.255 128.200 ;
        RECT 4.000 111.200 203.255 126.800 ;
        RECT 4.400 109.800 203.255 111.200 ;
        RECT 4.000 94.200 203.255 109.800 ;
        RECT 4.400 92.800 203.255 94.200 ;
        RECT 4.000 77.200 203.255 92.800 ;
        RECT 4.400 75.800 203.255 77.200 ;
        RECT 4.000 60.200 203.255 75.800 ;
        RECT 4.400 58.800 203.255 60.200 ;
        RECT 4.000 43.200 203.255 58.800 ;
        RECT 4.400 41.800 203.255 43.200 ;
        RECT 4.000 26.200 203.255 41.800 ;
        RECT 4.400 24.800 203.255 26.200 ;
        RECT 4.000 9.200 203.255 24.800 ;
        RECT 4.400 8.335 203.255 9.200 ;
      LAYER met4 ;
        RECT 35.255 47.775 97.440 237.825 ;
        RECT 99.840 47.775 174.240 237.825 ;
        RECT 176.640 47.775 191.985 237.825 ;
  END
END tms1x00_ram
END LIBRARY

