// This is the unpowered netlist.
module wrapped_tms1x00 (oram_csb,
    ram_csb,
    ram_web,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    io_in,
    io_oeb,
    io_out,
    oram_addr,
    oram_value,
    ram_adrb,
    ram_val,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o);
 output oram_csb;
 output ram_csb;
 output ram_web;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 output [8:0] oram_addr;
 input [31:0] oram_value;
 output [8:0] ram_adrb;
 input [31:0] ram_val;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;

 wire \K_override[0] ;
 wire \K_override[1] ;
 wire \K_override[2] ;
 wire \K_override[3] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire chip_sel_override;
 wire feedback_delay;
 wire net191;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net192;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net193;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire clknet_leaf_0_wb_clk_i;
 wire net178;
 wire net179;
 wire net180;
 wire net188;
 wire net189;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net190;
 wire \tms1x00.A[0] ;
 wire \tms1x00.A[1] ;
 wire \tms1x00.A[2] ;
 wire \tms1x00.A[3] ;
 wire \tms1x00.CL ;
 wire \tms1x00.K_in[0] ;
 wire \tms1x00.K_in[1] ;
 wire \tms1x00.K_in[2] ;
 wire \tms1x00.K_in[3] ;
 wire \tms1x00.K_latch[0] ;
 wire \tms1x00.K_latch[1] ;
 wire \tms1x00.K_latch[2] ;
 wire \tms1x00.K_latch[3] ;
 wire \tms1x00.N[0] ;
 wire \tms1x00.N[1] ;
 wire \tms1x00.N[2] ;
 wire \tms1x00.N[3] ;
 wire \tms1x00.PA[0] ;
 wire \tms1x00.PA[1] ;
 wire \tms1x00.PA[2] ;
 wire \tms1x00.PA[3] ;
 wire \tms1x00.PB[0] ;
 wire \tms1x00.PB[1] ;
 wire \tms1x00.PB[2] ;
 wire \tms1x00.PB[3] ;
 wire \tms1x00.PC[0] ;
 wire \tms1x00.PC[1] ;
 wire \tms1x00.PC[2] ;
 wire \tms1x00.PC[3] ;
 wire \tms1x00.PC[4] ;
 wire \tms1x00.PC[5] ;
 wire \tms1x00.P[0] ;
 wire \tms1x00.P[1] ;
 wire \tms1x00.P[2] ;
 wire \tms1x00.P[3] ;
 wire \tms1x00.RAM[0][0] ;
 wire \tms1x00.RAM[0][1] ;
 wire \tms1x00.RAM[0][2] ;
 wire \tms1x00.RAM[0][3] ;
 wire \tms1x00.RAM[100][0] ;
 wire \tms1x00.RAM[100][1] ;
 wire \tms1x00.RAM[100][2] ;
 wire \tms1x00.RAM[100][3] ;
 wire \tms1x00.RAM[101][0] ;
 wire \tms1x00.RAM[101][1] ;
 wire \tms1x00.RAM[101][2] ;
 wire \tms1x00.RAM[101][3] ;
 wire \tms1x00.RAM[102][0] ;
 wire \tms1x00.RAM[102][1] ;
 wire \tms1x00.RAM[102][2] ;
 wire \tms1x00.RAM[102][3] ;
 wire \tms1x00.RAM[103][0] ;
 wire \tms1x00.RAM[103][1] ;
 wire \tms1x00.RAM[103][2] ;
 wire \tms1x00.RAM[103][3] ;
 wire \tms1x00.RAM[104][0] ;
 wire \tms1x00.RAM[104][1] ;
 wire \tms1x00.RAM[104][2] ;
 wire \tms1x00.RAM[104][3] ;
 wire \tms1x00.RAM[105][0] ;
 wire \tms1x00.RAM[105][1] ;
 wire \tms1x00.RAM[105][2] ;
 wire \tms1x00.RAM[105][3] ;
 wire \tms1x00.RAM[106][0] ;
 wire \tms1x00.RAM[106][1] ;
 wire \tms1x00.RAM[106][2] ;
 wire \tms1x00.RAM[106][3] ;
 wire \tms1x00.RAM[107][0] ;
 wire \tms1x00.RAM[107][1] ;
 wire \tms1x00.RAM[107][2] ;
 wire \tms1x00.RAM[107][3] ;
 wire \tms1x00.RAM[108][0] ;
 wire \tms1x00.RAM[108][1] ;
 wire \tms1x00.RAM[108][2] ;
 wire \tms1x00.RAM[108][3] ;
 wire \tms1x00.RAM[109][0] ;
 wire \tms1x00.RAM[109][1] ;
 wire \tms1x00.RAM[109][2] ;
 wire \tms1x00.RAM[109][3] ;
 wire \tms1x00.RAM[10][0] ;
 wire \tms1x00.RAM[10][1] ;
 wire \tms1x00.RAM[10][2] ;
 wire \tms1x00.RAM[10][3] ;
 wire \tms1x00.RAM[110][0] ;
 wire \tms1x00.RAM[110][1] ;
 wire \tms1x00.RAM[110][2] ;
 wire \tms1x00.RAM[110][3] ;
 wire \tms1x00.RAM[111][0] ;
 wire \tms1x00.RAM[111][1] ;
 wire \tms1x00.RAM[111][2] ;
 wire \tms1x00.RAM[111][3] ;
 wire \tms1x00.RAM[112][0] ;
 wire \tms1x00.RAM[112][1] ;
 wire \tms1x00.RAM[112][2] ;
 wire \tms1x00.RAM[112][3] ;
 wire \tms1x00.RAM[113][0] ;
 wire \tms1x00.RAM[113][1] ;
 wire \tms1x00.RAM[113][2] ;
 wire \tms1x00.RAM[113][3] ;
 wire \tms1x00.RAM[114][0] ;
 wire \tms1x00.RAM[114][1] ;
 wire \tms1x00.RAM[114][2] ;
 wire \tms1x00.RAM[114][3] ;
 wire \tms1x00.RAM[115][0] ;
 wire \tms1x00.RAM[115][1] ;
 wire \tms1x00.RAM[115][2] ;
 wire \tms1x00.RAM[115][3] ;
 wire \tms1x00.RAM[116][0] ;
 wire \tms1x00.RAM[116][1] ;
 wire \tms1x00.RAM[116][2] ;
 wire \tms1x00.RAM[116][3] ;
 wire \tms1x00.RAM[117][0] ;
 wire \tms1x00.RAM[117][1] ;
 wire \tms1x00.RAM[117][2] ;
 wire \tms1x00.RAM[117][3] ;
 wire \tms1x00.RAM[118][0] ;
 wire \tms1x00.RAM[118][1] ;
 wire \tms1x00.RAM[118][2] ;
 wire \tms1x00.RAM[118][3] ;
 wire \tms1x00.RAM[119][0] ;
 wire \tms1x00.RAM[119][1] ;
 wire \tms1x00.RAM[119][2] ;
 wire \tms1x00.RAM[119][3] ;
 wire \tms1x00.RAM[11][0] ;
 wire \tms1x00.RAM[11][1] ;
 wire \tms1x00.RAM[11][2] ;
 wire \tms1x00.RAM[11][3] ;
 wire \tms1x00.RAM[120][0] ;
 wire \tms1x00.RAM[120][1] ;
 wire \tms1x00.RAM[120][2] ;
 wire \tms1x00.RAM[120][3] ;
 wire \tms1x00.RAM[121][0] ;
 wire \tms1x00.RAM[121][1] ;
 wire \tms1x00.RAM[121][2] ;
 wire \tms1x00.RAM[121][3] ;
 wire \tms1x00.RAM[122][0] ;
 wire \tms1x00.RAM[122][1] ;
 wire \tms1x00.RAM[122][2] ;
 wire \tms1x00.RAM[122][3] ;
 wire \tms1x00.RAM[123][0] ;
 wire \tms1x00.RAM[123][1] ;
 wire \tms1x00.RAM[123][2] ;
 wire \tms1x00.RAM[123][3] ;
 wire \tms1x00.RAM[124][0] ;
 wire \tms1x00.RAM[124][1] ;
 wire \tms1x00.RAM[124][2] ;
 wire \tms1x00.RAM[124][3] ;
 wire \tms1x00.RAM[125][0] ;
 wire \tms1x00.RAM[125][1] ;
 wire \tms1x00.RAM[125][2] ;
 wire \tms1x00.RAM[125][3] ;
 wire \tms1x00.RAM[126][0] ;
 wire \tms1x00.RAM[126][1] ;
 wire \tms1x00.RAM[126][2] ;
 wire \tms1x00.RAM[126][3] ;
 wire \tms1x00.RAM[127][0] ;
 wire \tms1x00.RAM[127][1] ;
 wire \tms1x00.RAM[127][2] ;
 wire \tms1x00.RAM[127][3] ;
 wire \tms1x00.RAM[12][0] ;
 wire \tms1x00.RAM[12][1] ;
 wire \tms1x00.RAM[12][2] ;
 wire \tms1x00.RAM[12][3] ;
 wire \tms1x00.RAM[13][0] ;
 wire \tms1x00.RAM[13][1] ;
 wire \tms1x00.RAM[13][2] ;
 wire \tms1x00.RAM[13][3] ;
 wire \tms1x00.RAM[14][0] ;
 wire \tms1x00.RAM[14][1] ;
 wire \tms1x00.RAM[14][2] ;
 wire \tms1x00.RAM[14][3] ;
 wire \tms1x00.RAM[15][0] ;
 wire \tms1x00.RAM[15][1] ;
 wire \tms1x00.RAM[15][2] ;
 wire \tms1x00.RAM[15][3] ;
 wire \tms1x00.RAM[16][0] ;
 wire \tms1x00.RAM[16][1] ;
 wire \tms1x00.RAM[16][2] ;
 wire \tms1x00.RAM[16][3] ;
 wire \tms1x00.RAM[17][0] ;
 wire \tms1x00.RAM[17][1] ;
 wire \tms1x00.RAM[17][2] ;
 wire \tms1x00.RAM[17][3] ;
 wire \tms1x00.RAM[18][0] ;
 wire \tms1x00.RAM[18][1] ;
 wire \tms1x00.RAM[18][2] ;
 wire \tms1x00.RAM[18][3] ;
 wire \tms1x00.RAM[19][0] ;
 wire \tms1x00.RAM[19][1] ;
 wire \tms1x00.RAM[19][2] ;
 wire \tms1x00.RAM[19][3] ;
 wire \tms1x00.RAM[1][0] ;
 wire \tms1x00.RAM[1][1] ;
 wire \tms1x00.RAM[1][2] ;
 wire \tms1x00.RAM[1][3] ;
 wire \tms1x00.RAM[20][0] ;
 wire \tms1x00.RAM[20][1] ;
 wire \tms1x00.RAM[20][2] ;
 wire \tms1x00.RAM[20][3] ;
 wire \tms1x00.RAM[21][0] ;
 wire \tms1x00.RAM[21][1] ;
 wire \tms1x00.RAM[21][2] ;
 wire \tms1x00.RAM[21][3] ;
 wire \tms1x00.RAM[22][0] ;
 wire \tms1x00.RAM[22][1] ;
 wire \tms1x00.RAM[22][2] ;
 wire \tms1x00.RAM[22][3] ;
 wire \tms1x00.RAM[23][0] ;
 wire \tms1x00.RAM[23][1] ;
 wire \tms1x00.RAM[23][2] ;
 wire \tms1x00.RAM[23][3] ;
 wire \tms1x00.RAM[24][0] ;
 wire \tms1x00.RAM[24][1] ;
 wire \tms1x00.RAM[24][2] ;
 wire \tms1x00.RAM[24][3] ;
 wire \tms1x00.RAM[25][0] ;
 wire \tms1x00.RAM[25][1] ;
 wire \tms1x00.RAM[25][2] ;
 wire \tms1x00.RAM[25][3] ;
 wire \tms1x00.RAM[26][0] ;
 wire \tms1x00.RAM[26][1] ;
 wire \tms1x00.RAM[26][2] ;
 wire \tms1x00.RAM[26][3] ;
 wire \tms1x00.RAM[27][0] ;
 wire \tms1x00.RAM[27][1] ;
 wire \tms1x00.RAM[27][2] ;
 wire \tms1x00.RAM[27][3] ;
 wire \tms1x00.RAM[28][0] ;
 wire \tms1x00.RAM[28][1] ;
 wire \tms1x00.RAM[28][2] ;
 wire \tms1x00.RAM[28][3] ;
 wire \tms1x00.RAM[29][0] ;
 wire \tms1x00.RAM[29][1] ;
 wire \tms1x00.RAM[29][2] ;
 wire \tms1x00.RAM[29][3] ;
 wire \tms1x00.RAM[2][0] ;
 wire \tms1x00.RAM[2][1] ;
 wire \tms1x00.RAM[2][2] ;
 wire \tms1x00.RAM[2][3] ;
 wire \tms1x00.RAM[30][0] ;
 wire \tms1x00.RAM[30][1] ;
 wire \tms1x00.RAM[30][2] ;
 wire \tms1x00.RAM[30][3] ;
 wire \tms1x00.RAM[31][0] ;
 wire \tms1x00.RAM[31][1] ;
 wire \tms1x00.RAM[31][2] ;
 wire \tms1x00.RAM[31][3] ;
 wire \tms1x00.RAM[32][0] ;
 wire \tms1x00.RAM[32][1] ;
 wire \tms1x00.RAM[32][2] ;
 wire \tms1x00.RAM[32][3] ;
 wire \tms1x00.RAM[33][0] ;
 wire \tms1x00.RAM[33][1] ;
 wire \tms1x00.RAM[33][2] ;
 wire \tms1x00.RAM[33][3] ;
 wire \tms1x00.RAM[34][0] ;
 wire \tms1x00.RAM[34][1] ;
 wire \tms1x00.RAM[34][2] ;
 wire \tms1x00.RAM[34][3] ;
 wire \tms1x00.RAM[35][0] ;
 wire \tms1x00.RAM[35][1] ;
 wire \tms1x00.RAM[35][2] ;
 wire \tms1x00.RAM[35][3] ;
 wire \tms1x00.RAM[36][0] ;
 wire \tms1x00.RAM[36][1] ;
 wire \tms1x00.RAM[36][2] ;
 wire \tms1x00.RAM[36][3] ;
 wire \tms1x00.RAM[37][0] ;
 wire \tms1x00.RAM[37][1] ;
 wire \tms1x00.RAM[37][2] ;
 wire \tms1x00.RAM[37][3] ;
 wire \tms1x00.RAM[38][0] ;
 wire \tms1x00.RAM[38][1] ;
 wire \tms1x00.RAM[38][2] ;
 wire \tms1x00.RAM[38][3] ;
 wire \tms1x00.RAM[39][0] ;
 wire \tms1x00.RAM[39][1] ;
 wire \tms1x00.RAM[39][2] ;
 wire \tms1x00.RAM[39][3] ;
 wire \tms1x00.RAM[3][0] ;
 wire \tms1x00.RAM[3][1] ;
 wire \tms1x00.RAM[3][2] ;
 wire \tms1x00.RAM[3][3] ;
 wire \tms1x00.RAM[40][0] ;
 wire \tms1x00.RAM[40][1] ;
 wire \tms1x00.RAM[40][2] ;
 wire \tms1x00.RAM[40][3] ;
 wire \tms1x00.RAM[41][0] ;
 wire \tms1x00.RAM[41][1] ;
 wire \tms1x00.RAM[41][2] ;
 wire \tms1x00.RAM[41][3] ;
 wire \tms1x00.RAM[42][0] ;
 wire \tms1x00.RAM[42][1] ;
 wire \tms1x00.RAM[42][2] ;
 wire \tms1x00.RAM[42][3] ;
 wire \tms1x00.RAM[43][0] ;
 wire \tms1x00.RAM[43][1] ;
 wire \tms1x00.RAM[43][2] ;
 wire \tms1x00.RAM[43][3] ;
 wire \tms1x00.RAM[44][0] ;
 wire \tms1x00.RAM[44][1] ;
 wire \tms1x00.RAM[44][2] ;
 wire \tms1x00.RAM[44][3] ;
 wire \tms1x00.RAM[45][0] ;
 wire \tms1x00.RAM[45][1] ;
 wire \tms1x00.RAM[45][2] ;
 wire \tms1x00.RAM[45][3] ;
 wire \tms1x00.RAM[46][0] ;
 wire \tms1x00.RAM[46][1] ;
 wire \tms1x00.RAM[46][2] ;
 wire \tms1x00.RAM[46][3] ;
 wire \tms1x00.RAM[47][0] ;
 wire \tms1x00.RAM[47][1] ;
 wire \tms1x00.RAM[47][2] ;
 wire \tms1x00.RAM[47][3] ;
 wire \tms1x00.RAM[48][0] ;
 wire \tms1x00.RAM[48][1] ;
 wire \tms1x00.RAM[48][2] ;
 wire \tms1x00.RAM[48][3] ;
 wire \tms1x00.RAM[49][0] ;
 wire \tms1x00.RAM[49][1] ;
 wire \tms1x00.RAM[49][2] ;
 wire \tms1x00.RAM[49][3] ;
 wire \tms1x00.RAM[4][0] ;
 wire \tms1x00.RAM[4][1] ;
 wire \tms1x00.RAM[4][2] ;
 wire \tms1x00.RAM[4][3] ;
 wire \tms1x00.RAM[50][0] ;
 wire \tms1x00.RAM[50][1] ;
 wire \tms1x00.RAM[50][2] ;
 wire \tms1x00.RAM[50][3] ;
 wire \tms1x00.RAM[51][0] ;
 wire \tms1x00.RAM[51][1] ;
 wire \tms1x00.RAM[51][2] ;
 wire \tms1x00.RAM[51][3] ;
 wire \tms1x00.RAM[52][0] ;
 wire \tms1x00.RAM[52][1] ;
 wire \tms1x00.RAM[52][2] ;
 wire \tms1x00.RAM[52][3] ;
 wire \tms1x00.RAM[53][0] ;
 wire \tms1x00.RAM[53][1] ;
 wire \tms1x00.RAM[53][2] ;
 wire \tms1x00.RAM[53][3] ;
 wire \tms1x00.RAM[54][0] ;
 wire \tms1x00.RAM[54][1] ;
 wire \tms1x00.RAM[54][2] ;
 wire \tms1x00.RAM[54][3] ;
 wire \tms1x00.RAM[55][0] ;
 wire \tms1x00.RAM[55][1] ;
 wire \tms1x00.RAM[55][2] ;
 wire \tms1x00.RAM[55][3] ;
 wire \tms1x00.RAM[56][0] ;
 wire \tms1x00.RAM[56][1] ;
 wire \tms1x00.RAM[56][2] ;
 wire \tms1x00.RAM[56][3] ;
 wire \tms1x00.RAM[57][0] ;
 wire \tms1x00.RAM[57][1] ;
 wire \tms1x00.RAM[57][2] ;
 wire \tms1x00.RAM[57][3] ;
 wire \tms1x00.RAM[58][0] ;
 wire \tms1x00.RAM[58][1] ;
 wire \tms1x00.RAM[58][2] ;
 wire \tms1x00.RAM[58][3] ;
 wire \tms1x00.RAM[59][0] ;
 wire \tms1x00.RAM[59][1] ;
 wire \tms1x00.RAM[59][2] ;
 wire \tms1x00.RAM[59][3] ;
 wire \tms1x00.RAM[5][0] ;
 wire \tms1x00.RAM[5][1] ;
 wire \tms1x00.RAM[5][2] ;
 wire \tms1x00.RAM[5][3] ;
 wire \tms1x00.RAM[60][0] ;
 wire \tms1x00.RAM[60][1] ;
 wire \tms1x00.RAM[60][2] ;
 wire \tms1x00.RAM[60][3] ;
 wire \tms1x00.RAM[61][0] ;
 wire \tms1x00.RAM[61][1] ;
 wire \tms1x00.RAM[61][2] ;
 wire \tms1x00.RAM[61][3] ;
 wire \tms1x00.RAM[62][0] ;
 wire \tms1x00.RAM[62][1] ;
 wire \tms1x00.RAM[62][2] ;
 wire \tms1x00.RAM[62][3] ;
 wire \tms1x00.RAM[63][0] ;
 wire \tms1x00.RAM[63][1] ;
 wire \tms1x00.RAM[63][2] ;
 wire \tms1x00.RAM[63][3] ;
 wire \tms1x00.RAM[64][0] ;
 wire \tms1x00.RAM[64][1] ;
 wire \tms1x00.RAM[64][2] ;
 wire \tms1x00.RAM[64][3] ;
 wire \tms1x00.RAM[65][0] ;
 wire \tms1x00.RAM[65][1] ;
 wire \tms1x00.RAM[65][2] ;
 wire \tms1x00.RAM[65][3] ;
 wire \tms1x00.RAM[66][0] ;
 wire \tms1x00.RAM[66][1] ;
 wire \tms1x00.RAM[66][2] ;
 wire \tms1x00.RAM[66][3] ;
 wire \tms1x00.RAM[67][0] ;
 wire \tms1x00.RAM[67][1] ;
 wire \tms1x00.RAM[67][2] ;
 wire \tms1x00.RAM[67][3] ;
 wire \tms1x00.RAM[68][0] ;
 wire \tms1x00.RAM[68][1] ;
 wire \tms1x00.RAM[68][2] ;
 wire \tms1x00.RAM[68][3] ;
 wire \tms1x00.RAM[69][0] ;
 wire \tms1x00.RAM[69][1] ;
 wire \tms1x00.RAM[69][2] ;
 wire \tms1x00.RAM[69][3] ;
 wire \tms1x00.RAM[6][0] ;
 wire \tms1x00.RAM[6][1] ;
 wire \tms1x00.RAM[6][2] ;
 wire \tms1x00.RAM[6][3] ;
 wire \tms1x00.RAM[70][0] ;
 wire \tms1x00.RAM[70][1] ;
 wire \tms1x00.RAM[70][2] ;
 wire \tms1x00.RAM[70][3] ;
 wire \tms1x00.RAM[71][0] ;
 wire \tms1x00.RAM[71][1] ;
 wire \tms1x00.RAM[71][2] ;
 wire \tms1x00.RAM[71][3] ;
 wire \tms1x00.RAM[72][0] ;
 wire \tms1x00.RAM[72][1] ;
 wire \tms1x00.RAM[72][2] ;
 wire \tms1x00.RAM[72][3] ;
 wire \tms1x00.RAM[73][0] ;
 wire \tms1x00.RAM[73][1] ;
 wire \tms1x00.RAM[73][2] ;
 wire \tms1x00.RAM[73][3] ;
 wire \tms1x00.RAM[74][0] ;
 wire \tms1x00.RAM[74][1] ;
 wire \tms1x00.RAM[74][2] ;
 wire \tms1x00.RAM[74][3] ;
 wire \tms1x00.RAM[75][0] ;
 wire \tms1x00.RAM[75][1] ;
 wire \tms1x00.RAM[75][2] ;
 wire \tms1x00.RAM[75][3] ;
 wire \tms1x00.RAM[76][0] ;
 wire \tms1x00.RAM[76][1] ;
 wire \tms1x00.RAM[76][2] ;
 wire \tms1x00.RAM[76][3] ;
 wire \tms1x00.RAM[77][0] ;
 wire \tms1x00.RAM[77][1] ;
 wire \tms1x00.RAM[77][2] ;
 wire \tms1x00.RAM[77][3] ;
 wire \tms1x00.RAM[78][0] ;
 wire \tms1x00.RAM[78][1] ;
 wire \tms1x00.RAM[78][2] ;
 wire \tms1x00.RAM[78][3] ;
 wire \tms1x00.RAM[79][0] ;
 wire \tms1x00.RAM[79][1] ;
 wire \tms1x00.RAM[79][2] ;
 wire \tms1x00.RAM[79][3] ;
 wire \tms1x00.RAM[7][0] ;
 wire \tms1x00.RAM[7][1] ;
 wire \tms1x00.RAM[7][2] ;
 wire \tms1x00.RAM[7][3] ;
 wire \tms1x00.RAM[80][0] ;
 wire \tms1x00.RAM[80][1] ;
 wire \tms1x00.RAM[80][2] ;
 wire \tms1x00.RAM[80][3] ;
 wire \tms1x00.RAM[81][0] ;
 wire \tms1x00.RAM[81][1] ;
 wire \tms1x00.RAM[81][2] ;
 wire \tms1x00.RAM[81][3] ;
 wire \tms1x00.RAM[82][0] ;
 wire \tms1x00.RAM[82][1] ;
 wire \tms1x00.RAM[82][2] ;
 wire \tms1x00.RAM[82][3] ;
 wire \tms1x00.RAM[83][0] ;
 wire \tms1x00.RAM[83][1] ;
 wire \tms1x00.RAM[83][2] ;
 wire \tms1x00.RAM[83][3] ;
 wire \tms1x00.RAM[84][0] ;
 wire \tms1x00.RAM[84][1] ;
 wire \tms1x00.RAM[84][2] ;
 wire \tms1x00.RAM[84][3] ;
 wire \tms1x00.RAM[85][0] ;
 wire \tms1x00.RAM[85][1] ;
 wire \tms1x00.RAM[85][2] ;
 wire \tms1x00.RAM[85][3] ;
 wire \tms1x00.RAM[86][0] ;
 wire \tms1x00.RAM[86][1] ;
 wire \tms1x00.RAM[86][2] ;
 wire \tms1x00.RAM[86][3] ;
 wire \tms1x00.RAM[87][0] ;
 wire \tms1x00.RAM[87][1] ;
 wire \tms1x00.RAM[87][2] ;
 wire \tms1x00.RAM[87][3] ;
 wire \tms1x00.RAM[88][0] ;
 wire \tms1x00.RAM[88][1] ;
 wire \tms1x00.RAM[88][2] ;
 wire \tms1x00.RAM[88][3] ;
 wire \tms1x00.RAM[89][0] ;
 wire \tms1x00.RAM[89][1] ;
 wire \tms1x00.RAM[89][2] ;
 wire \tms1x00.RAM[89][3] ;
 wire \tms1x00.RAM[8][0] ;
 wire \tms1x00.RAM[8][1] ;
 wire \tms1x00.RAM[8][2] ;
 wire \tms1x00.RAM[8][3] ;
 wire \tms1x00.RAM[90][0] ;
 wire \tms1x00.RAM[90][1] ;
 wire \tms1x00.RAM[90][2] ;
 wire \tms1x00.RAM[90][3] ;
 wire \tms1x00.RAM[91][0] ;
 wire \tms1x00.RAM[91][1] ;
 wire \tms1x00.RAM[91][2] ;
 wire \tms1x00.RAM[91][3] ;
 wire \tms1x00.RAM[92][0] ;
 wire \tms1x00.RAM[92][1] ;
 wire \tms1x00.RAM[92][2] ;
 wire \tms1x00.RAM[92][3] ;
 wire \tms1x00.RAM[93][0] ;
 wire \tms1x00.RAM[93][1] ;
 wire \tms1x00.RAM[93][2] ;
 wire \tms1x00.RAM[93][3] ;
 wire \tms1x00.RAM[94][0] ;
 wire \tms1x00.RAM[94][1] ;
 wire \tms1x00.RAM[94][2] ;
 wire \tms1x00.RAM[94][3] ;
 wire \tms1x00.RAM[95][0] ;
 wire \tms1x00.RAM[95][1] ;
 wire \tms1x00.RAM[95][2] ;
 wire \tms1x00.RAM[95][3] ;
 wire \tms1x00.RAM[96][0] ;
 wire \tms1x00.RAM[96][1] ;
 wire \tms1x00.RAM[96][2] ;
 wire \tms1x00.RAM[96][3] ;
 wire \tms1x00.RAM[97][0] ;
 wire \tms1x00.RAM[97][1] ;
 wire \tms1x00.RAM[97][2] ;
 wire \tms1x00.RAM[97][3] ;
 wire \tms1x00.RAM[98][0] ;
 wire \tms1x00.RAM[98][1] ;
 wire \tms1x00.RAM[98][2] ;
 wire \tms1x00.RAM[98][3] ;
 wire \tms1x00.RAM[99][0] ;
 wire \tms1x00.RAM[99][1] ;
 wire \tms1x00.RAM[99][2] ;
 wire \tms1x00.RAM[99][3] ;
 wire \tms1x00.RAM[9][0] ;
 wire \tms1x00.RAM[9][1] ;
 wire \tms1x00.RAM[9][2] ;
 wire \tms1x00.RAM[9][3] ;
 wire \tms1x00.SR[0] ;
 wire \tms1x00.SR[1] ;
 wire \tms1x00.SR[2] ;
 wire \tms1x00.SR[3] ;
 wire \tms1x00.SR[4] ;
 wire \tms1x00.SR[5] ;
 wire \tms1x00.X[0] ;
 wire \tms1x00.X[1] ;
 wire \tms1x00.X[2] ;
 wire \tms1x00.Y[0] ;
 wire \tms1x00.Y[1] ;
 wire \tms1x00.Y[2] ;
 wire \tms1x00.Y[3] ;
 wire \tms1x00.ins_in[0] ;
 wire \tms1x00.ins_in[1] ;
 wire \tms1x00.ins_in[2] ;
 wire \tms1x00.ins_in[3] ;
 wire \tms1x00.ins_in[4] ;
 wire \tms1x00.ins_in[5] ;
 wire \tms1x00.ins_in[6] ;
 wire \tms1x00.ins_in[7] ;
 wire \tms1x00.ram_addr_buff[0] ;
 wire \tms1x00.ram_addr_buff[1] ;
 wire \tms1x00.ram_addr_buff[2] ;
 wire \tms1x00.ram_addr_buff[3] ;
 wire \tms1x00.ram_addr_buff[4] ;
 wire \tms1x00.ram_addr_buff[5] ;
 wire \tms1x00.ram_addr_buff[6] ;
 wire \tms1x00.status ;
 wire \tms1x00.wb_step ;
 wire \tms1x00.wb_step_state ;
 wire valid;
 wire wb_rst_override;
 wire \wbs_o_buff[0] ;
 wire \wbs_o_buff[10] ;
 wire \wbs_o_buff[11] ;
 wire \wbs_o_buff[12] ;
 wire \wbs_o_buff[13] ;
 wire \wbs_o_buff[14] ;
 wire \wbs_o_buff[15] ;
 wire \wbs_o_buff[16] ;
 wire \wbs_o_buff[17] ;
 wire \wbs_o_buff[18] ;
 wire \wbs_o_buff[19] ;
 wire \wbs_o_buff[1] ;
 wire \wbs_o_buff[20] ;
 wire \wbs_o_buff[21] ;
 wire \wbs_o_buff[22] ;
 wire \wbs_o_buff[23] ;
 wire \wbs_o_buff[24] ;
 wire \wbs_o_buff[25] ;
 wire \wbs_o_buff[26] ;
 wire \wbs_o_buff[27] ;
 wire \wbs_o_buff[28] ;
 wire \wbs_o_buff[29] ;
 wire \wbs_o_buff[2] ;
 wire \wbs_o_buff[30] ;
 wire \wbs_o_buff[31] ;
 wire \wbs_o_buff[3] ;
 wire \wbs_o_buff[4] ;
 wire \wbs_o_buff[5] ;
 wire \wbs_o_buff[6] ;
 wire \wbs_o_buff[7] ;
 wire \wbs_o_buff[8] ;
 wire \wbs_o_buff[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire clknet_leaf_1_wb_clk_i;
 wire clknet_leaf_2_wb_clk_i;
 wire clknet_leaf_3_wb_clk_i;
 wire clknet_leaf_4_wb_clk_i;
 wire clknet_leaf_5_wb_clk_i;
 wire clknet_leaf_6_wb_clk_i;
 wire clknet_leaf_7_wb_clk_i;
 wire clknet_leaf_8_wb_clk_i;
 wire clknet_leaf_9_wb_clk_i;
 wire clknet_leaf_10_wb_clk_i;
 wire clknet_leaf_11_wb_clk_i;
 wire clknet_leaf_12_wb_clk_i;
 wire clknet_leaf_13_wb_clk_i;
 wire clknet_leaf_14_wb_clk_i;
 wire clknet_leaf_15_wb_clk_i;
 wire clknet_leaf_16_wb_clk_i;
 wire clknet_leaf_17_wb_clk_i;
 wire clknet_leaf_18_wb_clk_i;
 wire clknet_leaf_19_wb_clk_i;
 wire clknet_leaf_20_wb_clk_i;
 wire clknet_leaf_21_wb_clk_i;
 wire clknet_leaf_22_wb_clk_i;
 wire clknet_leaf_23_wb_clk_i;
 wire clknet_leaf_24_wb_clk_i;
 wire clknet_leaf_25_wb_clk_i;
 wire clknet_leaf_26_wb_clk_i;
 wire clknet_leaf_27_wb_clk_i;
 wire clknet_leaf_28_wb_clk_i;
 wire clknet_leaf_29_wb_clk_i;
 wire clknet_leaf_30_wb_clk_i;
 wire clknet_leaf_31_wb_clk_i;
 wire clknet_leaf_32_wb_clk_i;
 wire clknet_leaf_33_wb_clk_i;
 wire clknet_leaf_34_wb_clk_i;
 wire clknet_leaf_35_wb_clk_i;
 wire clknet_0_wb_clk_i;
 wire clknet_2_0__leaf_wb_clk_i;
 wire clknet_2_1__leaf_wb_clk_i;
 wire clknet_2_2__leaf_wb_clk_i;
 wire clknet_2_3__leaf_wb_clk_i;
 wire net200;

 sky130_fd_sc_hd__and2_1 _2179_ (.A(net67),
    .B(net58),
    .X(_0656_));
 sky130_fd_sc_hd__clkbuf_2 _2180_ (.A(_0656_),
    .X(valid));
 sky130_fd_sc_hd__clkbuf_4 _2181_ (.A(net49),
    .X(_0657_));
 sky130_fd_sc_hd__mux2_1 _2182_ (.A0(net14),
    .A1(\wbs_o_buff[0] ),
    .S(_0657_),
    .X(_0658_));
 sky130_fd_sc_hd__clkbuf_1 _2183_ (.A(_0658_),
    .X(net116));
 sky130_fd_sc_hd__mux2_1 _2184_ (.A0(net25),
    .A1(\wbs_o_buff[1] ),
    .S(_0657_),
    .X(_0659_));
 sky130_fd_sc_hd__clkbuf_1 _2185_ (.A(_0659_),
    .X(net127));
 sky130_fd_sc_hd__mux2_1 _2186_ (.A0(net36),
    .A1(\wbs_o_buff[2] ),
    .S(_0657_),
    .X(_0660_));
 sky130_fd_sc_hd__clkbuf_1 _2187_ (.A(_0660_),
    .X(net138));
 sky130_fd_sc_hd__mux2_1 _2188_ (.A0(net39),
    .A1(\wbs_o_buff[3] ),
    .S(_0657_),
    .X(_0661_));
 sky130_fd_sc_hd__clkbuf_1 _2189_ (.A(_0661_),
    .X(net141));
 sky130_fd_sc_hd__mux2_1 _2190_ (.A0(net40),
    .A1(\wbs_o_buff[4] ),
    .S(_0657_),
    .X(_0662_));
 sky130_fd_sc_hd__clkbuf_1 _2191_ (.A(_0662_),
    .X(net142));
 sky130_fd_sc_hd__mux2_1 _2192_ (.A0(net41),
    .A1(\wbs_o_buff[5] ),
    .S(_0657_),
    .X(_0663_));
 sky130_fd_sc_hd__clkbuf_1 _2193_ (.A(_0663_),
    .X(net143));
 sky130_fd_sc_hd__mux2_1 _2194_ (.A0(net42),
    .A1(\wbs_o_buff[6] ),
    .S(_0657_),
    .X(_0664_));
 sky130_fd_sc_hd__clkbuf_1 _2195_ (.A(_0664_),
    .X(net144));
 sky130_fd_sc_hd__mux2_1 _2196_ (.A0(net43),
    .A1(\wbs_o_buff[7] ),
    .S(_0657_),
    .X(_0665_));
 sky130_fd_sc_hd__clkbuf_1 _2197_ (.A(_0665_),
    .X(net145));
 sky130_fd_sc_hd__mux2_1 _2198_ (.A0(net44),
    .A1(\wbs_o_buff[8] ),
    .S(_0657_),
    .X(_0666_));
 sky130_fd_sc_hd__clkbuf_1 _2199_ (.A(_0666_),
    .X(net146));
 sky130_fd_sc_hd__mux2_1 _2200_ (.A0(net45),
    .A1(\wbs_o_buff[9] ),
    .S(_0657_),
    .X(_0667_));
 sky130_fd_sc_hd__clkbuf_1 _2201_ (.A(_0667_),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_4 _2202_ (.A(net49),
    .X(_0668_));
 sky130_fd_sc_hd__mux2_1 _2203_ (.A0(net15),
    .A1(\wbs_o_buff[10] ),
    .S(_0668_),
    .X(_0669_));
 sky130_fd_sc_hd__clkbuf_1 _2204_ (.A(_0669_),
    .X(net117));
 sky130_fd_sc_hd__mux2_1 _2205_ (.A0(net16),
    .A1(\wbs_o_buff[11] ),
    .S(_0668_),
    .X(_0670_));
 sky130_fd_sc_hd__clkbuf_1 _2206_ (.A(_0670_),
    .X(net118));
 sky130_fd_sc_hd__mux2_1 _2207_ (.A0(net17),
    .A1(\wbs_o_buff[12] ),
    .S(_0668_),
    .X(_0671_));
 sky130_fd_sc_hd__clkbuf_1 _2208_ (.A(_0671_),
    .X(net119));
 sky130_fd_sc_hd__mux2_1 _2209_ (.A0(net18),
    .A1(\wbs_o_buff[13] ),
    .S(_0668_),
    .X(_0672_));
 sky130_fd_sc_hd__clkbuf_1 _2210_ (.A(_0672_),
    .X(net120));
 sky130_fd_sc_hd__mux2_1 _2211_ (.A0(net19),
    .A1(\wbs_o_buff[14] ),
    .S(_0668_),
    .X(_0673_));
 sky130_fd_sc_hd__clkbuf_1 _2212_ (.A(_0673_),
    .X(net121));
 sky130_fd_sc_hd__mux2_1 _2213_ (.A0(net20),
    .A1(\wbs_o_buff[15] ),
    .S(_0668_),
    .X(_0674_));
 sky130_fd_sc_hd__clkbuf_1 _2214_ (.A(_0674_),
    .X(net122));
 sky130_fd_sc_hd__mux2_1 _2215_ (.A0(net21),
    .A1(\wbs_o_buff[16] ),
    .S(_0668_),
    .X(_0675_));
 sky130_fd_sc_hd__clkbuf_1 _2216_ (.A(_0675_),
    .X(net123));
 sky130_fd_sc_hd__mux2_1 _2217_ (.A0(net22),
    .A1(\wbs_o_buff[17] ),
    .S(_0668_),
    .X(_0676_));
 sky130_fd_sc_hd__clkbuf_1 _2218_ (.A(_0676_),
    .X(net124));
 sky130_fd_sc_hd__mux2_1 _2219_ (.A0(net23),
    .A1(\wbs_o_buff[18] ),
    .S(_0668_),
    .X(_0677_));
 sky130_fd_sc_hd__clkbuf_1 _2220_ (.A(_0677_),
    .X(net125));
 sky130_fd_sc_hd__mux2_1 _2221_ (.A0(net24),
    .A1(\wbs_o_buff[19] ),
    .S(_0668_),
    .X(_0678_));
 sky130_fd_sc_hd__clkbuf_1 _2222_ (.A(_0678_),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_4 _2223_ (.A(net49),
    .X(_0679_));
 sky130_fd_sc_hd__mux2_1 _2224_ (.A0(net26),
    .A1(\wbs_o_buff[20] ),
    .S(_0679_),
    .X(_0680_));
 sky130_fd_sc_hd__clkbuf_1 _2225_ (.A(_0680_),
    .X(net128));
 sky130_fd_sc_hd__mux2_1 _2226_ (.A0(net27),
    .A1(\wbs_o_buff[21] ),
    .S(_0679_),
    .X(_0681_));
 sky130_fd_sc_hd__clkbuf_1 _2227_ (.A(_0681_),
    .X(net129));
 sky130_fd_sc_hd__mux2_1 _2228_ (.A0(net28),
    .A1(\wbs_o_buff[22] ),
    .S(_0679_),
    .X(_0682_));
 sky130_fd_sc_hd__clkbuf_1 _2229_ (.A(_0682_),
    .X(net130));
 sky130_fd_sc_hd__mux2_1 _2230_ (.A0(net29),
    .A1(\wbs_o_buff[23] ),
    .S(_0679_),
    .X(_0683_));
 sky130_fd_sc_hd__clkbuf_1 _2231_ (.A(_0683_),
    .X(net131));
 sky130_fd_sc_hd__mux2_1 _2232_ (.A0(net30),
    .A1(\wbs_o_buff[24] ),
    .S(_0679_),
    .X(_0684_));
 sky130_fd_sc_hd__clkbuf_1 _2233_ (.A(_0684_),
    .X(net132));
 sky130_fd_sc_hd__mux2_1 _2234_ (.A0(net31),
    .A1(\wbs_o_buff[25] ),
    .S(_0679_),
    .X(_0685_));
 sky130_fd_sc_hd__clkbuf_1 _2235_ (.A(_0685_),
    .X(net133));
 sky130_fd_sc_hd__mux2_1 _2236_ (.A0(net32),
    .A1(\wbs_o_buff[26] ),
    .S(_0679_),
    .X(_0686_));
 sky130_fd_sc_hd__clkbuf_1 _2237_ (.A(_0686_),
    .X(net134));
 sky130_fd_sc_hd__mux2_1 _2238_ (.A0(net33),
    .A1(\wbs_o_buff[27] ),
    .S(_0679_),
    .X(_0687_));
 sky130_fd_sc_hd__clkbuf_1 _2239_ (.A(_0687_),
    .X(net135));
 sky130_fd_sc_hd__mux2_1 _2240_ (.A0(net34),
    .A1(\wbs_o_buff[28] ),
    .S(_0679_),
    .X(_0688_));
 sky130_fd_sc_hd__clkbuf_1 _2241_ (.A(_0688_),
    .X(net136));
 sky130_fd_sc_hd__mux2_1 _2242_ (.A0(net35),
    .A1(\wbs_o_buff[29] ),
    .S(_0679_),
    .X(_0689_));
 sky130_fd_sc_hd__clkbuf_1 _2243_ (.A(_0689_),
    .X(net137));
 sky130_fd_sc_hd__mux2_1 _2244_ (.A0(net37),
    .A1(\wbs_o_buff[30] ),
    .S(net49),
    .X(_0690_));
 sky130_fd_sc_hd__clkbuf_1 _2245_ (.A(_0690_),
    .X(net139));
 sky130_fd_sc_hd__mux2_1 _2246_ (.A0(net38),
    .A1(\wbs_o_buff[31] ),
    .S(net49),
    .X(_0691_));
 sky130_fd_sc_hd__clkbuf_1 _2247_ (.A(_0691_),
    .X(net140));
 sky130_fd_sc_hd__mux2_1 _2248_ (.A0(net2),
    .A1(\K_override[0] ),
    .S(net148),
    .X(_0692_));
 sky130_fd_sc_hd__clkbuf_1 _2249_ (.A(_0692_),
    .X(\tms1x00.K_in[0] ));
 sky130_fd_sc_hd__mux2_1 _2250_ (.A0(net3),
    .A1(\K_override[1] ),
    .S(net148),
    .X(_0693_));
 sky130_fd_sc_hd__clkbuf_1 _2251_ (.A(_0693_),
    .X(\tms1x00.K_in[1] ));
 sky130_fd_sc_hd__mux2_1 _2252_ (.A0(net4),
    .A1(\K_override[2] ),
    .S(net148),
    .X(_0694_));
 sky130_fd_sc_hd__clkbuf_1 _2253_ (.A(_0694_),
    .X(\tms1x00.K_in[2] ));
 sky130_fd_sc_hd__mux2_1 _2254_ (.A0(net5),
    .A1(\K_override[3] ),
    .S(net148),
    .X(_0695_));
 sky130_fd_sc_hd__clkbuf_1 _2255_ (.A(_0695_),
    .X(\tms1x00.K_in[3] ));
 sky130_fd_sc_hd__clkinv_2 _2256_ (.A(net68),
    .Y(net114));
 sky130_fd_sc_hd__and3_1 _2257_ (.A(net49),
    .B(net114),
    .C(valid),
    .X(_0696_));
 sky130_fd_sc_hd__buf_4 _2258_ (.A(_0696_),
    .X(_0697_));
 sky130_fd_sc_hd__buf_2 _2259_ (.A(_0697_),
    .X(_0698_));
 sky130_fd_sc_hd__nor2_4 _2260_ (.A(net46),
    .B(_0697_),
    .Y(_0699_));
 sky130_fd_sc_hd__buf_2 _2261_ (.A(_0699_),
    .X(_0700_));
 sky130_fd_sc_hd__a22o_1 _2262_ (.A1(net69),
    .A2(_0698_),
    .B1(_0700_),
    .B2(\wbs_o_buff[0] ),
    .X(_0003_));
 sky130_fd_sc_hd__a22o_1 _2263_ (.A1(net70),
    .A2(_0698_),
    .B1(_0700_),
    .B2(\wbs_o_buff[1] ),
    .X(_0014_));
 sky130_fd_sc_hd__a22o_1 _2264_ (.A1(net71),
    .A2(_0698_),
    .B1(_0700_),
    .B2(\wbs_o_buff[2] ),
    .X(_0025_));
 sky130_fd_sc_hd__a22o_1 _2265_ (.A1(net72),
    .A2(_0698_),
    .B1(_0700_),
    .B2(\wbs_o_buff[3] ),
    .X(_0028_));
 sky130_fd_sc_hd__a22o_1 _2266_ (.A1(net73),
    .A2(_0698_),
    .B1(_0700_),
    .B2(\wbs_o_buff[4] ),
    .X(_0029_));
 sky130_fd_sc_hd__clkbuf_4 _2267_ (.A(net74),
    .X(_0701_));
 sky130_fd_sc_hd__a22o_1 _2268_ (.A1(_0701_),
    .A2(_0698_),
    .B1(_0700_),
    .B2(\wbs_o_buff[5] ),
    .X(_0030_));
 sky130_fd_sc_hd__a22o_1 _2269_ (.A1(net75),
    .A2(_0698_),
    .B1(_0700_),
    .B2(\wbs_o_buff[6] ),
    .X(_0031_));
 sky130_fd_sc_hd__a22o_1 _2270_ (.A1(net76),
    .A2(_0698_),
    .B1(_0700_),
    .B2(\wbs_o_buff[7] ),
    .X(_0032_));
 sky130_fd_sc_hd__a22o_1 _2271_ (.A1(net77),
    .A2(_0698_),
    .B1(_0700_),
    .B2(\wbs_o_buff[8] ),
    .X(_0033_));
 sky130_fd_sc_hd__a22o_1 _2272_ (.A1(net78),
    .A2(_0698_),
    .B1(_0700_),
    .B2(\wbs_o_buff[9] ),
    .X(_0034_));
 sky130_fd_sc_hd__clkbuf_4 _2273_ (.A(_0697_),
    .X(_0702_));
 sky130_fd_sc_hd__clkbuf_4 _2274_ (.A(_0699_),
    .X(_0703_));
 sky130_fd_sc_hd__a22o_1 _2275_ (.A1(net79),
    .A2(_0702_),
    .B1(_0703_),
    .B2(\wbs_o_buff[10] ),
    .X(_0004_));
 sky130_fd_sc_hd__a22o_1 _2276_ (.A1(net80),
    .A2(_0702_),
    .B1(_0703_),
    .B2(\wbs_o_buff[11] ),
    .X(_0005_));
 sky130_fd_sc_hd__a22o_1 _2277_ (.A1(net81),
    .A2(_0702_),
    .B1(_0703_),
    .B2(\wbs_o_buff[12] ),
    .X(_0006_));
 sky130_fd_sc_hd__a22o_1 _2278_ (.A1(net82),
    .A2(_0702_),
    .B1(_0703_),
    .B2(\wbs_o_buff[13] ),
    .X(_0007_));
 sky130_fd_sc_hd__a22o_1 _2279_ (.A1(net83),
    .A2(_0702_),
    .B1(_0703_),
    .B2(\wbs_o_buff[14] ),
    .X(_0008_));
 sky130_fd_sc_hd__a22o_1 _2280_ (.A1(net84),
    .A2(_0702_),
    .B1(_0703_),
    .B2(\wbs_o_buff[15] ),
    .X(_0009_));
 sky130_fd_sc_hd__a22o_1 _2281_ (.A1(net85),
    .A2(_0702_),
    .B1(_0703_),
    .B2(\wbs_o_buff[16] ),
    .X(_0010_));
 sky130_fd_sc_hd__a22o_1 _2282_ (.A1(net86),
    .A2(_0702_),
    .B1(_0703_),
    .B2(\wbs_o_buff[17] ),
    .X(_0011_));
 sky130_fd_sc_hd__a22o_1 _2283_ (.A1(net87),
    .A2(_0702_),
    .B1(_0703_),
    .B2(\wbs_o_buff[18] ),
    .X(_0012_));
 sky130_fd_sc_hd__a22o_1 _2284_ (.A1(net88),
    .A2(_0702_),
    .B1(_0703_),
    .B2(\wbs_o_buff[19] ),
    .X(_0013_));
 sky130_fd_sc_hd__buf_2 _2285_ (.A(_0699_),
    .X(_0704_));
 sky130_fd_sc_hd__a22o_1 _2286_ (.A1(net89),
    .A2(_0697_),
    .B1(_0704_),
    .B2(\wbs_o_buff[20] ),
    .X(_0015_));
 sky130_fd_sc_hd__a22o_1 _2287_ (.A1(net90),
    .A2(_0697_),
    .B1(_0704_),
    .B2(\wbs_o_buff[21] ),
    .X(_0016_));
 sky130_fd_sc_hd__a22o_1 _2288_ (.A1(net91),
    .A2(_0697_),
    .B1(_0704_),
    .B2(\wbs_o_buff[22] ),
    .X(_0017_));
 sky130_fd_sc_hd__a22o_1 _2289_ (.A1(net92),
    .A2(_0697_),
    .B1(_0704_),
    .B2(\wbs_o_buff[23] ),
    .X(_0018_));
 sky130_fd_sc_hd__and2_1 _2290_ (.A(\wbs_o_buff[24] ),
    .B(_0704_),
    .X(_0705_));
 sky130_fd_sc_hd__clkbuf_1 _2291_ (.A(_0705_),
    .X(_0019_));
 sky130_fd_sc_hd__and2_1 _2292_ (.A(\wbs_o_buff[25] ),
    .B(_0704_),
    .X(_0706_));
 sky130_fd_sc_hd__clkbuf_1 _2293_ (.A(_0706_),
    .X(_0020_));
 sky130_fd_sc_hd__and2_1 _2294_ (.A(\wbs_o_buff[26] ),
    .B(_0704_),
    .X(_0707_));
 sky130_fd_sc_hd__clkbuf_1 _2295_ (.A(_0707_),
    .X(_0021_));
 sky130_fd_sc_hd__and2_1 _2296_ (.A(\wbs_o_buff[27] ),
    .B(_0704_),
    .X(_0708_));
 sky130_fd_sc_hd__clkbuf_1 _2297_ (.A(_0708_),
    .X(_0022_));
 sky130_fd_sc_hd__and2_1 _2298_ (.A(\wbs_o_buff[28] ),
    .B(_0704_),
    .X(_0709_));
 sky130_fd_sc_hd__clkbuf_1 _2299_ (.A(_0709_),
    .X(_0023_));
 sky130_fd_sc_hd__and2_1 _2300_ (.A(\wbs_o_buff[29] ),
    .B(_0704_),
    .X(_0710_));
 sky130_fd_sc_hd__clkbuf_1 _2301_ (.A(_0710_),
    .X(_0024_));
 sky130_fd_sc_hd__and2_1 _2302_ (.A(\wbs_o_buff[30] ),
    .B(_0699_),
    .X(_0711_));
 sky130_fd_sc_hd__clkbuf_1 _2303_ (.A(_0711_),
    .X(_0026_));
 sky130_fd_sc_hd__and2_1 _2304_ (.A(\wbs_o_buff[31] ),
    .B(_0699_),
    .X(_0712_));
 sky130_fd_sc_hd__clkbuf_1 _2305_ (.A(_0712_),
    .X(_0027_));
 sky130_fd_sc_hd__inv_2 _2306_ (.A(net46),
    .Y(_0713_));
 sky130_fd_sc_hd__nand3_2 _2307_ (.A(net49),
    .B(net68),
    .C(valid),
    .Y(_0714_));
 sky130_fd_sc_hd__and3_2 _2308_ (.A(net49),
    .B(net68),
    .C(valid),
    .X(_0715_));
 sky130_fd_sc_hd__and2_1 _2309_ (.A(net59),
    .B(_0715_),
    .X(_0716_));
 sky130_fd_sc_hd__a32o_1 _2310_ (.A1(wb_rst_override),
    .A2(_0713_),
    .A3(_0714_),
    .B1(_0716_),
    .B2(net62),
    .X(_0001_));
 sky130_fd_sc_hd__a32o_1 _2311_ (.A1(\tms1x00.wb_step ),
    .A2(_0713_),
    .A3(_0714_),
    .B1(_0716_),
    .B2(net63),
    .X(_0002_));
 sky130_fd_sc_hd__a31o_1 _2312_ (.A1(_0713_),
    .A2(net148),
    .A3(_0714_),
    .B1(_0716_),
    .X(_0000_));
 sky130_fd_sc_hd__clkbuf_4 _2313_ (.A(\tms1x00.ram_addr_buff[0] ),
    .X(_0717_));
 sky130_fd_sc_hd__nor2_8 _2314_ (.A(wb_rst_override),
    .B(net46),
    .Y(_0718_));
 sky130_fd_sc_hd__inv_2 _2315_ (.A(net76),
    .Y(_0719_));
 sky130_fd_sc_hd__nor2_2 _2316_ (.A(_0719_),
    .B(net75),
    .Y(_0720_));
 sky130_fd_sc_hd__xnor2_2 _2317_ (.A(\tms1x00.wb_step ),
    .B(\tms1x00.wb_step_state ),
    .Y(_0721_));
 sky130_fd_sc_hd__nand2_1 _2318_ (.A(net148),
    .B(_0721_),
    .Y(_0722_));
 sky130_fd_sc_hd__and3b_1 _2319_ (.A_N(_0701_),
    .B(_0720_),
    .C(_0722_),
    .X(_0723_));
 sky130_fd_sc_hd__clkbuf_4 _2320_ (.A(_0723_),
    .X(_0724_));
 sky130_fd_sc_hd__nand2_2 _2321_ (.A(_0718_),
    .B(_0724_),
    .Y(_0725_));
 sky130_fd_sc_hd__buf_4 _2322_ (.A(_0725_),
    .X(_0726_));
 sky130_fd_sc_hd__mux2_1 _2323_ (.A0(\tms1x00.Y[0] ),
    .A1(_0717_),
    .S(_0726_),
    .X(_0727_));
 sky130_fd_sc_hd__clkbuf_1 _2324_ (.A(_0727_),
    .X(_0042_));
 sky130_fd_sc_hd__clkbuf_4 _2325_ (.A(\tms1x00.ram_addr_buff[1] ),
    .X(_0728_));
 sky130_fd_sc_hd__mux2_1 _2326_ (.A0(\tms1x00.Y[1] ),
    .A1(_0728_),
    .S(_0726_),
    .X(_0729_));
 sky130_fd_sc_hd__clkbuf_1 _2327_ (.A(_0729_),
    .X(_0043_));
 sky130_fd_sc_hd__buf_2 _2328_ (.A(\tms1x00.Y[2] ),
    .X(_0730_));
 sky130_fd_sc_hd__mux2_1 _2329_ (.A0(_0730_),
    .A1(\tms1x00.ram_addr_buff[2] ),
    .S(_0726_),
    .X(_0731_));
 sky130_fd_sc_hd__clkbuf_1 _2330_ (.A(_0731_),
    .X(_0044_));
 sky130_fd_sc_hd__buf_2 _2331_ (.A(\tms1x00.Y[3] ),
    .X(_0732_));
 sky130_fd_sc_hd__buf_2 _2332_ (.A(_0732_),
    .X(_0733_));
 sky130_fd_sc_hd__mux2_1 _2333_ (.A0(_0733_),
    .A1(\tms1x00.ram_addr_buff[3] ),
    .S(_0726_),
    .X(_0734_));
 sky130_fd_sc_hd__clkbuf_1 _2334_ (.A(_0734_),
    .X(_0045_));
 sky130_fd_sc_hd__mux2_1 _2335_ (.A0(\tms1x00.X[2] ),
    .A1(\tms1x00.ram_addr_buff[4] ),
    .S(_0726_),
    .X(_0735_));
 sky130_fd_sc_hd__clkbuf_1 _2336_ (.A(_0735_),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_1 _2337_ (.A0(\tms1x00.X[0] ),
    .A1(\tms1x00.ram_addr_buff[5] ),
    .S(_0726_),
    .X(_0736_));
 sky130_fd_sc_hd__clkbuf_1 _2338_ (.A(_0736_),
    .X(_0047_));
 sky130_fd_sc_hd__mux2_1 _2339_ (.A0(\tms1x00.X[1] ),
    .A1(\tms1x00.ram_addr_buff[6] ),
    .S(_0726_),
    .X(_0737_));
 sky130_fd_sc_hd__clkbuf_1 _2340_ (.A(_0737_),
    .X(_0048_));
 sky130_fd_sc_hd__clkinv_4 _2341_ (.A(_0718_),
    .Y(_0738_));
 sky130_fd_sc_hd__clkbuf_4 _2342_ (.A(_0738_),
    .X(net103));
 sky130_fd_sc_hd__nand2_1 _2343_ (.A(net48),
    .B(valid),
    .Y(net113));
 sky130_fd_sc_hd__clkinv_2 _2344_ (.A(\tms1x00.Y[2] ),
    .Y(_0739_));
 sky130_fd_sc_hd__nor2_1 _2345_ (.A(\tms1x00.Y[1] ),
    .B(\tms1x00.Y[0] ),
    .Y(_0740_));
 sky130_fd_sc_hd__nand2_1 _2346_ (.A(_0739_),
    .B(_0740_),
    .Y(_0741_));
 sky130_fd_sc_hd__buf_2 _2347_ (.A(\tms1x00.ins_in[0] ),
    .X(_0742_));
 sky130_fd_sc_hd__buf_2 _2348_ (.A(\tms1x00.ins_in[3] ),
    .X(_0743_));
 sky130_fd_sc_hd__nand2_1 _2349_ (.A(_0743_),
    .B(\tms1x00.ins_in[2] ),
    .Y(_0744_));
 sky130_fd_sc_hd__nand3b_1 _2350_ (.A_N(net76),
    .B(net75),
    .C(net74),
    .Y(_0745_));
 sky130_fd_sc_hd__a21o_2 _2351_ (.A1(net148),
    .A2(_0721_),
    .B1(_0745_),
    .X(_0746_));
 sky130_fd_sc_hd__clkbuf_4 _2352_ (.A(\tms1x00.ins_in[7] ),
    .X(_0747_));
 sky130_fd_sc_hd__clkbuf_4 _2353_ (.A(\tms1x00.ins_in[6] ),
    .X(_0748_));
 sky130_fd_sc_hd__or3_1 _2354_ (.A(_0747_),
    .B(_0748_),
    .C(\tms1x00.ins_in[5] ),
    .X(_0749_));
 sky130_fd_sc_hd__or2_1 _2355_ (.A(\tms1x00.ins_in[4] ),
    .B(_0749_),
    .X(_0750_));
 sky130_fd_sc_hd__or2_1 _2356_ (.A(_0746_),
    .B(_0750_),
    .X(_0751_));
 sky130_fd_sc_hd__or4_4 _2357_ (.A(\tms1x00.ins_in[1] ),
    .B(_0742_),
    .C(_0744_),
    .D(_0751_),
    .X(_0752_));
 sky130_fd_sc_hd__buf_2 _2358_ (.A(_0752_),
    .X(_0753_));
 sky130_fd_sc_hd__inv_2 _2359_ (.A(\tms1x00.Y[3] ),
    .Y(_0754_));
 sky130_fd_sc_hd__clkbuf_2 _2360_ (.A(_0754_),
    .X(_0755_));
 sky130_fd_sc_hd__and2_1 _2361_ (.A(_0739_),
    .B(_0740_),
    .X(_0756_));
 sky130_fd_sc_hd__or3b_1 _2362_ (.A(_0744_),
    .B(\tms1x00.ins_in[1] ),
    .C_N(_0742_),
    .X(_0757_));
 sky130_fd_sc_hd__inv_2 _2363_ (.A(_0749_),
    .Y(_0758_));
 sky130_fd_sc_hd__and2_1 _2364_ (.A(net148),
    .B(_0721_),
    .X(_0759_));
 sky130_fd_sc_hd__buf_2 _2365_ (.A(_0759_),
    .X(_0760_));
 sky130_fd_sc_hd__nor2_1 _2366_ (.A(_0760_),
    .B(_0745_),
    .Y(_0761_));
 sky130_fd_sc_hd__clkinv_2 _2367_ (.A(\tms1x00.ins_in[4] ),
    .Y(_0762_));
 sky130_fd_sc_hd__and4b_2 _2368_ (.A_N(_0757_),
    .B(_0758_),
    .C(_0761_),
    .D(_0762_),
    .X(_0763_));
 sky130_fd_sc_hd__buf_2 _2369_ (.A(_0763_),
    .X(_0764_));
 sky130_fd_sc_hd__a31o_1 _2370_ (.A1(_0755_),
    .A2(_0756_),
    .A3(_0764_),
    .B1(net77),
    .X(_0765_));
 sky130_fd_sc_hd__clkbuf_4 _2371_ (.A(_0718_),
    .X(_0766_));
 sky130_fd_sc_hd__o311a_1 _2372_ (.A1(_0733_),
    .A2(_0741_),
    .A3(_0753_),
    .B1(_0765_),
    .C1(_0766_),
    .X(_0049_));
 sky130_fd_sc_hd__a22o_1 _2373_ (.A1(chip_sel_override),
    .A2(_0714_),
    .B1(_0716_),
    .B2(net64),
    .X(_0050_));
 sky130_fd_sc_hd__or4b_1 _2374_ (.A(net76),
    .B(net74),
    .C(\tms1x00.ins_in[1] ),
    .D_N(net75),
    .X(_0767_));
 sky130_fd_sc_hd__inv_2 _2375_ (.A(\tms1x00.ins_in[2] ),
    .Y(_0768_));
 sky130_fd_sc_hd__and4b_1 _2376_ (.A_N(\tms1x00.ins_in[5] ),
    .B(\tms1x00.ins_in[4] ),
    .C(\tms1x00.ins_in[7] ),
    .D(\tms1x00.ins_in[6] ),
    .X(_0769_));
 sky130_fd_sc_hd__or3b_1 _2377_ (.A(\tms1x00.ins_in[3] ),
    .B(_0768_),
    .C_N(_0769_),
    .X(_0770_));
 sky130_fd_sc_hd__or4_2 _2378_ (.A(_0738_),
    .B(_0760_),
    .C(_0767_),
    .D(_0770_),
    .X(_0771_));
 sky130_fd_sc_hd__or2_1 _2379_ (.A(_0747_),
    .B(_0748_),
    .X(_0772_));
 sky130_fd_sc_hd__clkinv_2 _2380_ (.A(_0040_),
    .Y(_0773_));
 sky130_fd_sc_hd__inv_2 _2381_ (.A(_0038_),
    .Y(_0774_));
 sky130_fd_sc_hd__clkbuf_4 _2382_ (.A(_0774_),
    .X(_0775_));
 sky130_fd_sc_hd__clkbuf_4 _2383_ (.A(_0775_),
    .X(_0776_));
 sky130_fd_sc_hd__buf_6 _2384_ (.A(_0035_),
    .X(_0777_));
 sky130_fd_sc_hd__buf_4 _2385_ (.A(_0777_),
    .X(_0778_));
 sky130_fd_sc_hd__clkbuf_8 _2386_ (.A(_0036_),
    .X(_0779_));
 sky130_fd_sc_hd__buf_6 _2387_ (.A(_0779_),
    .X(_0780_));
 sky130_fd_sc_hd__mux4_1 _2388_ (.A0(\tms1x00.RAM[80][0] ),
    .A1(\tms1x00.RAM[81][0] ),
    .A2(\tms1x00.RAM[82][0] ),
    .A3(\tms1x00.RAM[83][0] ),
    .S0(_0778_),
    .S1(_0780_),
    .X(_0781_));
 sky130_fd_sc_hd__mux4_1 _2389_ (.A0(\tms1x00.RAM[84][0] ),
    .A1(\tms1x00.RAM[85][0] ),
    .A2(\tms1x00.RAM[86][0] ),
    .A3(\tms1x00.RAM[87][0] ),
    .S0(_0778_),
    .S1(_0780_),
    .X(_0782_));
 sky130_fd_sc_hd__clkbuf_4 _2390_ (.A(_0037_),
    .X(_0783_));
 sky130_fd_sc_hd__mux2_1 _2391_ (.A0(_0781_),
    .A1(_0782_),
    .S(_0783_),
    .X(_0784_));
 sky130_fd_sc_hd__inv_2 _2392_ (.A(_0036_),
    .Y(_0785_));
 sky130_fd_sc_hd__clkbuf_4 _2393_ (.A(_0785_),
    .X(_0786_));
 sky130_fd_sc_hd__buf_4 _2394_ (.A(_0786_),
    .X(_0787_));
 sky130_fd_sc_hd__buf_6 _2395_ (.A(_0777_),
    .X(_0788_));
 sky130_fd_sc_hd__buf_4 _2396_ (.A(_0788_),
    .X(_0789_));
 sky130_fd_sc_hd__mux2_1 _2397_ (.A0(\tms1x00.RAM[92][0] ),
    .A1(\tms1x00.RAM[93][0] ),
    .S(_0789_),
    .X(_0790_));
 sky130_fd_sc_hd__buf_6 _2398_ (.A(_0780_),
    .X(_0791_));
 sky130_fd_sc_hd__mux2_1 _2399_ (.A0(\tms1x00.RAM[94][0] ),
    .A1(\tms1x00.RAM[95][0] ),
    .S(_0788_),
    .X(_0792_));
 sky130_fd_sc_hd__inv_2 _2400_ (.A(_0037_),
    .Y(_0793_));
 sky130_fd_sc_hd__clkbuf_4 _2401_ (.A(_0793_),
    .X(_0794_));
 sky130_fd_sc_hd__a21o_1 _2402_ (.A1(_0791_),
    .A2(_0792_),
    .B1(_0794_),
    .X(_0795_));
 sky130_fd_sc_hd__a21o_1 _2403_ (.A1(_0787_),
    .A2(_0790_),
    .B1(_0795_),
    .X(_0796_));
 sky130_fd_sc_hd__buf_2 _2404_ (.A(_0037_),
    .X(_0797_));
 sky130_fd_sc_hd__clkbuf_4 _2405_ (.A(_0797_),
    .X(_0798_));
 sky130_fd_sc_hd__clkbuf_16 _2406_ (.A(_0777_),
    .X(_0799_));
 sky130_fd_sc_hd__buf_6 _2407_ (.A(_0779_),
    .X(_0800_));
 sky130_fd_sc_hd__mux4_1 _2408_ (.A0(\tms1x00.RAM[88][0] ),
    .A1(\tms1x00.RAM[89][0] ),
    .A2(\tms1x00.RAM[90][0] ),
    .A3(\tms1x00.RAM[91][0] ),
    .S0(_0799_),
    .S1(_0800_),
    .X(_0801_));
 sky130_fd_sc_hd__clkbuf_4 _2409_ (.A(_0038_),
    .X(_0802_));
 sky130_fd_sc_hd__o21a_1 _2410_ (.A1(_0798_),
    .A2(_0801_),
    .B1(_0802_),
    .X(_0803_));
 sky130_fd_sc_hd__inv_2 _2411_ (.A(_0039_),
    .Y(_0804_));
 sky130_fd_sc_hd__a221o_1 _2412_ (.A1(_0776_),
    .A2(_0784_),
    .B1(_0796_),
    .B2(_0803_),
    .C1(_0804_),
    .X(_0805_));
 sky130_fd_sc_hd__clkbuf_4 _2413_ (.A(_0038_),
    .X(_0806_));
 sky130_fd_sc_hd__clkbuf_4 _2414_ (.A(_0797_),
    .X(_0807_));
 sky130_fd_sc_hd__buf_8 _2415_ (.A(_0777_),
    .X(_0808_));
 sky130_fd_sc_hd__mux4_1 _2416_ (.A0(\tms1x00.RAM[72][0] ),
    .A1(\tms1x00.RAM[73][0] ),
    .A2(\tms1x00.RAM[74][0] ),
    .A3(\tms1x00.RAM[75][0] ),
    .S0(_0808_),
    .S1(_0780_),
    .X(_0809_));
 sky130_fd_sc_hd__or2_1 _2417_ (.A(_0807_),
    .B(_0809_),
    .X(_0810_));
 sky130_fd_sc_hd__or2b_1 _2418_ (.A(\tms1x00.RAM[79][0] ),
    .B_N(_0789_),
    .X(_0811_));
 sky130_fd_sc_hd__buf_6 _2419_ (.A(_0036_),
    .X(_0812_));
 sky130_fd_sc_hd__buf_6 _2420_ (.A(_0812_),
    .X(_0813_));
 sky130_fd_sc_hd__o21a_1 _2421_ (.A1(_0789_),
    .A2(\tms1x00.RAM[78][0] ),
    .B1(_0813_),
    .X(_0814_));
 sky130_fd_sc_hd__buf_8 _2422_ (.A(_0035_),
    .X(_0815_));
 sky130_fd_sc_hd__buf_6 _2423_ (.A(_0815_),
    .X(_0816_));
 sky130_fd_sc_hd__mux2_1 _2424_ (.A0(\tms1x00.RAM[76][0] ),
    .A1(\tms1x00.RAM[77][0] ),
    .S(_0816_),
    .X(_0817_));
 sky130_fd_sc_hd__clkbuf_4 _2425_ (.A(_0785_),
    .X(_0818_));
 sky130_fd_sc_hd__clkbuf_4 _2426_ (.A(_0793_),
    .X(_0819_));
 sky130_fd_sc_hd__a221o_1 _2427_ (.A1(_0811_),
    .A2(_0814_),
    .B1(_0817_),
    .B2(_0818_),
    .C1(_0819_),
    .X(_0820_));
 sky130_fd_sc_hd__clkbuf_4 _2428_ (.A(_0039_),
    .X(_0821_));
 sky130_fd_sc_hd__buf_6 _2429_ (.A(_0812_),
    .X(_0822_));
 sky130_fd_sc_hd__buf_6 _2430_ (.A(_0035_),
    .X(_0823_));
 sky130_fd_sc_hd__mux2_1 _2431_ (.A0(\tms1x00.RAM[70][0] ),
    .A1(\tms1x00.RAM[71][0] ),
    .S(_0823_),
    .X(_0824_));
 sky130_fd_sc_hd__and2_1 _2432_ (.A(_0822_),
    .B(_0824_),
    .X(_0825_));
 sky130_fd_sc_hd__buf_6 _2433_ (.A(_0035_),
    .X(_0826_));
 sky130_fd_sc_hd__mux2_1 _2434_ (.A0(\tms1x00.RAM[68][0] ),
    .A1(\tms1x00.RAM[69][0] ),
    .S(_0826_),
    .X(_0827_));
 sky130_fd_sc_hd__clkbuf_4 _2435_ (.A(_0793_),
    .X(_0828_));
 sky130_fd_sc_hd__a21o_1 _2436_ (.A1(_0786_),
    .A2(_0827_),
    .B1(_0828_),
    .X(_0829_));
 sky130_fd_sc_hd__buf_6 _2437_ (.A(_0777_),
    .X(_0830_));
 sky130_fd_sc_hd__buf_6 _2438_ (.A(_0779_),
    .X(_0831_));
 sky130_fd_sc_hd__mux4_1 _2439_ (.A0(\tms1x00.RAM[64][0] ),
    .A1(\tms1x00.RAM[65][0] ),
    .A2(\tms1x00.RAM[66][0] ),
    .A3(\tms1x00.RAM[67][0] ),
    .S0(_0830_),
    .S1(_0831_),
    .X(_0832_));
 sky130_fd_sc_hd__o221a_1 _2440_ (.A1(_0825_),
    .A2(_0829_),
    .B1(_0832_),
    .B2(_0807_),
    .C1(_0775_),
    .X(_0833_));
 sky130_fd_sc_hd__a311o_1 _2441_ (.A1(_0806_),
    .A2(_0810_),
    .A3(_0820_),
    .B1(_0821_),
    .C1(_0833_),
    .X(_0834_));
 sky130_fd_sc_hd__inv_2 _2442_ (.A(_0041_),
    .Y(_0835_));
 sky130_fd_sc_hd__mux4_1 _2443_ (.A0(\tms1x00.RAM[108][0] ),
    .A1(\tms1x00.RAM[109][0] ),
    .A2(\tms1x00.RAM[110][0] ),
    .A3(\tms1x00.RAM[111][0] ),
    .S0(_0799_),
    .S1(_0800_),
    .X(_0836_));
 sky130_fd_sc_hd__mux4_1 _2444_ (.A0(\tms1x00.RAM[104][0] ),
    .A1(\tms1x00.RAM[105][0] ),
    .A2(\tms1x00.RAM[106][0] ),
    .A3(\tms1x00.RAM[107][0] ),
    .S0(_0777_),
    .S1(_0779_),
    .X(_0837_));
 sky130_fd_sc_hd__or2_1 _2445_ (.A(_0797_),
    .B(_0837_),
    .X(_0838_));
 sky130_fd_sc_hd__o211a_1 _2446_ (.A1(_0819_),
    .A2(_0836_),
    .B1(_0838_),
    .C1(_0802_),
    .X(_0839_));
 sky130_fd_sc_hd__buf_8 _2447_ (.A(_0815_),
    .X(_0840_));
 sky130_fd_sc_hd__mux4_2 _2448_ (.A0(\tms1x00.RAM[96][0] ),
    .A1(\tms1x00.RAM[97][0] ),
    .A2(\tms1x00.RAM[98][0] ),
    .A3(\tms1x00.RAM[99][0] ),
    .S0(_0840_),
    .S1(_0813_),
    .X(_0841_));
 sky130_fd_sc_hd__mux4_1 _2449_ (.A0(\tms1x00.RAM[100][0] ),
    .A1(\tms1x00.RAM[101][0] ),
    .A2(\tms1x00.RAM[102][0] ),
    .A3(\tms1x00.RAM[103][0] ),
    .S0(_0815_),
    .S1(_0779_),
    .X(_0842_));
 sky130_fd_sc_hd__or2_1 _2450_ (.A(_0828_),
    .B(_0842_),
    .X(_0843_));
 sky130_fd_sc_hd__o211a_1 _2451_ (.A1(_0798_),
    .A2(_0841_),
    .B1(_0843_),
    .C1(_0775_),
    .X(_0844_));
 sky130_fd_sc_hd__mux4_1 _2452_ (.A0(\tms1x00.RAM[120][0] ),
    .A1(\tms1x00.RAM[121][0] ),
    .A2(\tms1x00.RAM[122][0] ),
    .A3(\tms1x00.RAM[123][0] ),
    .S0(_0815_),
    .S1(_0812_),
    .X(_0845_));
 sky130_fd_sc_hd__or2_1 _2453_ (.A(_0797_),
    .B(_0845_),
    .X(_0846_));
 sky130_fd_sc_hd__mux4_1 _2454_ (.A0(\tms1x00.RAM[124][0] ),
    .A1(\tms1x00.RAM[125][0] ),
    .A2(\tms1x00.RAM[126][0] ),
    .A3(\tms1x00.RAM[127][0] ),
    .S0(_0815_),
    .S1(_0812_),
    .X(_0847_));
 sky130_fd_sc_hd__o21a_1 _2455_ (.A1(_0794_),
    .A2(_0847_),
    .B1(_0038_),
    .X(_0848_));
 sky130_fd_sc_hd__or2b_1 _2456_ (.A(\tms1x00.RAM[119][0] ),
    .B_N(_0808_),
    .X(_0849_));
 sky130_fd_sc_hd__buf_6 _2457_ (.A(_0779_),
    .X(_0850_));
 sky130_fd_sc_hd__o21a_1 _2458_ (.A1(_0808_),
    .A2(\tms1x00.RAM[118][0] ),
    .B1(_0850_),
    .X(_0851_));
 sky130_fd_sc_hd__mux2_1 _2459_ (.A0(\tms1x00.RAM[116][0] ),
    .A1(\tms1x00.RAM[117][0] ),
    .S(_0788_),
    .X(_0852_));
 sky130_fd_sc_hd__a221o_1 _2460_ (.A1(_0849_),
    .A2(_0851_),
    .B1(_0852_),
    .B2(_0786_),
    .C1(_0828_),
    .X(_0853_));
 sky130_fd_sc_hd__mux4_2 _2461_ (.A0(\tms1x00.RAM[112][0] ),
    .A1(\tms1x00.RAM[113][0] ),
    .A2(\tms1x00.RAM[114][0] ),
    .A3(\tms1x00.RAM[115][0] ),
    .S0(_0815_),
    .S1(_0812_),
    .X(_0854_));
 sky130_fd_sc_hd__o21a_1 _2462_ (.A1(_0797_),
    .A2(_0854_),
    .B1(_0774_),
    .X(_0855_));
 sky130_fd_sc_hd__a221o_1 _2463_ (.A1(_0846_),
    .A2(_0848_),
    .B1(_0853_),
    .B2(_0855_),
    .C1(_0804_),
    .X(_0856_));
 sky130_fd_sc_hd__o311a_1 _2464_ (.A1(_0821_),
    .A2(_0839_),
    .A3(_0844_),
    .B1(_0856_),
    .C1(_0040_),
    .X(_0857_));
 sky130_fd_sc_hd__a311o_2 _2465_ (.A1(_0773_),
    .A2(_0805_),
    .A3(_0834_),
    .B1(_0835_),
    .C1(_0857_),
    .X(_0858_));
 sky130_fd_sc_hd__mux4_1 _2466_ (.A0(\tms1x00.RAM[16][0] ),
    .A1(\tms1x00.RAM[17][0] ),
    .A2(\tms1x00.RAM[18][0] ),
    .A3(\tms1x00.RAM[19][0] ),
    .S0(_0830_),
    .S1(_0831_),
    .X(_0859_));
 sky130_fd_sc_hd__mux4_2 _2467_ (.A0(\tms1x00.RAM[20][0] ),
    .A1(\tms1x00.RAM[21][0] ),
    .A2(\tms1x00.RAM[22][0] ),
    .A3(\tms1x00.RAM[23][0] ),
    .S0(_0830_),
    .S1(_0831_),
    .X(_0860_));
 sky130_fd_sc_hd__mux2_1 _2468_ (.A0(_0859_),
    .A1(_0860_),
    .S(_0783_),
    .X(_0861_));
 sky130_fd_sc_hd__mux2_1 _2469_ (.A0(\tms1x00.RAM[30][0] ),
    .A1(\tms1x00.RAM[31][0] ),
    .S(_0823_),
    .X(_0862_));
 sky130_fd_sc_hd__and2_1 _2470_ (.A(_0822_),
    .B(_0862_),
    .X(_0863_));
 sky130_fd_sc_hd__mux2_1 _2471_ (.A0(\tms1x00.RAM[28][0] ),
    .A1(\tms1x00.RAM[29][0] ),
    .S(_0826_),
    .X(_0864_));
 sky130_fd_sc_hd__a21o_1 _2472_ (.A1(_0786_),
    .A2(_0864_),
    .B1(_0828_),
    .X(_0865_));
 sky130_fd_sc_hd__mux4_2 _2473_ (.A0(\tms1x00.RAM[24][0] ),
    .A1(\tms1x00.RAM[25][0] ),
    .A2(\tms1x00.RAM[26][0] ),
    .A3(\tms1x00.RAM[27][0] ),
    .S0(_0830_),
    .S1(_0800_),
    .X(_0866_));
 sky130_fd_sc_hd__o221a_1 _2474_ (.A1(_0863_),
    .A2(_0865_),
    .B1(_0866_),
    .B2(_0798_),
    .C1(_0802_),
    .X(_0867_));
 sky130_fd_sc_hd__a211o_1 _2475_ (.A1(_0776_),
    .A2(_0861_),
    .B1(_0867_),
    .C1(_0804_),
    .X(_0868_));
 sky130_fd_sc_hd__mux4_1 _2476_ (.A0(\tms1x00.RAM[8][0] ),
    .A1(\tms1x00.RAM[9][0] ),
    .A2(\tms1x00.RAM[10][0] ),
    .A3(\tms1x00.RAM[11][0] ),
    .S0(_0808_),
    .S1(_0780_),
    .X(_0869_));
 sky130_fd_sc_hd__or2_1 _2477_ (.A(_0807_),
    .B(_0869_),
    .X(_0870_));
 sky130_fd_sc_hd__or2b_1 _2478_ (.A(\tms1x00.RAM[15][0] ),
    .B_N(_0789_),
    .X(_0871_));
 sky130_fd_sc_hd__o21a_1 _2479_ (.A1(_0789_),
    .A2(\tms1x00.RAM[14][0] ),
    .B1(_0813_),
    .X(_0872_));
 sky130_fd_sc_hd__buf_6 _2480_ (.A(_0815_),
    .X(_0873_));
 sky130_fd_sc_hd__mux2_1 _2481_ (.A0(\tms1x00.RAM[12][0] ),
    .A1(\tms1x00.RAM[13][0] ),
    .S(_0873_),
    .X(_0874_));
 sky130_fd_sc_hd__a221o_1 _2482_ (.A1(_0871_),
    .A2(_0872_),
    .B1(_0874_),
    .B2(_0818_),
    .C1(_0819_),
    .X(_0875_));
 sky130_fd_sc_hd__mux2_1 _2483_ (.A0(\tms1x00.RAM[6][0] ),
    .A1(\tms1x00.RAM[7][0] ),
    .S(_0823_),
    .X(_0876_));
 sky130_fd_sc_hd__and2_1 _2484_ (.A(_0822_),
    .B(_0876_),
    .X(_0877_));
 sky130_fd_sc_hd__mux2_1 _2485_ (.A0(\tms1x00.RAM[4][0] ),
    .A1(\tms1x00.RAM[5][0] ),
    .S(_0826_),
    .X(_0878_));
 sky130_fd_sc_hd__a21o_1 _2486_ (.A1(_0786_),
    .A2(_0878_),
    .B1(_0828_),
    .X(_0879_));
 sky130_fd_sc_hd__mux4_1 _2487_ (.A0(\tms1x00.RAM[0][0] ),
    .A1(\tms1x00.RAM[1][0] ),
    .A2(\tms1x00.RAM[2][0] ),
    .A3(\tms1x00.RAM[3][0] ),
    .S0(_0830_),
    .S1(_0831_),
    .X(_0880_));
 sky130_fd_sc_hd__o221a_1 _2488_ (.A1(_0877_),
    .A2(_0879_),
    .B1(_0880_),
    .B2(_0807_),
    .C1(_0775_),
    .X(_0881_));
 sky130_fd_sc_hd__a311o_1 _2489_ (.A1(_0806_),
    .A2(_0870_),
    .A3(_0875_),
    .B1(_0039_),
    .C1(_0881_),
    .X(_0882_));
 sky130_fd_sc_hd__mux4_2 _2490_ (.A0(\tms1x00.RAM[44][0] ),
    .A1(\tms1x00.RAM[45][0] ),
    .A2(\tms1x00.RAM[46][0] ),
    .A3(\tms1x00.RAM[47][0] ),
    .S0(_0808_),
    .S1(_0831_),
    .X(_0883_));
 sky130_fd_sc_hd__mux4_1 _2491_ (.A0(\tms1x00.RAM[40][0] ),
    .A1(\tms1x00.RAM[41][0] ),
    .A2(\tms1x00.RAM[42][0] ),
    .A3(\tms1x00.RAM[43][0] ),
    .S0(_0777_),
    .S1(_0779_),
    .X(_0884_));
 sky130_fd_sc_hd__or2_1 _2492_ (.A(_0797_),
    .B(_0884_),
    .X(_0885_));
 sky130_fd_sc_hd__o211a_1 _2493_ (.A1(_0819_),
    .A2(_0883_),
    .B1(_0885_),
    .C1(_0802_),
    .X(_0886_));
 sky130_fd_sc_hd__mux4_2 _2494_ (.A0(\tms1x00.RAM[32][0] ),
    .A1(\tms1x00.RAM[33][0] ),
    .A2(\tms1x00.RAM[34][0] ),
    .A3(\tms1x00.RAM[35][0] ),
    .S0(_0799_),
    .S1(_0800_),
    .X(_0887_));
 sky130_fd_sc_hd__mux4_1 _2495_ (.A0(\tms1x00.RAM[36][0] ),
    .A1(\tms1x00.RAM[37][0] ),
    .A2(\tms1x00.RAM[38][0] ),
    .A3(\tms1x00.RAM[39][0] ),
    .S0(_0777_),
    .S1(_0779_),
    .X(_0888_));
 sky130_fd_sc_hd__or2_1 _2496_ (.A(_0828_),
    .B(_0888_),
    .X(_0889_));
 sky130_fd_sc_hd__o211a_1 _2497_ (.A1(_0798_),
    .A2(_0887_),
    .B1(_0889_),
    .C1(_0775_),
    .X(_0890_));
 sky130_fd_sc_hd__mux4_1 _2498_ (.A0(\tms1x00.RAM[56][0] ),
    .A1(\tms1x00.RAM[57][0] ),
    .A2(\tms1x00.RAM[58][0] ),
    .A3(\tms1x00.RAM[59][0] ),
    .S0(_0777_),
    .S1(_0779_),
    .X(_0891_));
 sky130_fd_sc_hd__or2_1 _2499_ (.A(_0797_),
    .B(_0891_),
    .X(_0892_));
 sky130_fd_sc_hd__mux4_1 _2500_ (.A0(\tms1x00.RAM[60][0] ),
    .A1(\tms1x00.RAM[61][0] ),
    .A2(\tms1x00.RAM[62][0] ),
    .A3(\tms1x00.RAM[63][0] ),
    .S0(_0777_),
    .S1(_0779_),
    .X(_0893_));
 sky130_fd_sc_hd__o21a_1 _2501_ (.A1(_0828_),
    .A2(_0893_),
    .B1(_0038_),
    .X(_0894_));
 sky130_fd_sc_hd__or2b_1 _2502_ (.A(\tms1x00.RAM[55][0] ),
    .B_N(_0778_),
    .X(_0895_));
 sky130_fd_sc_hd__o21a_1 _2503_ (.A1(_0778_),
    .A2(\tms1x00.RAM[54][0] ),
    .B1(_0812_),
    .X(_0896_));
 sky130_fd_sc_hd__mux2_1 _2504_ (.A0(\tms1x00.RAM[52][0] ),
    .A1(\tms1x00.RAM[53][0] ),
    .S(_0826_),
    .X(_0897_));
 sky130_fd_sc_hd__a221o_1 _2505_ (.A1(_0895_),
    .A2(_0896_),
    .B1(_0897_),
    .B2(_0785_),
    .C1(_0828_),
    .X(_0898_));
 sky130_fd_sc_hd__mux4_1 _2506_ (.A0(\tms1x00.RAM[48][0] ),
    .A1(\tms1x00.RAM[49][0] ),
    .A2(\tms1x00.RAM[50][0] ),
    .A3(\tms1x00.RAM[51][0] ),
    .S0(_0815_),
    .S1(_0812_),
    .X(_0899_));
 sky130_fd_sc_hd__o21a_1 _2507_ (.A1(_0797_),
    .A2(_0899_),
    .B1(_0774_),
    .X(_0900_));
 sky130_fd_sc_hd__a221o_1 _2508_ (.A1(_0892_),
    .A2(_0894_),
    .B1(_0898_),
    .B2(_0900_),
    .C1(_0804_),
    .X(_0901_));
 sky130_fd_sc_hd__o311a_1 _2509_ (.A1(_0039_),
    .A2(_0886_),
    .A3(_0890_),
    .B1(_0901_),
    .C1(_0040_),
    .X(_0902_));
 sky130_fd_sc_hd__a311o_1 _2510_ (.A1(_0773_),
    .A2(_0868_),
    .A3(_0882_),
    .B1(_0902_),
    .C1(_0041_),
    .X(_0903_));
 sky130_fd_sc_hd__or4b_1 _2511_ (.A(_0747_),
    .B(_0762_),
    .C(_0748_),
    .D_N(\tms1x00.ins_in[5] ),
    .X(_0904_));
 sky130_fd_sc_hd__or4_1 _2512_ (.A(\tms1x00.ins_in[3] ),
    .B(_0738_),
    .C(_0746_),
    .D(_0904_),
    .X(_0905_));
 sky130_fd_sc_hd__nor2_1 _2513_ (.A(\tms1x00.ins_in[2] ),
    .B(_0905_),
    .Y(_0906_));
 sky130_fd_sc_hd__a31o_1 _2514_ (.A1(_0772_),
    .A2(_0858_),
    .A3(_0903_),
    .B1(_0906_),
    .X(_0907_));
 sky130_fd_sc_hd__nor2_1 _2515_ (.A(\tms1x00.ins_in[1] ),
    .B(_0742_),
    .Y(_0908_));
 sky130_fd_sc_hd__and2b_1 _2516_ (.A_N(_0771_),
    .B(_0908_),
    .X(_0909_));
 sky130_fd_sc_hd__a22o_1 _2517_ (.A1(_0771_),
    .A2(_0907_),
    .B1(_0909_),
    .B2(\tms1x00.A[0] ),
    .X(_0910_));
 sky130_fd_sc_hd__buf_4 _2518_ (.A(_0910_),
    .X(_0911_));
 sky130_fd_sc_hd__clkbuf_4 _2519_ (.A(_0911_),
    .X(_0912_));
 sky130_fd_sc_hd__nand3b_4 _2520_ (.A_N(\tms1x00.ram_addr_buff[4] ),
    .B(\tms1x00.ram_addr_buff[5] ),
    .C(\tms1x00.ram_addr_buff[6] ),
    .Y(_0913_));
 sky130_fd_sc_hd__clkbuf_8 _2521_ (.A(_0913_),
    .X(_0914_));
 sky130_fd_sc_hd__and2_1 _2522_ (.A(_0905_),
    .B(_0771_),
    .X(_0915_));
 sky130_fd_sc_hd__and3b_2 _2523_ (.A_N(_0915_),
    .B(\tms1x00.ram_addr_buff[3] ),
    .C(\tms1x00.ram_addr_buff[2] ),
    .X(_0916_));
 sky130_fd_sc_hd__nand3b_4 _2524_ (.A_N(_0728_),
    .B(_0916_),
    .C(_0717_),
    .Y(_0917_));
 sky130_fd_sc_hd__or2_2 _2525_ (.A(_0914_),
    .B(_0917_),
    .X(_0918_));
 sky130_fd_sc_hd__mux2_1 _2526_ (.A0(_0912_),
    .A1(\tms1x00.RAM[109][0] ),
    .S(_0918_),
    .X(_0919_));
 sky130_fd_sc_hd__clkbuf_1 _2527_ (.A(_0919_),
    .X(_0051_));
 sky130_fd_sc_hd__clkbuf_4 _2528_ (.A(_0804_),
    .X(_0920_));
 sky130_fd_sc_hd__clkbuf_4 _2529_ (.A(_0797_),
    .X(_0921_));
 sky130_fd_sc_hd__clkbuf_4 _2530_ (.A(_0921_),
    .X(_0922_));
 sky130_fd_sc_hd__buf_6 _2531_ (.A(_0826_),
    .X(_0923_));
 sky130_fd_sc_hd__buf_6 _2532_ (.A(_0923_),
    .X(_0924_));
 sky130_fd_sc_hd__mux2_1 _2533_ (.A0(\tms1x00.RAM[68][1] ),
    .A1(\tms1x00.RAM[69][1] ),
    .S(_0924_),
    .X(_0925_));
 sky130_fd_sc_hd__nand2_1 _2534_ (.A(_0787_),
    .B(_0925_),
    .Y(_0926_));
 sky130_fd_sc_hd__buf_4 _2535_ (.A(_0850_),
    .X(_0927_));
 sky130_fd_sc_hd__buf_4 _2536_ (.A(_0927_),
    .X(_0928_));
 sky130_fd_sc_hd__mux2_1 _2537_ (.A0(\tms1x00.RAM[70][1] ),
    .A1(\tms1x00.RAM[71][1] ),
    .S(_0924_),
    .X(_0929_));
 sky130_fd_sc_hd__nand2_1 _2538_ (.A(_0928_),
    .B(_0929_),
    .Y(_0930_));
 sky130_fd_sc_hd__buf_6 _2539_ (.A(_0840_),
    .X(_0931_));
 sky130_fd_sc_hd__clkbuf_8 _2540_ (.A(_0822_),
    .X(_0932_));
 sky130_fd_sc_hd__mux4_1 _2541_ (.A0(\tms1x00.RAM[64][1] ),
    .A1(\tms1x00.RAM[65][1] ),
    .A2(\tms1x00.RAM[66][1] ),
    .A3(\tms1x00.RAM[67][1] ),
    .S0(_0931_),
    .S1(_0932_),
    .X(_0933_));
 sky130_fd_sc_hd__o21ai_1 _2542_ (.A1(_0922_),
    .A2(_0933_),
    .B1(_0776_),
    .Y(_0934_));
 sky130_fd_sc_hd__a31o_1 _2543_ (.A1(_0922_),
    .A2(_0926_),
    .A3(_0930_),
    .B1(_0934_),
    .X(_0935_));
 sky130_fd_sc_hd__mux4_1 _2544_ (.A0(\tms1x00.RAM[72][1] ),
    .A1(\tms1x00.RAM[73][1] ),
    .A2(\tms1x00.RAM[74][1] ),
    .A3(\tms1x00.RAM[75][1] ),
    .S0(_0924_),
    .S1(_0928_),
    .X(_0936_));
 sky130_fd_sc_hd__or2b_1 _2545_ (.A(\tms1x00.RAM[79][1] ),
    .B_N(_0924_),
    .X(_0937_));
 sky130_fd_sc_hd__o21a_1 _2546_ (.A1(_0924_),
    .A2(\tms1x00.RAM[78][1] ),
    .B1(_0932_),
    .X(_0938_));
 sky130_fd_sc_hd__mux2_1 _2547_ (.A0(\tms1x00.RAM[76][1] ),
    .A1(\tms1x00.RAM[77][1] ),
    .S(_0924_),
    .X(_0939_));
 sky130_fd_sc_hd__clkbuf_4 _2548_ (.A(_0819_),
    .X(_0940_));
 sky130_fd_sc_hd__a221o_1 _2549_ (.A1(_0937_),
    .A2(_0938_),
    .B1(_0939_),
    .B2(_0787_),
    .C1(_0940_),
    .X(_0941_));
 sky130_fd_sc_hd__clkbuf_4 _2550_ (.A(_0802_),
    .X(_0942_));
 sky130_fd_sc_hd__o211ai_1 _2551_ (.A1(_0922_),
    .A2(_0936_),
    .B1(_0941_),
    .C1(_0942_),
    .Y(_0943_));
 sky130_fd_sc_hd__clkbuf_4 _2552_ (.A(_0775_),
    .X(_0944_));
 sky130_fd_sc_hd__buf_8 _2553_ (.A(_0808_),
    .X(_0945_));
 sky130_fd_sc_hd__mux4_1 _2554_ (.A0(\tms1x00.RAM[80][1] ),
    .A1(\tms1x00.RAM[81][1] ),
    .A2(\tms1x00.RAM[82][1] ),
    .A3(\tms1x00.RAM[83][1] ),
    .S0(_0945_),
    .S1(_0791_),
    .X(_0946_));
 sky130_fd_sc_hd__mux4_1 _2555_ (.A0(\tms1x00.RAM[84][1] ),
    .A1(\tms1x00.RAM[85][1] ),
    .A2(\tms1x00.RAM[86][1] ),
    .A3(\tms1x00.RAM[87][1] ),
    .S0(_0945_),
    .S1(_0791_),
    .X(_0947_));
 sky130_fd_sc_hd__clkbuf_4 _2556_ (.A(_0783_),
    .X(_0948_));
 sky130_fd_sc_hd__mux2_1 _2557_ (.A0(_0946_),
    .A1(_0947_),
    .S(_0948_),
    .X(_0949_));
 sky130_fd_sc_hd__mux2_1 _2558_ (.A0(\tms1x00.RAM[92][1] ),
    .A1(\tms1x00.RAM[93][1] ),
    .S(_0816_),
    .X(_0950_));
 sky130_fd_sc_hd__and2_1 _2559_ (.A(_0818_),
    .B(_0950_),
    .X(_0951_));
 sky130_fd_sc_hd__mux2_1 _2560_ (.A0(\tms1x00.RAM[94][1] ),
    .A1(\tms1x00.RAM[95][1] ),
    .S(_0923_),
    .X(_0952_));
 sky130_fd_sc_hd__buf_4 _2561_ (.A(_0794_),
    .X(_0953_));
 sky130_fd_sc_hd__a21o_1 _2562_ (.A1(_0928_),
    .A2(_0952_),
    .B1(_0953_),
    .X(_0954_));
 sky130_fd_sc_hd__buf_8 _2563_ (.A(_0799_),
    .X(_0955_));
 sky130_fd_sc_hd__buf_6 _2564_ (.A(_0800_),
    .X(_0956_));
 sky130_fd_sc_hd__mux4_1 _2565_ (.A0(\tms1x00.RAM[88][1] ),
    .A1(\tms1x00.RAM[89][1] ),
    .A2(\tms1x00.RAM[90][1] ),
    .A3(\tms1x00.RAM[91][1] ),
    .S0(_0955_),
    .S1(_0956_),
    .X(_0957_));
 sky130_fd_sc_hd__o221a_1 _2566_ (.A1(_0951_),
    .A2(_0954_),
    .B1(_0957_),
    .B2(_0948_),
    .C1(_0942_),
    .X(_0958_));
 sky130_fd_sc_hd__a211oi_1 _2567_ (.A1(_0944_),
    .A2(_0949_),
    .B1(_0958_),
    .C1(_0920_),
    .Y(_0959_));
 sky130_fd_sc_hd__a311o_1 _2568_ (.A1(_0920_),
    .A2(_0935_),
    .A3(_0943_),
    .B1(_0040_),
    .C1(_0959_),
    .X(_0960_));
 sky130_fd_sc_hd__mux4_1 _2569_ (.A0(\tms1x00.RAM[100][1] ),
    .A1(\tms1x00.RAM[101][1] ),
    .A2(\tms1x00.RAM[102][1] ),
    .A3(\tms1x00.RAM[103][1] ),
    .S0(_0945_),
    .S1(_0791_),
    .X(_0961_));
 sky130_fd_sc_hd__or2_1 _2570_ (.A(_0940_),
    .B(_0961_),
    .X(_0962_));
 sky130_fd_sc_hd__mux4_1 _2571_ (.A0(\tms1x00.RAM[96][1] ),
    .A1(\tms1x00.RAM[97][1] ),
    .A2(\tms1x00.RAM[98][1] ),
    .A3(\tms1x00.RAM[99][1] ),
    .S0(_0945_),
    .S1(_0791_),
    .X(_0963_));
 sky130_fd_sc_hd__or2_1 _2572_ (.A(_0948_),
    .B(_0963_),
    .X(_0964_));
 sky130_fd_sc_hd__mux4_1 _2573_ (.A0(\tms1x00.RAM[108][1] ),
    .A1(\tms1x00.RAM[109][1] ),
    .A2(\tms1x00.RAM[110][1] ),
    .A3(\tms1x00.RAM[111][1] ),
    .S0(_0955_),
    .S1(_0956_),
    .X(_0965_));
 sky130_fd_sc_hd__mux4_1 _2574_ (.A0(\tms1x00.RAM[104][1] ),
    .A1(\tms1x00.RAM[105][1] ),
    .A2(\tms1x00.RAM[106][1] ),
    .A3(\tms1x00.RAM[107][1] ),
    .S0(_0799_),
    .S1(_0813_),
    .X(_0966_));
 sky130_fd_sc_hd__or2_1 _2575_ (.A(_0798_),
    .B(_0966_),
    .X(_0967_));
 sky130_fd_sc_hd__o211a_1 _2576_ (.A1(_0940_),
    .A2(_0965_),
    .B1(_0967_),
    .C1(_0942_),
    .X(_0968_));
 sky130_fd_sc_hd__a311o_1 _2577_ (.A1(_0944_),
    .A2(_0962_),
    .A3(_0964_),
    .B1(_0821_),
    .C1(_0968_),
    .X(_0969_));
 sky130_fd_sc_hd__mux4_1 _2578_ (.A0(\tms1x00.RAM[124][1] ),
    .A1(\tms1x00.RAM[125][1] ),
    .A2(\tms1x00.RAM[126][1] ),
    .A3(\tms1x00.RAM[127][1] ),
    .S0(_0945_),
    .S1(_0956_),
    .X(_0970_));
 sky130_fd_sc_hd__mux4_2 _2579_ (.A0(\tms1x00.RAM[120][1] ),
    .A1(\tms1x00.RAM[121][1] ),
    .A2(\tms1x00.RAM[122][1] ),
    .A3(\tms1x00.RAM[123][1] ),
    .S0(_0808_),
    .S1(_0831_),
    .X(_0971_));
 sky130_fd_sc_hd__or2_1 _2580_ (.A(_0807_),
    .B(_0971_),
    .X(_0972_));
 sky130_fd_sc_hd__o211a_1 _2581_ (.A1(_0940_),
    .A2(_0970_),
    .B1(_0972_),
    .C1(_0806_),
    .X(_0973_));
 sky130_fd_sc_hd__mux4_2 _2582_ (.A0(\tms1x00.RAM[112][1] ),
    .A1(\tms1x00.RAM[113][1] ),
    .A2(\tms1x00.RAM[114][1] ),
    .A3(\tms1x00.RAM[115][1] ),
    .S0(_0955_),
    .S1(_0956_),
    .X(_0974_));
 sky130_fd_sc_hd__clkbuf_8 _2583_ (.A(_0778_),
    .X(_0975_));
 sky130_fd_sc_hd__or2b_1 _2584_ (.A(\tms1x00.RAM[119][1] ),
    .B_N(_0975_),
    .X(_0976_));
 sky130_fd_sc_hd__buf_6 _2585_ (.A(_0850_),
    .X(_0977_));
 sky130_fd_sc_hd__o21a_1 _2586_ (.A1(_0975_),
    .A2(\tms1x00.RAM[118][1] ),
    .B1(_0977_),
    .X(_0978_));
 sky130_fd_sc_hd__mux2_1 _2587_ (.A0(\tms1x00.RAM[116][1] ),
    .A1(\tms1x00.RAM[117][1] ),
    .S(_0923_),
    .X(_0979_));
 sky130_fd_sc_hd__a221o_1 _2588_ (.A1(_0976_),
    .A2(_0978_),
    .B1(_0979_),
    .B2(_0818_),
    .C1(_0819_),
    .X(_0980_));
 sky130_fd_sc_hd__o211a_1 _2589_ (.A1(_0948_),
    .A2(_0974_),
    .B1(_0980_),
    .C1(_0776_),
    .X(_0981_));
 sky130_fd_sc_hd__o31a_1 _2590_ (.A1(_0920_),
    .A2(_0973_),
    .A3(_0981_),
    .B1(_0040_),
    .X(_0982_));
 sky130_fd_sc_hd__a21oi_1 _2591_ (.A1(_0969_),
    .A2(_0982_),
    .B1(_0835_),
    .Y(_0983_));
 sky130_fd_sc_hd__mux4_1 _2592_ (.A0(\tms1x00.RAM[16][1] ),
    .A1(\tms1x00.RAM[17][1] ),
    .A2(\tms1x00.RAM[18][1] ),
    .A3(\tms1x00.RAM[19][1] ),
    .S0(_0975_),
    .S1(_0791_),
    .X(_0984_));
 sky130_fd_sc_hd__mux4_2 _2593_ (.A0(\tms1x00.RAM[20][1] ),
    .A1(\tms1x00.RAM[21][1] ),
    .A2(\tms1x00.RAM[22][1] ),
    .A3(\tms1x00.RAM[23][1] ),
    .S0(_0975_),
    .S1(_0791_),
    .X(_0985_));
 sky130_fd_sc_hd__mux2_1 _2594_ (.A0(_0984_),
    .A1(_0985_),
    .S(_0921_),
    .X(_0986_));
 sky130_fd_sc_hd__mux2_1 _2595_ (.A0(\tms1x00.RAM[28][1] ),
    .A1(\tms1x00.RAM[29][1] ),
    .S(_0873_),
    .X(_0987_));
 sky130_fd_sc_hd__and2_1 _2596_ (.A(_0818_),
    .B(_0987_),
    .X(_0988_));
 sky130_fd_sc_hd__mux2_1 _2597_ (.A0(\tms1x00.RAM[30][1] ),
    .A1(\tms1x00.RAM[31][1] ),
    .S(_0816_),
    .X(_0989_));
 sky130_fd_sc_hd__a21o_1 _2598_ (.A1(_0932_),
    .A2(_0989_),
    .B1(_0819_),
    .X(_0990_));
 sky130_fd_sc_hd__mux4_2 _2599_ (.A0(\tms1x00.RAM[24][1] ),
    .A1(\tms1x00.RAM[25][1] ),
    .A2(\tms1x00.RAM[26][1] ),
    .A3(\tms1x00.RAM[27][1] ),
    .S0(_0945_),
    .S1(_0791_),
    .X(_0991_));
 sky130_fd_sc_hd__o221a_1 _2600_ (.A1(_0988_),
    .A2(_0990_),
    .B1(_0991_),
    .B2(_0948_),
    .C1(_0806_),
    .X(_0992_));
 sky130_fd_sc_hd__a211oi_1 _2601_ (.A1(_0944_),
    .A2(_0986_),
    .B1(_0992_),
    .C1(_0920_),
    .Y(_0993_));
 sky130_fd_sc_hd__mux2_1 _2602_ (.A0(\tms1x00.RAM[4][1] ),
    .A1(\tms1x00.RAM[5][1] ),
    .S(_0924_),
    .X(_0994_));
 sky130_fd_sc_hd__mux2_1 _2603_ (.A0(\tms1x00.RAM[6][1] ),
    .A1(\tms1x00.RAM[7][1] ),
    .S(_0975_),
    .X(_0995_));
 sky130_fd_sc_hd__clkbuf_4 _2604_ (.A(_0794_),
    .X(_0996_));
 sky130_fd_sc_hd__a21o_1 _2605_ (.A1(_0928_),
    .A2(_0995_),
    .B1(_0996_),
    .X(_0997_));
 sky130_fd_sc_hd__a21oi_1 _2606_ (.A1(_0787_),
    .A2(_0994_),
    .B1(_0997_),
    .Y(_0998_));
 sky130_fd_sc_hd__mux4_1 _2607_ (.A0(\tms1x00.RAM[0][1] ),
    .A1(\tms1x00.RAM[1][1] ),
    .A2(\tms1x00.RAM[2][1] ),
    .A3(\tms1x00.RAM[3][1] ),
    .S0(_0955_),
    .S1(_0956_),
    .X(_0999_));
 sky130_fd_sc_hd__o21ai_1 _2608_ (.A1(_0948_),
    .A2(_0999_),
    .B1(_0776_),
    .Y(_1000_));
 sky130_fd_sc_hd__mux2_1 _2609_ (.A0(\tms1x00.RAM[14][1] ),
    .A1(\tms1x00.RAM[15][1] ),
    .S(_0924_),
    .X(_1001_));
 sky130_fd_sc_hd__mux2_1 _2610_ (.A0(\tms1x00.RAM[12][1] ),
    .A1(\tms1x00.RAM[13][1] ),
    .S(_0975_),
    .X(_1002_));
 sky130_fd_sc_hd__a21o_1 _2611_ (.A1(_0787_),
    .A2(_1002_),
    .B1(_0996_),
    .X(_1003_));
 sky130_fd_sc_hd__a21oi_1 _2612_ (.A1(_0928_),
    .A2(_1001_),
    .B1(_1003_),
    .Y(_1004_));
 sky130_fd_sc_hd__mux4_1 _2613_ (.A0(\tms1x00.RAM[8][1] ),
    .A1(\tms1x00.RAM[9][1] ),
    .A2(\tms1x00.RAM[10][1] ),
    .A3(\tms1x00.RAM[11][1] ),
    .S0(_0931_),
    .S1(_0956_),
    .X(_1005_));
 sky130_fd_sc_hd__o21ai_1 _2614_ (.A1(_0948_),
    .A2(_1005_),
    .B1(_0942_),
    .Y(_1006_));
 sky130_fd_sc_hd__o221a_1 _2615_ (.A1(_0998_),
    .A2(_1000_),
    .B1(_1004_),
    .B2(_1006_),
    .C1(_0920_),
    .X(_1007_));
 sky130_fd_sc_hd__mux4_1 _2616_ (.A0(\tms1x00.RAM[44][1] ),
    .A1(\tms1x00.RAM[45][1] ),
    .A2(\tms1x00.RAM[46][1] ),
    .A3(\tms1x00.RAM[47][1] ),
    .S0(_0799_),
    .S1(_0800_),
    .X(_1008_));
 sky130_fd_sc_hd__nor2_1 _2617_ (.A(_0953_),
    .B(_1008_),
    .Y(_1009_));
 sky130_fd_sc_hd__mux4_1 _2618_ (.A0(\tms1x00.RAM[40][1] ),
    .A1(\tms1x00.RAM[41][1] ),
    .A2(\tms1x00.RAM[42][1] ),
    .A3(\tms1x00.RAM[43][1] ),
    .S0(_0808_),
    .S1(_0780_),
    .X(_1010_));
 sky130_fd_sc_hd__o21ai_1 _2619_ (.A1(_0807_),
    .A2(_1010_),
    .B1(_0802_),
    .Y(_1011_));
 sky130_fd_sc_hd__mux4_1 _2620_ (.A0(\tms1x00.RAM[32][1] ),
    .A1(\tms1x00.RAM[33][1] ),
    .A2(\tms1x00.RAM[34][1] ),
    .A3(\tms1x00.RAM[35][1] ),
    .S0(_0840_),
    .S1(_0813_),
    .X(_1012_));
 sky130_fd_sc_hd__nor2_1 _2621_ (.A(_0798_),
    .B(_1012_),
    .Y(_1013_));
 sky130_fd_sc_hd__mux4_2 _2622_ (.A0(\tms1x00.RAM[36][1] ),
    .A1(\tms1x00.RAM[37][1] ),
    .A2(\tms1x00.RAM[38][1] ),
    .A3(\tms1x00.RAM[39][1] ),
    .S0(_0808_),
    .S1(_0831_),
    .X(_1014_));
 sky130_fd_sc_hd__o21ai_1 _2623_ (.A1(_0819_),
    .A2(_1014_),
    .B1(_0775_),
    .Y(_1015_));
 sky130_fd_sc_hd__o221a_1 _2624_ (.A1(_1009_),
    .A2(_1011_),
    .B1(_1013_),
    .B2(_1015_),
    .C1(_0804_),
    .X(_1016_));
 sky130_fd_sc_hd__mux4_1 _2625_ (.A0(\tms1x00.RAM[56][1] ),
    .A1(\tms1x00.RAM[57][1] ),
    .A2(\tms1x00.RAM[58][1] ),
    .A3(\tms1x00.RAM[59][1] ),
    .S0(_0823_),
    .S1(_0850_),
    .X(_1017_));
 sky130_fd_sc_hd__or2_1 _2626_ (.A(_0783_),
    .B(_1017_),
    .X(_1018_));
 sky130_fd_sc_hd__mux4_1 _2627_ (.A0(\tms1x00.RAM[60][1] ),
    .A1(\tms1x00.RAM[61][1] ),
    .A2(\tms1x00.RAM[62][1] ),
    .A3(\tms1x00.RAM[63][1] ),
    .S0(_0826_),
    .S1(_0850_),
    .X(_1019_));
 sky130_fd_sc_hd__o21a_1 _2628_ (.A1(_0794_),
    .A2(_1019_),
    .B1(_0038_),
    .X(_1020_));
 sky130_fd_sc_hd__or2b_1 _2629_ (.A(\tms1x00.RAM[55][1] ),
    .B_N(_0873_),
    .X(_1021_));
 sky130_fd_sc_hd__o21a_1 _2630_ (.A1(_0840_),
    .A2(\tms1x00.RAM[54][1] ),
    .B1(_0780_),
    .X(_1022_));
 sky130_fd_sc_hd__mux2_1 _2631_ (.A0(\tms1x00.RAM[52][1] ),
    .A1(\tms1x00.RAM[53][1] ),
    .S(_0778_),
    .X(_1023_));
 sky130_fd_sc_hd__a221o_1 _2632_ (.A1(_1021_),
    .A2(_1022_),
    .B1(_1023_),
    .B2(_0818_),
    .C1(_0794_),
    .X(_1024_));
 sky130_fd_sc_hd__mux4_1 _2633_ (.A0(\tms1x00.RAM[48][1] ),
    .A1(\tms1x00.RAM[49][1] ),
    .A2(\tms1x00.RAM[50][1] ),
    .A3(\tms1x00.RAM[51][1] ),
    .S0(_0788_),
    .S1(_0780_),
    .X(_1025_));
 sky130_fd_sc_hd__o21a_1 _2634_ (.A1(_0783_),
    .A2(_1025_),
    .B1(_0774_),
    .X(_1026_));
 sky130_fd_sc_hd__a221o_1 _2635_ (.A1(_1018_),
    .A2(_1020_),
    .B1(_1024_),
    .B2(_1026_),
    .C1(_0804_),
    .X(_1027_));
 sky130_fd_sc_hd__or3b_1 _2636_ (.A(_0773_),
    .B(_1016_),
    .C_N(_1027_),
    .X(_1028_));
 sky130_fd_sc_hd__o311a_1 _2637_ (.A1(_0040_),
    .A2(_0993_),
    .A3(_1007_),
    .B1(_1028_),
    .C1(_0835_),
    .X(_1029_));
 sky130_fd_sc_hd__a21oi_2 _2638_ (.A1(_0960_),
    .A2(_0983_),
    .B1(_1029_),
    .Y(_1030_));
 sky130_fd_sc_hd__and2b_1 _2639_ (.A_N(_0747_),
    .B(_0748_),
    .X(_1031_));
 sky130_fd_sc_hd__inv_2 _2640_ (.A(_1031_),
    .Y(_1032_));
 sky130_fd_sc_hd__a32o_1 _2641_ (.A1(_0771_),
    .A2(_1030_),
    .A3(_1032_),
    .B1(_0909_),
    .B2(\tms1x00.A[1] ),
    .X(_1033_));
 sky130_fd_sc_hd__buf_4 _2642_ (.A(_1033_),
    .X(_1034_));
 sky130_fd_sc_hd__clkbuf_4 _2643_ (.A(_1034_),
    .X(_1035_));
 sky130_fd_sc_hd__mux2_1 _2644_ (.A0(_1035_),
    .A1(\tms1x00.RAM[109][1] ),
    .S(_0918_),
    .X(_1036_));
 sky130_fd_sc_hd__clkbuf_1 _2645_ (.A(_1036_),
    .X(_0052_));
 sky130_fd_sc_hd__mux4_2 _2646_ (.A0(\tms1x00.RAM[44][2] ),
    .A1(\tms1x00.RAM[45][2] ),
    .A2(\tms1x00.RAM[46][2] ),
    .A3(\tms1x00.RAM[47][2] ),
    .S0(_0955_),
    .S1(_0956_),
    .X(_1037_));
 sky130_fd_sc_hd__mux4_1 _2647_ (.A0(\tms1x00.RAM[40][2] ),
    .A1(\tms1x00.RAM[41][2] ),
    .A2(\tms1x00.RAM[42][2] ),
    .A3(\tms1x00.RAM[43][2] ),
    .S0(_0830_),
    .S1(_0831_),
    .X(_1038_));
 sky130_fd_sc_hd__or2_1 _2648_ (.A(_0807_),
    .B(_1038_),
    .X(_1039_));
 sky130_fd_sc_hd__o211a_1 _2649_ (.A1(_0940_),
    .A2(_1037_),
    .B1(_1039_),
    .C1(_0942_),
    .X(_1040_));
 sky130_fd_sc_hd__mux4_2 _2650_ (.A0(\tms1x00.RAM[32][2] ),
    .A1(\tms1x00.RAM[33][2] ),
    .A2(\tms1x00.RAM[34][2] ),
    .A3(\tms1x00.RAM[35][2] ),
    .S0(_0955_),
    .S1(_0956_),
    .X(_1041_));
 sky130_fd_sc_hd__mux4_2 _2651_ (.A0(\tms1x00.RAM[36][2] ),
    .A1(\tms1x00.RAM[37][2] ),
    .A2(\tms1x00.RAM[38][2] ),
    .A3(\tms1x00.RAM[39][2] ),
    .S0(_0799_),
    .S1(_0800_),
    .X(_1042_));
 sky130_fd_sc_hd__or2_1 _2652_ (.A(_0819_),
    .B(_1042_),
    .X(_1043_));
 sky130_fd_sc_hd__o211a_1 _2653_ (.A1(_0948_),
    .A2(_1041_),
    .B1(_1043_),
    .C1(_0776_),
    .X(_1044_));
 sky130_fd_sc_hd__or2b_1 _2654_ (.A(\tms1x00.RAM[55][2] ),
    .B_N(_0975_),
    .X(_1045_));
 sky130_fd_sc_hd__o21a_1 _2655_ (.A1(_0975_),
    .A2(\tms1x00.RAM[54][2] ),
    .B1(_0977_),
    .X(_1046_));
 sky130_fd_sc_hd__mux2_1 _2656_ (.A0(\tms1x00.RAM[52][2] ),
    .A1(\tms1x00.RAM[53][2] ),
    .S(_0923_),
    .X(_1047_));
 sky130_fd_sc_hd__a221o_1 _2657_ (.A1(_1045_),
    .A2(_1046_),
    .B1(_1047_),
    .B2(_0818_),
    .C1(_0953_),
    .X(_1048_));
 sky130_fd_sc_hd__mux4_2 _2658_ (.A0(\tms1x00.RAM[48][2] ),
    .A1(\tms1x00.RAM[49][2] ),
    .A2(\tms1x00.RAM[50][2] ),
    .A3(\tms1x00.RAM[51][2] ),
    .S0(_0799_),
    .S1(_0800_),
    .X(_1049_));
 sky130_fd_sc_hd__or2_1 _2659_ (.A(_0798_),
    .B(_1049_),
    .X(_1050_));
 sky130_fd_sc_hd__mux4_1 _2660_ (.A0(\tms1x00.RAM[60][2] ),
    .A1(\tms1x00.RAM[61][2] ),
    .A2(\tms1x00.RAM[62][2] ),
    .A3(\tms1x00.RAM[63][2] ),
    .S0(_0840_),
    .S1(_0822_),
    .X(_1051_));
 sky130_fd_sc_hd__mux4_1 _2661_ (.A0(\tms1x00.RAM[56][2] ),
    .A1(\tms1x00.RAM[57][2] ),
    .A2(\tms1x00.RAM[58][2] ),
    .A3(\tms1x00.RAM[59][2] ),
    .S0(_0815_),
    .S1(_0812_),
    .X(_1052_));
 sky130_fd_sc_hd__or2_1 _2662_ (.A(_0797_),
    .B(_1052_),
    .X(_1053_));
 sky130_fd_sc_hd__o211a_1 _2663_ (.A1(_0953_),
    .A2(_1051_),
    .B1(_1053_),
    .C1(_0802_),
    .X(_1054_));
 sky130_fd_sc_hd__a311o_1 _2664_ (.A1(_0776_),
    .A2(_1048_),
    .A3(_1050_),
    .B1(_0804_),
    .C1(_1054_),
    .X(_1055_));
 sky130_fd_sc_hd__o311a_1 _2665_ (.A1(_0821_),
    .A2(_1040_),
    .A3(_1044_),
    .B1(_0040_),
    .C1(_1055_),
    .X(_1056_));
 sky130_fd_sc_hd__mux4_2 _2666_ (.A0(\tms1x00.RAM[16][2] ),
    .A1(\tms1x00.RAM[17][2] ),
    .A2(\tms1x00.RAM[18][2] ),
    .A3(\tms1x00.RAM[19][2] ),
    .S0(_0955_),
    .S1(_0956_),
    .X(_1057_));
 sky130_fd_sc_hd__mux4_2 _2667_ (.A0(\tms1x00.RAM[20][2] ),
    .A1(\tms1x00.RAM[21][2] ),
    .A2(\tms1x00.RAM[22][2] ),
    .A3(\tms1x00.RAM[23][2] ),
    .S0(_0799_),
    .S1(_0800_),
    .X(_1058_));
 sky130_fd_sc_hd__or2_1 _2668_ (.A(_0819_),
    .B(_1058_),
    .X(_1059_));
 sky130_fd_sc_hd__o211a_1 _2669_ (.A1(_0948_),
    .A2(_1057_),
    .B1(_1059_),
    .C1(_0776_),
    .X(_1060_));
 sky130_fd_sc_hd__mux2_1 _2670_ (.A0(\tms1x00.RAM[30][2] ),
    .A1(\tms1x00.RAM[31][2] ),
    .S(_0923_),
    .X(_1061_));
 sky130_fd_sc_hd__and2_1 _2671_ (.A(_0932_),
    .B(_1061_),
    .X(_1062_));
 sky130_fd_sc_hd__mux2_1 _2672_ (.A0(\tms1x00.RAM[28][2] ),
    .A1(\tms1x00.RAM[29][2] ),
    .S(_0789_),
    .X(_1063_));
 sky130_fd_sc_hd__a21o_1 _2673_ (.A1(_0818_),
    .A2(_1063_),
    .B1(_0953_),
    .X(_1064_));
 sky130_fd_sc_hd__mux4_2 _2674_ (.A0(\tms1x00.RAM[24][2] ),
    .A1(\tms1x00.RAM[25][2] ),
    .A2(\tms1x00.RAM[26][2] ),
    .A3(\tms1x00.RAM[27][2] ),
    .S0(_0955_),
    .S1(_0956_),
    .X(_1065_));
 sky130_fd_sc_hd__o221a_1 _2675_ (.A1(_1062_),
    .A2(_1064_),
    .B1(_1065_),
    .B2(_0948_),
    .C1(_0942_),
    .X(_1066_));
 sky130_fd_sc_hd__mux2_1 _2676_ (.A0(\tms1x00.RAM[6][2] ),
    .A1(\tms1x00.RAM[7][2] ),
    .S(_0815_),
    .X(_1067_));
 sky130_fd_sc_hd__and2_1 _2677_ (.A(_0813_),
    .B(_1067_),
    .X(_1068_));
 sky130_fd_sc_hd__mux2_1 _2678_ (.A0(\tms1x00.RAM[4][2] ),
    .A1(\tms1x00.RAM[5][2] ),
    .S(_0823_),
    .X(_1069_));
 sky130_fd_sc_hd__a21o_1 _2679_ (.A1(_0785_),
    .A2(_1069_),
    .B1(_0793_),
    .X(_1070_));
 sky130_fd_sc_hd__mux4_1 _2680_ (.A0(\tms1x00.RAM[0][2] ),
    .A1(\tms1x00.RAM[1][2] ),
    .A2(\tms1x00.RAM[2][2] ),
    .A3(\tms1x00.RAM[3][2] ),
    .S0(_0808_),
    .S1(_0831_),
    .X(_1071_));
 sky130_fd_sc_hd__o221a_1 _2681_ (.A1(_1068_),
    .A2(_1070_),
    .B1(_1071_),
    .B2(_0807_),
    .C1(_0774_),
    .X(_1072_));
 sky130_fd_sc_hd__mux4_1 _2682_ (.A0(\tms1x00.RAM[8][2] ),
    .A1(\tms1x00.RAM[9][2] ),
    .A2(\tms1x00.RAM[10][2] ),
    .A3(\tms1x00.RAM[11][2] ),
    .S0(_0830_),
    .S1(_0800_),
    .X(_1073_));
 sky130_fd_sc_hd__or2b_1 _2683_ (.A(\tms1x00.RAM[15][2] ),
    .B_N(_0788_),
    .X(_1074_));
 sky130_fd_sc_hd__o21a_1 _2684_ (.A1(_0788_),
    .A2(\tms1x00.RAM[14][2] ),
    .B1(_0812_),
    .X(_1075_));
 sky130_fd_sc_hd__mux2_1 _2685_ (.A0(\tms1x00.RAM[12][2] ),
    .A1(\tms1x00.RAM[13][2] ),
    .S(_0823_),
    .X(_1076_));
 sky130_fd_sc_hd__a221o_1 _2686_ (.A1(_1074_),
    .A2(_1075_),
    .B1(_1076_),
    .B2(_0785_),
    .C1(_0793_),
    .X(_1077_));
 sky130_fd_sc_hd__o211a_1 _2687_ (.A1(_0807_),
    .A2(_1073_),
    .B1(_1077_),
    .C1(_0802_),
    .X(_1078_));
 sky130_fd_sc_hd__or3_1 _2688_ (.A(_0039_),
    .B(_1072_),
    .C(_1078_),
    .X(_1079_));
 sky130_fd_sc_hd__o311a_1 _2689_ (.A1(_0920_),
    .A2(_1060_),
    .A3(_1066_),
    .B1(_1079_),
    .C1(_0773_),
    .X(_1080_));
 sky130_fd_sc_hd__mux4_2 _2690_ (.A0(\tms1x00.RAM[80][2] ),
    .A1(\tms1x00.RAM[81][2] ),
    .A2(\tms1x00.RAM[82][2] ),
    .A3(\tms1x00.RAM[83][2] ),
    .S0(_0931_),
    .S1(_0932_),
    .X(_1081_));
 sky130_fd_sc_hd__mux4_1 _2691_ (.A0(\tms1x00.RAM[84][2] ),
    .A1(\tms1x00.RAM[85][2] ),
    .A2(\tms1x00.RAM[86][2] ),
    .A3(\tms1x00.RAM[87][2] ),
    .S0(_0873_),
    .S1(_0977_),
    .X(_1082_));
 sky130_fd_sc_hd__or2_1 _2692_ (.A(_0953_),
    .B(_1082_),
    .X(_1083_));
 sky130_fd_sc_hd__o211a_1 _2693_ (.A1(_0922_),
    .A2(_1081_),
    .B1(_1083_),
    .C1(_0944_),
    .X(_1084_));
 sky130_fd_sc_hd__mux2_1 _2694_ (.A0(\tms1x00.RAM[94][2] ),
    .A1(\tms1x00.RAM[95][2] ),
    .S(_0789_),
    .X(_1085_));
 sky130_fd_sc_hd__and2_1 _2695_ (.A(_0928_),
    .B(_1085_),
    .X(_1086_));
 sky130_fd_sc_hd__mux2_1 _2696_ (.A0(\tms1x00.RAM[92][2] ),
    .A1(\tms1x00.RAM[93][2] ),
    .S(_0975_),
    .X(_1087_));
 sky130_fd_sc_hd__a21o_1 _2697_ (.A1(_0787_),
    .A2(_1087_),
    .B1(_0996_),
    .X(_1088_));
 sky130_fd_sc_hd__mux4_1 _2698_ (.A0(\tms1x00.RAM[88][2] ),
    .A1(\tms1x00.RAM[89][2] ),
    .A2(\tms1x00.RAM[90][2] ),
    .A3(\tms1x00.RAM[91][2] ),
    .S0(_0931_),
    .S1(_0932_),
    .X(_1089_));
 sky130_fd_sc_hd__o221a_1 _2699_ (.A1(_1086_),
    .A2(_1088_),
    .B1(_1089_),
    .B2(_0922_),
    .C1(_0942_),
    .X(_1090_));
 sky130_fd_sc_hd__mux2_1 _2700_ (.A0(\tms1x00.RAM[70][2] ),
    .A1(\tms1x00.RAM[71][2] ),
    .S(_0788_),
    .X(_1091_));
 sky130_fd_sc_hd__and2_1 _2701_ (.A(_0977_),
    .B(_1091_),
    .X(_1092_));
 sky130_fd_sc_hd__mux2_1 _2702_ (.A0(\tms1x00.RAM[68][2] ),
    .A1(\tms1x00.RAM[69][2] ),
    .S(_0788_),
    .X(_1093_));
 sky130_fd_sc_hd__a21o_1 _2703_ (.A1(_0786_),
    .A2(_1093_),
    .B1(_0794_),
    .X(_1094_));
 sky130_fd_sc_hd__mux4_1 _2704_ (.A0(\tms1x00.RAM[64][2] ),
    .A1(\tms1x00.RAM[65][2] ),
    .A2(\tms1x00.RAM[66][2] ),
    .A3(\tms1x00.RAM[67][2] ),
    .S0(_0840_),
    .S1(_0813_),
    .X(_1095_));
 sky130_fd_sc_hd__o221a_1 _2705_ (.A1(_1092_),
    .A2(_1094_),
    .B1(_1095_),
    .B2(_0798_),
    .C1(_0775_),
    .X(_1096_));
 sky130_fd_sc_hd__mux4_1 _2706_ (.A0(\tms1x00.RAM[72][2] ),
    .A1(\tms1x00.RAM[73][2] ),
    .A2(\tms1x00.RAM[74][2] ),
    .A3(\tms1x00.RAM[75][2] ),
    .S0(_0873_),
    .S1(_0822_),
    .X(_1097_));
 sky130_fd_sc_hd__or2b_1 _2707_ (.A(\tms1x00.RAM[79][2] ),
    .B_N(_0830_),
    .X(_1098_));
 sky130_fd_sc_hd__o21a_1 _2708_ (.A1(_0830_),
    .A2(\tms1x00.RAM[78][2] ),
    .B1(_0850_),
    .X(_1099_));
 sky130_fd_sc_hd__mux2_1 _2709_ (.A0(\tms1x00.RAM[76][2] ),
    .A1(\tms1x00.RAM[77][2] ),
    .S(_0788_),
    .X(_1100_));
 sky130_fd_sc_hd__a221o_1 _2710_ (.A1(_1098_),
    .A2(_1099_),
    .B1(_1100_),
    .B2(_0786_),
    .C1(_0794_),
    .X(_1101_));
 sky130_fd_sc_hd__o211a_1 _2711_ (.A1(_0921_),
    .A2(_1097_),
    .B1(_1101_),
    .C1(_0802_),
    .X(_1102_));
 sky130_fd_sc_hd__or3_1 _2712_ (.A(_0821_),
    .B(_1096_),
    .C(_1102_),
    .X(_1103_));
 sky130_fd_sc_hd__o311a_1 _2713_ (.A1(_0920_),
    .A2(_1084_),
    .A3(_1090_),
    .B1(_1103_),
    .C1(_0773_),
    .X(_1104_));
 sky130_fd_sc_hd__or2b_1 _2714_ (.A(\tms1x00.RAM[119][2] ),
    .B_N(_0945_),
    .X(_1105_));
 sky130_fd_sc_hd__o21a_1 _2715_ (.A1(_0945_),
    .A2(\tms1x00.RAM[118][2] ),
    .B1(_0927_),
    .X(_1106_));
 sky130_fd_sc_hd__mux2_1 _2716_ (.A0(\tms1x00.RAM[116][2] ),
    .A1(\tms1x00.RAM[117][2] ),
    .S(_0789_),
    .X(_1107_));
 sky130_fd_sc_hd__a221o_1 _2717_ (.A1(_1105_),
    .A2(_1106_),
    .B1(_1107_),
    .B2(_0818_),
    .C1(_0953_),
    .X(_1108_));
 sky130_fd_sc_hd__mux4_1 _2718_ (.A0(\tms1x00.RAM[112][2] ),
    .A1(\tms1x00.RAM[113][2] ),
    .A2(\tms1x00.RAM[114][2] ),
    .A3(\tms1x00.RAM[115][2] ),
    .S0(_0873_),
    .S1(_0822_),
    .X(_1109_));
 sky130_fd_sc_hd__or2_1 _2719_ (.A(_0921_),
    .B(_1109_),
    .X(_1110_));
 sky130_fd_sc_hd__mux4_1 _2720_ (.A0(\tms1x00.RAM[124][2] ),
    .A1(\tms1x00.RAM[125][2] ),
    .A2(\tms1x00.RAM[126][2] ),
    .A3(\tms1x00.RAM[127][2] ),
    .S0(_0816_),
    .S1(_0977_),
    .X(_1111_));
 sky130_fd_sc_hd__mux4_1 _2721_ (.A0(\tms1x00.RAM[120][2] ),
    .A1(\tms1x00.RAM[121][2] ),
    .A2(\tms1x00.RAM[122][2] ),
    .A3(\tms1x00.RAM[123][2] ),
    .S0(_0823_),
    .S1(_0850_),
    .X(_1112_));
 sky130_fd_sc_hd__or2_1 _2722_ (.A(_0783_),
    .B(_1112_),
    .X(_1113_));
 sky130_fd_sc_hd__o211a_1 _2723_ (.A1(_0996_),
    .A2(_1111_),
    .B1(_1113_),
    .C1(_0806_),
    .X(_1114_));
 sky130_fd_sc_hd__a311o_1 _2724_ (.A1(_0944_),
    .A2(_1108_),
    .A3(_1110_),
    .B1(_0804_),
    .C1(_1114_),
    .X(_1115_));
 sky130_fd_sc_hd__mux4_1 _2725_ (.A0(\tms1x00.RAM[100][2] ),
    .A1(\tms1x00.RAM[101][2] ),
    .A2(\tms1x00.RAM[102][2] ),
    .A3(\tms1x00.RAM[103][2] ),
    .S0(_0873_),
    .S1(_0822_),
    .X(_1116_));
 sky130_fd_sc_hd__or2_1 _2726_ (.A(_0953_),
    .B(_1116_),
    .X(_1117_));
 sky130_fd_sc_hd__mux4_2 _2727_ (.A0(\tms1x00.RAM[96][2] ),
    .A1(\tms1x00.RAM[97][2] ),
    .A2(\tms1x00.RAM[98][2] ),
    .A3(\tms1x00.RAM[99][2] ),
    .S0(_0873_),
    .S1(_0822_),
    .X(_1118_));
 sky130_fd_sc_hd__or2_1 _2728_ (.A(_0921_),
    .B(_1118_),
    .X(_1119_));
 sky130_fd_sc_hd__mux4_1 _2729_ (.A0(\tms1x00.RAM[108][2] ),
    .A1(\tms1x00.RAM[109][2] ),
    .A2(\tms1x00.RAM[110][2] ),
    .A3(\tms1x00.RAM[111][2] ),
    .S0(_0816_),
    .S1(_0977_),
    .X(_1120_));
 sky130_fd_sc_hd__mux4_1 _2730_ (.A0(\tms1x00.RAM[104][2] ),
    .A1(\tms1x00.RAM[105][2] ),
    .A2(\tms1x00.RAM[106][2] ),
    .A3(\tms1x00.RAM[107][2] ),
    .S0(_0823_),
    .S1(_0850_),
    .X(_1121_));
 sky130_fd_sc_hd__or2_1 _2731_ (.A(_0783_),
    .B(_1121_),
    .X(_1122_));
 sky130_fd_sc_hd__o211a_1 _2732_ (.A1(_0996_),
    .A2(_1120_),
    .B1(_1122_),
    .C1(_0806_),
    .X(_1123_));
 sky130_fd_sc_hd__a311o_1 _2733_ (.A1(_0776_),
    .A2(_1117_),
    .A3(_1119_),
    .B1(_0821_),
    .C1(_1123_),
    .X(_1124_));
 sky130_fd_sc_hd__a31o_1 _2734_ (.A1(_0040_),
    .A2(_1115_),
    .A3(_1124_),
    .B1(_0835_),
    .X(_1125_));
 sky130_fd_sc_hd__o32a_1 _2735_ (.A1(_0041_),
    .A2(_1056_),
    .A3(_1080_),
    .B1(_1104_),
    .B2(_1125_),
    .X(_1126_));
 sky130_fd_sc_hd__or2b_1 _2736_ (.A(_0748_),
    .B_N(_0747_),
    .X(_1127_));
 sky130_fd_sc_hd__a32o_1 _2737_ (.A1(_0771_),
    .A2(_1126_),
    .A3(_1127_),
    .B1(_0909_),
    .B2(\tms1x00.A[2] ),
    .X(_1128_));
 sky130_fd_sc_hd__buf_4 _2738_ (.A(_1128_),
    .X(_1129_));
 sky130_fd_sc_hd__buf_4 _2739_ (.A(_1129_),
    .X(_1130_));
 sky130_fd_sc_hd__mux2_1 _2740_ (.A0(_1130_),
    .A1(\tms1x00.RAM[109][2] ),
    .S(_0918_),
    .X(_1131_));
 sky130_fd_sc_hd__clkbuf_1 _2741_ (.A(_1131_),
    .X(_0053_));
 sky130_fd_sc_hd__mux4_1 _2742_ (.A0(\tms1x00.RAM[80][3] ),
    .A1(\tms1x00.RAM[81][3] ),
    .A2(\tms1x00.RAM[82][3] ),
    .A3(\tms1x00.RAM[83][3] ),
    .S0(_0931_),
    .S1(_0932_),
    .X(_1132_));
 sky130_fd_sc_hd__mux4_1 _2743_ (.A0(\tms1x00.RAM[84][3] ),
    .A1(\tms1x00.RAM[85][3] ),
    .A2(\tms1x00.RAM[86][3] ),
    .A3(\tms1x00.RAM[87][3] ),
    .S0(_0840_),
    .S1(_0813_),
    .X(_1133_));
 sky130_fd_sc_hd__or2_1 _2744_ (.A(_0953_),
    .B(_1133_),
    .X(_1134_));
 sky130_fd_sc_hd__o211a_1 _2745_ (.A1(_0922_),
    .A2(_1132_),
    .B1(_1134_),
    .C1(_0776_),
    .X(_1135_));
 sky130_fd_sc_hd__mux2_1 _2746_ (.A0(\tms1x00.RAM[94][3] ),
    .A1(\tms1x00.RAM[95][3] ),
    .S(_0923_),
    .X(_1136_));
 sky130_fd_sc_hd__and2_1 _2747_ (.A(_0928_),
    .B(_1136_),
    .X(_1137_));
 sky130_fd_sc_hd__mux2_1 _2748_ (.A0(\tms1x00.RAM[92][3] ),
    .A1(\tms1x00.RAM[93][3] ),
    .S(_0789_),
    .X(_1138_));
 sky130_fd_sc_hd__a21o_1 _2749_ (.A1(_0787_),
    .A2(_1138_),
    .B1(_0953_),
    .X(_1139_));
 sky130_fd_sc_hd__mux4_1 _2750_ (.A0(\tms1x00.RAM[88][3] ),
    .A1(\tms1x00.RAM[89][3] ),
    .A2(\tms1x00.RAM[90][3] ),
    .A3(\tms1x00.RAM[91][3] ),
    .S0(_0931_),
    .S1(_0932_),
    .X(_1140_));
 sky130_fd_sc_hd__o221a_1 _2751_ (.A1(_1137_),
    .A2(_1139_),
    .B1(_1140_),
    .B2(_0922_),
    .C1(_0942_),
    .X(_1141_));
 sky130_fd_sc_hd__mux2_1 _2752_ (.A0(\tms1x00.RAM[70][3] ),
    .A1(\tms1x00.RAM[71][3] ),
    .S(_0823_),
    .X(_1142_));
 sky130_fd_sc_hd__and2_1 _2753_ (.A(_0822_),
    .B(_1142_),
    .X(_1143_));
 sky130_fd_sc_hd__mux2_1 _2754_ (.A0(\tms1x00.RAM[68][3] ),
    .A1(\tms1x00.RAM[69][3] ),
    .S(_0826_),
    .X(_1144_));
 sky130_fd_sc_hd__a21o_1 _2755_ (.A1(_0786_),
    .A2(_1144_),
    .B1(_0828_),
    .X(_1145_));
 sky130_fd_sc_hd__mux4_1 _2756_ (.A0(\tms1x00.RAM[64][3] ),
    .A1(\tms1x00.RAM[65][3] ),
    .A2(\tms1x00.RAM[66][3] ),
    .A3(\tms1x00.RAM[67][3] ),
    .S0(_0830_),
    .S1(_0831_),
    .X(_1146_));
 sky130_fd_sc_hd__o221a_1 _2757_ (.A1(_1143_),
    .A2(_1145_),
    .B1(_1146_),
    .B2(_0807_),
    .C1(_0775_),
    .X(_1147_));
 sky130_fd_sc_hd__mux4_1 _2758_ (.A0(\tms1x00.RAM[72][3] ),
    .A1(\tms1x00.RAM[73][3] ),
    .A2(\tms1x00.RAM[74][3] ),
    .A3(\tms1x00.RAM[75][3] ),
    .S0(_0799_),
    .S1(_0813_),
    .X(_1148_));
 sky130_fd_sc_hd__or2b_1 _2759_ (.A(\tms1x00.RAM[79][3] ),
    .B_N(_0778_),
    .X(_1149_));
 sky130_fd_sc_hd__o21a_1 _2760_ (.A1(_0778_),
    .A2(\tms1x00.RAM[78][3] ),
    .B1(_0812_),
    .X(_1150_));
 sky130_fd_sc_hd__mux2_1 _2761_ (.A0(\tms1x00.RAM[76][3] ),
    .A1(\tms1x00.RAM[77][3] ),
    .S(_0826_),
    .X(_1151_));
 sky130_fd_sc_hd__a221o_1 _2762_ (.A1(_1149_),
    .A2(_1150_),
    .B1(_1151_),
    .B2(_0786_),
    .C1(_0828_),
    .X(_1152_));
 sky130_fd_sc_hd__o211a_1 _2763_ (.A1(_0798_),
    .A2(_1148_),
    .B1(_1152_),
    .C1(_0802_),
    .X(_1153_));
 sky130_fd_sc_hd__or3_1 _2764_ (.A(_0821_),
    .B(_1147_),
    .C(_1153_),
    .X(_1154_));
 sky130_fd_sc_hd__o311a_1 _2765_ (.A1(_0920_),
    .A2(_1135_),
    .A3(_1141_),
    .B1(_1154_),
    .C1(_0773_),
    .X(_1155_));
 sky130_fd_sc_hd__mux4_1 _2766_ (.A0(\tms1x00.RAM[108][3] ),
    .A1(\tms1x00.RAM[109][3] ),
    .A2(\tms1x00.RAM[110][3] ),
    .A3(\tms1x00.RAM[111][3] ),
    .S0(_0931_),
    .S1(_0932_),
    .X(_1156_));
 sky130_fd_sc_hd__mux4_1 _2767_ (.A0(\tms1x00.RAM[104][3] ),
    .A1(\tms1x00.RAM[105][3] ),
    .A2(\tms1x00.RAM[106][3] ),
    .A3(\tms1x00.RAM[107][3] ),
    .S0(_0840_),
    .S1(_0813_),
    .X(_1157_));
 sky130_fd_sc_hd__or2_1 _2768_ (.A(_0798_),
    .B(_1157_),
    .X(_1158_));
 sky130_fd_sc_hd__o211a_1 _2769_ (.A1(_0940_),
    .A2(_1156_),
    .B1(_1158_),
    .C1(_0942_),
    .X(_1159_));
 sky130_fd_sc_hd__mux4_2 _2770_ (.A0(\tms1x00.RAM[96][3] ),
    .A1(\tms1x00.RAM[97][3] ),
    .A2(\tms1x00.RAM[98][3] ),
    .A3(\tms1x00.RAM[99][3] ),
    .S0(_0931_),
    .S1(_0932_),
    .X(_1160_));
 sky130_fd_sc_hd__mux4_1 _2771_ (.A0(\tms1x00.RAM[100][3] ),
    .A1(\tms1x00.RAM[101][3] ),
    .A2(\tms1x00.RAM[102][3] ),
    .A3(\tms1x00.RAM[103][3] ),
    .S0(_0873_),
    .S1(_0977_),
    .X(_1161_));
 sky130_fd_sc_hd__or2_1 _2772_ (.A(_0996_),
    .B(_1161_),
    .X(_1162_));
 sky130_fd_sc_hd__o211a_1 _2773_ (.A1(_0922_),
    .A2(_1160_),
    .B1(_1162_),
    .C1(_0944_),
    .X(_1163_));
 sky130_fd_sc_hd__or2b_1 _2774_ (.A(\tms1x00.RAM[119][3] ),
    .B_N(_0955_),
    .X(_1164_));
 sky130_fd_sc_hd__o21a_1 _2775_ (.A1(_0955_),
    .A2(\tms1x00.RAM[118][3] ),
    .B1(_0927_),
    .X(_1165_));
 sky130_fd_sc_hd__mux2_1 _2776_ (.A0(\tms1x00.RAM[116][3] ),
    .A1(\tms1x00.RAM[117][3] ),
    .S(_0789_),
    .X(_1166_));
 sky130_fd_sc_hd__a221o_1 _2777_ (.A1(_1164_),
    .A2(_1165_),
    .B1(_1166_),
    .B2(_0787_),
    .C1(_0996_),
    .X(_1167_));
 sky130_fd_sc_hd__mux4_1 _2778_ (.A0(\tms1x00.RAM[112][3] ),
    .A1(\tms1x00.RAM[113][3] ),
    .A2(\tms1x00.RAM[114][3] ),
    .A3(\tms1x00.RAM[115][3] ),
    .S0(_0873_),
    .S1(_0977_),
    .X(_1168_));
 sky130_fd_sc_hd__or2_1 _2779_ (.A(_0921_),
    .B(_1168_),
    .X(_1169_));
 sky130_fd_sc_hd__mux4_1 _2780_ (.A0(\tms1x00.RAM[124][3] ),
    .A1(\tms1x00.RAM[125][3] ),
    .A2(\tms1x00.RAM[126][3] ),
    .A3(\tms1x00.RAM[127][3] ),
    .S0(_0923_),
    .S1(_0927_),
    .X(_1170_));
 sky130_fd_sc_hd__mux4_1 _2781_ (.A0(\tms1x00.RAM[120][3] ),
    .A1(\tms1x00.RAM[121][3] ),
    .A2(\tms1x00.RAM[122][3] ),
    .A3(\tms1x00.RAM[123][3] ),
    .S0(_0823_),
    .S1(_0850_),
    .X(_1171_));
 sky130_fd_sc_hd__or2_1 _2782_ (.A(_0783_),
    .B(_1171_),
    .X(_1172_));
 sky130_fd_sc_hd__o211a_1 _2783_ (.A1(_0940_),
    .A2(_1170_),
    .B1(_1172_),
    .C1(_0806_),
    .X(_1173_));
 sky130_fd_sc_hd__a311o_1 _2784_ (.A1(_0944_),
    .A2(_1167_),
    .A3(_1169_),
    .B1(_0804_),
    .C1(_1173_),
    .X(_1174_));
 sky130_fd_sc_hd__o311a_1 _2785_ (.A1(_0821_),
    .A2(_1159_),
    .A3(_1163_),
    .B1(_0040_),
    .C1(_1174_),
    .X(_1175_));
 sky130_fd_sc_hd__mux4_1 _2786_ (.A0(\tms1x00.RAM[16][3] ),
    .A1(\tms1x00.RAM[17][3] ),
    .A2(\tms1x00.RAM[18][3] ),
    .A3(\tms1x00.RAM[19][3] ),
    .S0(_0924_),
    .S1(_0928_),
    .X(_1176_));
 sky130_fd_sc_hd__mux4_2 _2787_ (.A0(\tms1x00.RAM[20][3] ),
    .A1(\tms1x00.RAM[21][3] ),
    .A2(\tms1x00.RAM[22][3] ),
    .A3(\tms1x00.RAM[23][3] ),
    .S0(_0923_),
    .S1(_0927_),
    .X(_1177_));
 sky130_fd_sc_hd__or2_1 _2788_ (.A(_0996_),
    .B(_1177_),
    .X(_1178_));
 sky130_fd_sc_hd__o211a_1 _2789_ (.A1(_0922_),
    .A2(_1176_),
    .B1(_1178_),
    .C1(_0944_),
    .X(_1179_));
 sky130_fd_sc_hd__mux2_1 _2790_ (.A0(\tms1x00.RAM[30][3] ),
    .A1(\tms1x00.RAM[31][3] ),
    .S(_0945_),
    .X(_1180_));
 sky130_fd_sc_hd__and2_1 _2791_ (.A(_0928_),
    .B(_1180_),
    .X(_1181_));
 sky130_fd_sc_hd__mux2_1 _2792_ (.A0(\tms1x00.RAM[28][3] ),
    .A1(\tms1x00.RAM[29][3] ),
    .S(_0945_),
    .X(_1182_));
 sky130_fd_sc_hd__a21o_1 _2793_ (.A1(_0787_),
    .A2(_1182_),
    .B1(_0940_),
    .X(_1183_));
 sky130_fd_sc_hd__mux4_2 _2794_ (.A0(\tms1x00.RAM[24][3] ),
    .A1(\tms1x00.RAM[25][3] ),
    .A2(\tms1x00.RAM[26][3] ),
    .A3(\tms1x00.RAM[27][3] ),
    .S0(_0924_),
    .S1(_0928_),
    .X(_1184_));
 sky130_fd_sc_hd__o221a_1 _2795_ (.A1(_1181_),
    .A2(_1183_),
    .B1(_1184_),
    .B2(_0922_),
    .C1(_0942_),
    .X(_1185_));
 sky130_fd_sc_hd__mux2_1 _2796_ (.A0(\tms1x00.RAM[6][3] ),
    .A1(\tms1x00.RAM[7][3] ),
    .S(_0788_),
    .X(_1186_));
 sky130_fd_sc_hd__and2_1 _2797_ (.A(_0927_),
    .B(_1186_),
    .X(_1187_));
 sky130_fd_sc_hd__mux2_1 _2798_ (.A0(\tms1x00.RAM[4][3] ),
    .A1(\tms1x00.RAM[5][3] ),
    .S(_0778_),
    .X(_1188_));
 sky130_fd_sc_hd__a21o_1 _2799_ (.A1(_0818_),
    .A2(_1188_),
    .B1(_0794_),
    .X(_1189_));
 sky130_fd_sc_hd__mux4_2 _2800_ (.A0(\tms1x00.RAM[0][3] ),
    .A1(\tms1x00.RAM[1][3] ),
    .A2(\tms1x00.RAM[2][3] ),
    .A3(\tms1x00.RAM[3][3] ),
    .S0(_0816_),
    .S1(_0977_),
    .X(_1190_));
 sky130_fd_sc_hd__o221a_1 _2801_ (.A1(_1187_),
    .A2(_1189_),
    .B1(_1190_),
    .B2(_0921_),
    .C1(_0775_),
    .X(_1191_));
 sky130_fd_sc_hd__mux4_1 _2802_ (.A0(\tms1x00.RAM[8][3] ),
    .A1(\tms1x00.RAM[9][3] ),
    .A2(\tms1x00.RAM[10][3] ),
    .A3(\tms1x00.RAM[11][3] ),
    .S0(_0816_),
    .S1(_0927_),
    .X(_1192_));
 sky130_fd_sc_hd__or2b_1 _2803_ (.A(\tms1x00.RAM[15][3] ),
    .B_N(_0840_),
    .X(_1193_));
 sky130_fd_sc_hd__o21a_1 _2804_ (.A1(_0840_),
    .A2(\tms1x00.RAM[14][3] ),
    .B1(_0780_),
    .X(_1194_));
 sky130_fd_sc_hd__mux2_1 _2805_ (.A0(\tms1x00.RAM[12][3] ),
    .A1(\tms1x00.RAM[13][3] ),
    .S(_0778_),
    .X(_1195_));
 sky130_fd_sc_hd__a221o_1 _2806_ (.A1(_1193_),
    .A2(_1194_),
    .B1(_1195_),
    .B2(_0786_),
    .C1(_0794_),
    .X(_1196_));
 sky130_fd_sc_hd__o211a_1 _2807_ (.A1(_0921_),
    .A2(_1192_),
    .B1(_1196_),
    .C1(_0806_),
    .X(_1197_));
 sky130_fd_sc_hd__or3_1 _2808_ (.A(_0821_),
    .B(_1191_),
    .C(_1197_),
    .X(_1198_));
 sky130_fd_sc_hd__o311a_1 _2809_ (.A1(_0920_),
    .A2(_1179_),
    .A3(_1185_),
    .B1(_1198_),
    .C1(_0773_),
    .X(_1199_));
 sky130_fd_sc_hd__mux4_1 _2810_ (.A0(\tms1x00.RAM[36][3] ),
    .A1(\tms1x00.RAM[37][3] ),
    .A2(\tms1x00.RAM[38][3] ),
    .A3(\tms1x00.RAM[39][3] ),
    .S0(_0816_),
    .S1(_0927_),
    .X(_1200_));
 sky130_fd_sc_hd__or2_1 _2811_ (.A(_0996_),
    .B(_1200_),
    .X(_1201_));
 sky130_fd_sc_hd__mux4_2 _2812_ (.A0(\tms1x00.RAM[32][3] ),
    .A1(\tms1x00.RAM[33][3] ),
    .A2(\tms1x00.RAM[34][3] ),
    .A3(\tms1x00.RAM[35][3] ),
    .S0(_0816_),
    .S1(_0927_),
    .X(_1202_));
 sky130_fd_sc_hd__or2_1 _2813_ (.A(_0921_),
    .B(_1202_),
    .X(_1203_));
 sky130_fd_sc_hd__mux4_2 _2814_ (.A0(\tms1x00.RAM[44][3] ),
    .A1(\tms1x00.RAM[45][3] ),
    .A2(\tms1x00.RAM[46][3] ),
    .A3(\tms1x00.RAM[47][3] ),
    .S0(_0923_),
    .S1(_0791_),
    .X(_1204_));
 sky130_fd_sc_hd__mux4_1 _2815_ (.A0(\tms1x00.RAM[40][3] ),
    .A1(\tms1x00.RAM[41][3] ),
    .A2(\tms1x00.RAM[42][3] ),
    .A3(\tms1x00.RAM[43][3] ),
    .S0(_0826_),
    .S1(_0780_),
    .X(_1205_));
 sky130_fd_sc_hd__or2_1 _2816_ (.A(_0783_),
    .B(_1205_),
    .X(_1206_));
 sky130_fd_sc_hd__o211a_1 _2817_ (.A1(_0940_),
    .A2(_1204_),
    .B1(_1206_),
    .C1(_0806_),
    .X(_1207_));
 sky130_fd_sc_hd__a311o_1 _2818_ (.A1(_0944_),
    .A2(_1201_),
    .A3(_1203_),
    .B1(_0821_),
    .C1(_1207_),
    .X(_1208_));
 sky130_fd_sc_hd__or2b_1 _2819_ (.A(\tms1x00.RAM[55][3] ),
    .B_N(_0931_),
    .X(_1209_));
 sky130_fd_sc_hd__o21a_1 _2820_ (.A1(_0931_),
    .A2(\tms1x00.RAM[54][3] ),
    .B1(_0791_),
    .X(_1210_));
 sky130_fd_sc_hd__mux2_1 _2821_ (.A0(\tms1x00.RAM[52][3] ),
    .A1(\tms1x00.RAM[53][3] ),
    .S(_0975_),
    .X(_1211_));
 sky130_fd_sc_hd__a221o_1 _2822_ (.A1(_1209_),
    .A2(_1210_),
    .B1(_1211_),
    .B2(_0787_),
    .C1(_0996_),
    .X(_1212_));
 sky130_fd_sc_hd__mux4_2 _2823_ (.A0(\tms1x00.RAM[48][3] ),
    .A1(\tms1x00.RAM[49][3] ),
    .A2(\tms1x00.RAM[50][3] ),
    .A3(\tms1x00.RAM[51][3] ),
    .S0(_0816_),
    .S1(_0977_),
    .X(_1213_));
 sky130_fd_sc_hd__or2_1 _2824_ (.A(_0921_),
    .B(_1213_),
    .X(_1214_));
 sky130_fd_sc_hd__mux4_1 _2825_ (.A0(\tms1x00.RAM[60][3] ),
    .A1(\tms1x00.RAM[61][3] ),
    .A2(\tms1x00.RAM[62][3] ),
    .A3(\tms1x00.RAM[63][3] ),
    .S0(_0923_),
    .S1(_0927_),
    .X(_1215_));
 sky130_fd_sc_hd__mux4_1 _2826_ (.A0(\tms1x00.RAM[56][3] ),
    .A1(\tms1x00.RAM[57][3] ),
    .A2(\tms1x00.RAM[58][3] ),
    .A3(\tms1x00.RAM[59][3] ),
    .S0(_0826_),
    .S1(_0850_),
    .X(_1216_));
 sky130_fd_sc_hd__or2_1 _2827_ (.A(_0783_),
    .B(_1216_),
    .X(_1217_));
 sky130_fd_sc_hd__o211a_1 _2828_ (.A1(_0940_),
    .A2(_1215_),
    .B1(_1217_),
    .C1(_0806_),
    .X(_1218_));
 sky130_fd_sc_hd__a311o_1 _2829_ (.A1(_0944_),
    .A2(_1212_),
    .A3(_1214_),
    .B1(_0920_),
    .C1(_1218_),
    .X(_1219_));
 sky130_fd_sc_hd__a31o_1 _2830_ (.A1(_0040_),
    .A2(_1208_),
    .A3(_1219_),
    .B1(_0041_),
    .X(_1220_));
 sky130_fd_sc_hd__o32a_2 _2831_ (.A1(_0835_),
    .A2(_1155_),
    .A3(_1175_),
    .B1(_1199_),
    .B2(_1220_),
    .X(_1221_));
 sky130_fd_sc_hd__nand2_1 _2832_ (.A(_0747_),
    .B(_0748_),
    .Y(_1222_));
 sky130_fd_sc_hd__a22o_1 _2833_ (.A1(\tms1x00.A[3] ),
    .A2(_0909_),
    .B1(_1221_),
    .B2(_1222_),
    .X(_1223_));
 sky130_fd_sc_hd__clkbuf_4 _2834_ (.A(_1223_),
    .X(_1224_));
 sky130_fd_sc_hd__clkbuf_4 _2835_ (.A(_1224_),
    .X(_1225_));
 sky130_fd_sc_hd__mux2_1 _2836_ (.A0(_1225_),
    .A1(\tms1x00.RAM[109][3] ),
    .S(_0918_),
    .X(_1226_));
 sky130_fd_sc_hd__clkbuf_1 _2837_ (.A(_1226_),
    .X(_0054_));
 sky130_fd_sc_hd__nand2_1 _2838_ (.A(\tms1x00.ram_addr_buff[0] ),
    .B(\tms1x00.ram_addr_buff[1] ),
    .Y(_1227_));
 sky130_fd_sc_hd__or3_1 _2839_ (.A(\tms1x00.ram_addr_buff[2] ),
    .B(\tms1x00.ram_addr_buff[3] ),
    .C(_0915_),
    .X(_1228_));
 sky130_fd_sc_hd__or2_4 _2840_ (.A(_1227_),
    .B(_1228_),
    .X(_1229_));
 sky130_fd_sc_hd__or2_2 _2841_ (.A(_0914_),
    .B(_1229_),
    .X(_1230_));
 sky130_fd_sc_hd__mux2_1 _2842_ (.A0(_0912_),
    .A1(\tms1x00.RAM[99][0] ),
    .S(_1230_),
    .X(_1231_));
 sky130_fd_sc_hd__clkbuf_1 _2843_ (.A(_1231_),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _2844_ (.A0(_1035_),
    .A1(\tms1x00.RAM[99][1] ),
    .S(_1230_),
    .X(_1232_));
 sky130_fd_sc_hd__clkbuf_1 _2845_ (.A(_1232_),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _2846_ (.A0(_1130_),
    .A1(\tms1x00.RAM[99][2] ),
    .S(_1230_),
    .X(_1233_));
 sky130_fd_sc_hd__clkbuf_1 _2847_ (.A(_1233_),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _2848_ (.A0(_1225_),
    .A1(\tms1x00.RAM[99][3] ),
    .S(_1230_),
    .X(_1234_));
 sky130_fd_sc_hd__clkbuf_1 _2849_ (.A(_1234_),
    .X(_0058_));
 sky130_fd_sc_hd__clkbuf_4 _2850_ (.A(_0911_),
    .X(_1235_));
 sky130_fd_sc_hd__or3b_4 _2851_ (.A(\tms1x00.ram_addr_buff[4] ),
    .B(\tms1x00.ram_addr_buff[5] ),
    .C_N(\tms1x00.ram_addr_buff[6] ),
    .X(_1236_));
 sky130_fd_sc_hd__buf_4 _2852_ (.A(_1236_),
    .X(_1237_));
 sky130_fd_sc_hd__or3b_1 _2853_ (.A(\tms1x00.ram_addr_buff[3] ),
    .B(_0915_),
    .C_N(\tms1x00.ram_addr_buff[2] ),
    .X(_1238_));
 sky130_fd_sc_hd__or3b_1 _2854_ (.A(\tms1x00.ram_addr_buff[1] ),
    .B(_1238_),
    .C_N(_0717_),
    .X(_1239_));
 sky130_fd_sc_hd__buf_4 _2855_ (.A(_1239_),
    .X(_1240_));
 sky130_fd_sc_hd__nor2_2 _2856_ (.A(_1237_),
    .B(_1240_),
    .Y(_1241_));
 sky130_fd_sc_hd__mux2_1 _2857_ (.A0(\tms1x00.RAM[69][0] ),
    .A1(_1235_),
    .S(_1241_),
    .X(_1242_));
 sky130_fd_sc_hd__clkbuf_1 _2858_ (.A(_1242_),
    .X(_0059_));
 sky130_fd_sc_hd__buf_4 _2859_ (.A(_1034_),
    .X(_1243_));
 sky130_fd_sc_hd__mux2_1 _2860_ (.A0(\tms1x00.RAM[69][1] ),
    .A1(_1243_),
    .S(_1241_),
    .X(_1244_));
 sky130_fd_sc_hd__clkbuf_1 _2861_ (.A(_1244_),
    .X(_0060_));
 sky130_fd_sc_hd__buf_4 _2862_ (.A(_1129_),
    .X(_1245_));
 sky130_fd_sc_hd__mux2_1 _2863_ (.A0(\tms1x00.RAM[69][2] ),
    .A1(_1245_),
    .S(_1241_),
    .X(_1246_));
 sky130_fd_sc_hd__clkbuf_1 _2864_ (.A(_1246_),
    .X(_0061_));
 sky130_fd_sc_hd__buf_4 _2865_ (.A(_1224_),
    .X(_1247_));
 sky130_fd_sc_hd__mux2_1 _2866_ (.A0(\tms1x00.RAM[69][3] ),
    .A1(_1247_),
    .S(_1241_),
    .X(_1248_));
 sky130_fd_sc_hd__clkbuf_1 _2867_ (.A(_1248_),
    .X(_0062_));
 sky130_fd_sc_hd__or3b_4 _2868_ (.A(\tms1x00.ram_addr_buff[5] ),
    .B(\tms1x00.ram_addr_buff[6] ),
    .C_N(\tms1x00.ram_addr_buff[4] ),
    .X(_1249_));
 sky130_fd_sc_hd__buf_4 _2869_ (.A(_1249_),
    .X(_1250_));
 sky130_fd_sc_hd__or3b_4 _2870_ (.A(_0728_),
    .B(_1228_),
    .C_N(_0717_),
    .X(_1251_));
 sky130_fd_sc_hd__or2_2 _2871_ (.A(_1250_),
    .B(_1251_),
    .X(_1252_));
 sky130_fd_sc_hd__mux2_1 _2872_ (.A0(_0912_),
    .A1(\tms1x00.RAM[17][0] ),
    .S(_1252_),
    .X(_1253_));
 sky130_fd_sc_hd__clkbuf_1 _2873_ (.A(_1253_),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _2874_ (.A0(_1035_),
    .A1(\tms1x00.RAM[17][1] ),
    .S(_1252_),
    .X(_1254_));
 sky130_fd_sc_hd__clkbuf_1 _2875_ (.A(_1254_),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _2876_ (.A0(_1130_),
    .A1(\tms1x00.RAM[17][2] ),
    .S(_1252_),
    .X(_1255_));
 sky130_fd_sc_hd__clkbuf_1 _2877_ (.A(_1255_),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _2878_ (.A0(_1225_),
    .A1(\tms1x00.RAM[17][3] ),
    .S(_1252_),
    .X(_1256_));
 sky130_fd_sc_hd__clkbuf_1 _2879_ (.A(_1256_),
    .X(_0066_));
 sky130_fd_sc_hd__nand3b_4 _2880_ (.A_N(\tms1x00.ram_addr_buff[5] ),
    .B(\tms1x00.ram_addr_buff[6] ),
    .C(\tms1x00.ram_addr_buff[4] ),
    .Y(_1257_));
 sky130_fd_sc_hd__buf_6 _2881_ (.A(_1257_),
    .X(_1258_));
 sky130_fd_sc_hd__or3b_1 _2882_ (.A(\tms1x00.ram_addr_buff[2] ),
    .B(_0915_),
    .C_N(\tms1x00.ram_addr_buff[3] ),
    .X(_1259_));
 sky130_fd_sc_hd__or3b_1 _2883_ (.A(\tms1x00.ram_addr_buff[1] ),
    .B(_1259_),
    .C_N(\tms1x00.ram_addr_buff[0] ),
    .X(_1260_));
 sky130_fd_sc_hd__buf_6 _2884_ (.A(_1260_),
    .X(_1261_));
 sky130_fd_sc_hd__nor2_2 _2885_ (.A(_1258_),
    .B(_1261_),
    .Y(_1262_));
 sky130_fd_sc_hd__mux2_1 _2886_ (.A0(\tms1x00.RAM[89][0] ),
    .A1(_1235_),
    .S(_1262_),
    .X(_1263_));
 sky130_fd_sc_hd__clkbuf_1 _2887_ (.A(_1263_),
    .X(_0067_));
 sky130_fd_sc_hd__mux2_1 _2888_ (.A0(\tms1x00.RAM[89][1] ),
    .A1(_1243_),
    .S(_1262_),
    .X(_1264_));
 sky130_fd_sc_hd__clkbuf_1 _2889_ (.A(_1264_),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _2890_ (.A0(\tms1x00.RAM[89][2] ),
    .A1(_1245_),
    .S(_1262_),
    .X(_1265_));
 sky130_fd_sc_hd__clkbuf_1 _2891_ (.A(_1265_),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_1 _2892_ (.A0(\tms1x00.RAM[89][3] ),
    .A1(_1247_),
    .S(_1262_),
    .X(_1266_));
 sky130_fd_sc_hd__clkbuf_1 _2893_ (.A(_1266_),
    .X(_0070_));
 sky130_fd_sc_hd__nand3_4 _2894_ (.A(_0717_),
    .B(_0728_),
    .C(_0916_),
    .Y(_1267_));
 sky130_fd_sc_hd__or2_2 _2895_ (.A(_1237_),
    .B(_1267_),
    .X(_1268_));
 sky130_fd_sc_hd__mux2_1 _2896_ (.A0(_0912_),
    .A1(\tms1x00.RAM[79][0] ),
    .S(_1268_),
    .X(_1269_));
 sky130_fd_sc_hd__clkbuf_1 _2897_ (.A(_1269_),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _2898_ (.A0(_1035_),
    .A1(\tms1x00.RAM[79][1] ),
    .S(_1268_),
    .X(_1270_));
 sky130_fd_sc_hd__clkbuf_1 _2899_ (.A(_1270_),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_1 _2900_ (.A0(_1130_),
    .A1(\tms1x00.RAM[79][2] ),
    .S(_1268_),
    .X(_1271_));
 sky130_fd_sc_hd__clkbuf_1 _2901_ (.A(_1271_),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _2902_ (.A0(_1225_),
    .A1(\tms1x00.RAM[79][3] ),
    .S(_1268_),
    .X(_1272_));
 sky130_fd_sc_hd__clkbuf_1 _2903_ (.A(_1272_),
    .X(_0074_));
 sky130_fd_sc_hd__or3b_4 _2904_ (.A(_1228_),
    .B(_0717_),
    .C_N(_0728_),
    .X(_1273_));
 sky130_fd_sc_hd__or2_2 _2905_ (.A(_1250_),
    .B(_1273_),
    .X(_1274_));
 sky130_fd_sc_hd__mux2_1 _2906_ (.A0(_0912_),
    .A1(\tms1x00.RAM[18][0] ),
    .S(_1274_),
    .X(_1275_));
 sky130_fd_sc_hd__clkbuf_1 _2907_ (.A(_1275_),
    .X(_0075_));
 sky130_fd_sc_hd__mux2_1 _2908_ (.A0(_1035_),
    .A1(\tms1x00.RAM[18][1] ),
    .S(_1274_),
    .X(_1276_));
 sky130_fd_sc_hd__clkbuf_1 _2909_ (.A(_1276_),
    .X(_0076_));
 sky130_fd_sc_hd__mux2_1 _2910_ (.A0(_1130_),
    .A1(\tms1x00.RAM[18][2] ),
    .S(_1274_),
    .X(_1277_));
 sky130_fd_sc_hd__clkbuf_1 _2911_ (.A(_1277_),
    .X(_0077_));
 sky130_fd_sc_hd__mux2_1 _2912_ (.A0(_1225_),
    .A1(\tms1x00.RAM[18][3] ),
    .S(_1274_),
    .X(_1278_));
 sky130_fd_sc_hd__clkbuf_1 _2913_ (.A(_1278_),
    .X(_0078_));
 sky130_fd_sc_hd__mux2_1 _2914_ (.A0(\K_override[0] ),
    .A1(net65),
    .S(_0715_),
    .X(_1279_));
 sky130_fd_sc_hd__clkbuf_1 _2915_ (.A(_1279_),
    .X(_0079_));
 sky130_fd_sc_hd__mux2_1 _2916_ (.A0(\K_override[1] ),
    .A1(net66),
    .S(_0715_),
    .X(_1280_));
 sky130_fd_sc_hd__clkbuf_1 _2917_ (.A(_1280_),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _2918_ (.A0(\K_override[2] ),
    .A1(net60),
    .S(_0715_),
    .X(_1281_));
 sky130_fd_sc_hd__clkbuf_1 _2919_ (.A(_1281_),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_1 _2920_ (.A0(\K_override[3] ),
    .A1(net61),
    .S(_0715_),
    .X(_1282_));
 sky130_fd_sc_hd__clkbuf_1 _2921_ (.A(_1282_),
    .X(_0082_));
 sky130_fd_sc_hd__nand3b_4 _2922_ (.A_N(\tms1x00.ram_addr_buff[6] ),
    .B(\tms1x00.ram_addr_buff[5] ),
    .C(\tms1x00.ram_addr_buff[4] ),
    .Y(_1283_));
 sky130_fd_sc_hd__clkbuf_8 _2923_ (.A(_1283_),
    .X(_1284_));
 sky130_fd_sc_hd__or2_1 _2924_ (.A(_1227_),
    .B(_1259_),
    .X(_1285_));
 sky130_fd_sc_hd__buf_6 _2925_ (.A(_1285_),
    .X(_1286_));
 sky130_fd_sc_hd__nor2_2 _2926_ (.A(_1284_),
    .B(_1286_),
    .Y(_1287_));
 sky130_fd_sc_hd__mux2_1 _2927_ (.A0(\tms1x00.RAM[59][0] ),
    .A1(_1235_),
    .S(_1287_),
    .X(_1288_));
 sky130_fd_sc_hd__clkbuf_1 _2928_ (.A(_1288_),
    .X(_0083_));
 sky130_fd_sc_hd__mux2_1 _2929_ (.A0(\tms1x00.RAM[59][1] ),
    .A1(_1243_),
    .S(_1287_),
    .X(_1289_));
 sky130_fd_sc_hd__clkbuf_1 _2930_ (.A(_1289_),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_1 _2931_ (.A0(\tms1x00.RAM[59][2] ),
    .A1(_1245_),
    .S(_1287_),
    .X(_1290_));
 sky130_fd_sc_hd__clkbuf_1 _2932_ (.A(_1290_),
    .X(_0085_));
 sky130_fd_sc_hd__mux2_1 _2933_ (.A0(\tms1x00.RAM[59][3] ),
    .A1(_1247_),
    .S(_1287_),
    .X(_1291_));
 sky130_fd_sc_hd__clkbuf_1 _2934_ (.A(_1291_),
    .X(_0086_));
 sky130_fd_sc_hd__or2_2 _2935_ (.A(_1251_),
    .B(_1283_),
    .X(_1292_));
 sky130_fd_sc_hd__mux2_1 _2936_ (.A0(_0912_),
    .A1(\tms1x00.RAM[49][0] ),
    .S(_1292_),
    .X(_1293_));
 sky130_fd_sc_hd__clkbuf_1 _2937_ (.A(_1293_),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_1 _2938_ (.A0(_1035_),
    .A1(\tms1x00.RAM[49][1] ),
    .S(_1292_),
    .X(_1294_));
 sky130_fd_sc_hd__clkbuf_1 _2939_ (.A(_1294_),
    .X(_0088_));
 sky130_fd_sc_hd__mux2_1 _2940_ (.A0(_1130_),
    .A1(\tms1x00.RAM[49][2] ),
    .S(_1292_),
    .X(_1295_));
 sky130_fd_sc_hd__clkbuf_1 _2941_ (.A(_1295_),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _2942_ (.A0(_1225_),
    .A1(\tms1x00.RAM[49][3] ),
    .S(_1292_),
    .X(_1296_));
 sky130_fd_sc_hd__clkbuf_1 _2943_ (.A(_1296_),
    .X(_0090_));
 sky130_fd_sc_hd__or2_2 _2944_ (.A(_1229_),
    .B(_1249_),
    .X(_1297_));
 sky130_fd_sc_hd__mux2_1 _2945_ (.A0(_0912_),
    .A1(\tms1x00.RAM[19][0] ),
    .S(_1297_),
    .X(_1298_));
 sky130_fd_sc_hd__clkbuf_1 _2946_ (.A(_1298_),
    .X(_0091_));
 sky130_fd_sc_hd__mux2_1 _2947_ (.A0(_1035_),
    .A1(\tms1x00.RAM[19][1] ),
    .S(_1297_),
    .X(_1299_));
 sky130_fd_sc_hd__clkbuf_1 _2948_ (.A(_1299_),
    .X(_0092_));
 sky130_fd_sc_hd__mux2_1 _2949_ (.A0(_1130_),
    .A1(\tms1x00.RAM[19][2] ),
    .S(_1297_),
    .X(_1300_));
 sky130_fd_sc_hd__clkbuf_1 _2950_ (.A(_1300_),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _2951_ (.A0(_1225_),
    .A1(\tms1x00.RAM[19][3] ),
    .S(_1297_),
    .X(_1301_));
 sky130_fd_sc_hd__clkbuf_1 _2952_ (.A(_1301_),
    .X(_0094_));
 sky130_fd_sc_hd__or3_1 _2953_ (.A(\tms1x00.ram_addr_buff[0] ),
    .B(\tms1x00.ram_addr_buff[1] ),
    .C(_1259_),
    .X(_1302_));
 sky130_fd_sc_hd__buf_6 _2954_ (.A(_1302_),
    .X(_1303_));
 sky130_fd_sc_hd__nor2_2 _2955_ (.A(_0914_),
    .B(_1303_),
    .Y(_1304_));
 sky130_fd_sc_hd__mux2_1 _2956_ (.A0(\tms1x00.RAM[104][0] ),
    .A1(_1235_),
    .S(_1304_),
    .X(_1305_));
 sky130_fd_sc_hd__clkbuf_1 _2957_ (.A(_1305_),
    .X(_0095_));
 sky130_fd_sc_hd__mux2_1 _2958_ (.A0(\tms1x00.RAM[104][1] ),
    .A1(_1243_),
    .S(_1304_),
    .X(_1306_));
 sky130_fd_sc_hd__clkbuf_1 _2959_ (.A(_1306_),
    .X(_0096_));
 sky130_fd_sc_hd__mux2_1 _2960_ (.A0(\tms1x00.RAM[104][2] ),
    .A1(_1245_),
    .S(_1304_),
    .X(_1307_));
 sky130_fd_sc_hd__clkbuf_1 _2961_ (.A(_1307_),
    .X(_0097_));
 sky130_fd_sc_hd__mux2_1 _2962_ (.A0(\tms1x00.RAM[104][3] ),
    .A1(_1247_),
    .S(_1304_),
    .X(_1308_));
 sky130_fd_sc_hd__clkbuf_1 _2963_ (.A(_1308_),
    .X(_0098_));
 sky130_fd_sc_hd__or2_1 _2964_ (.A(_1227_),
    .B(_1238_),
    .X(_1309_));
 sky130_fd_sc_hd__clkbuf_8 _2965_ (.A(_1309_),
    .X(_1310_));
 sky130_fd_sc_hd__nor2_2 _2966_ (.A(_0914_),
    .B(_1310_),
    .Y(_1311_));
 sky130_fd_sc_hd__mux2_1 _2967_ (.A0(\tms1x00.RAM[103][0] ),
    .A1(_1235_),
    .S(_1311_),
    .X(_1312_));
 sky130_fd_sc_hd__clkbuf_1 _2968_ (.A(_1312_),
    .X(_0099_));
 sky130_fd_sc_hd__mux2_1 _2969_ (.A0(\tms1x00.RAM[103][1] ),
    .A1(_1243_),
    .S(_1311_),
    .X(_1313_));
 sky130_fd_sc_hd__clkbuf_1 _2970_ (.A(_1313_),
    .X(_0100_));
 sky130_fd_sc_hd__mux2_1 _2971_ (.A0(\tms1x00.RAM[103][2] ),
    .A1(_1245_),
    .S(_1311_),
    .X(_1314_));
 sky130_fd_sc_hd__clkbuf_1 _2972_ (.A(_1314_),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _2973_ (.A0(\tms1x00.RAM[103][3] ),
    .A1(_1247_),
    .S(_1311_),
    .X(_1315_));
 sky130_fd_sc_hd__clkbuf_1 _2974_ (.A(_1315_),
    .X(_0102_));
 sky130_fd_sc_hd__or3b_1 _2975_ (.A(_1238_),
    .B(\tms1x00.ram_addr_buff[0] ),
    .C_N(_0728_),
    .X(_1316_));
 sky130_fd_sc_hd__buf_4 _2976_ (.A(_1316_),
    .X(_1317_));
 sky130_fd_sc_hd__nor2_2 _2977_ (.A(_0914_),
    .B(_1317_),
    .Y(_1318_));
 sky130_fd_sc_hd__mux2_1 _2978_ (.A0(\tms1x00.RAM[102][0] ),
    .A1(_1235_),
    .S(_1318_),
    .X(_1319_));
 sky130_fd_sc_hd__clkbuf_1 _2979_ (.A(_1319_),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _2980_ (.A0(\tms1x00.RAM[102][1] ),
    .A1(_1243_),
    .S(_1318_),
    .X(_1320_));
 sky130_fd_sc_hd__clkbuf_1 _2981_ (.A(_1320_),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _2982_ (.A0(\tms1x00.RAM[102][2] ),
    .A1(_1245_),
    .S(_1318_),
    .X(_1321_));
 sky130_fd_sc_hd__clkbuf_1 _2983_ (.A(_1321_),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _2984_ (.A0(\tms1x00.RAM[102][3] ),
    .A1(_1247_),
    .S(_1318_),
    .X(_1322_));
 sky130_fd_sc_hd__clkbuf_1 _2985_ (.A(_1322_),
    .X(_0106_));
 sky130_fd_sc_hd__clkbuf_4 _2986_ (.A(_0910_),
    .X(_1323_));
 sky130_fd_sc_hd__buf_2 _2987_ (.A(_1323_),
    .X(_1324_));
 sky130_fd_sc_hd__nor2_2 _2988_ (.A(_0914_),
    .B(_1240_),
    .Y(_1325_));
 sky130_fd_sc_hd__mux2_1 _2989_ (.A0(\tms1x00.RAM[101][0] ),
    .A1(_1324_),
    .S(_1325_),
    .X(_1326_));
 sky130_fd_sc_hd__clkbuf_1 _2990_ (.A(_1326_),
    .X(_0107_));
 sky130_fd_sc_hd__clkbuf_4 _2991_ (.A(_1033_),
    .X(_1327_));
 sky130_fd_sc_hd__buf_2 _2992_ (.A(_1327_),
    .X(_1328_));
 sky130_fd_sc_hd__mux2_1 _2993_ (.A0(\tms1x00.RAM[101][1] ),
    .A1(_1328_),
    .S(_1325_),
    .X(_1329_));
 sky130_fd_sc_hd__clkbuf_1 _2994_ (.A(_1329_),
    .X(_0108_));
 sky130_fd_sc_hd__clkbuf_4 _2995_ (.A(_1128_),
    .X(_1330_));
 sky130_fd_sc_hd__clkbuf_4 _2996_ (.A(_1330_),
    .X(_1331_));
 sky130_fd_sc_hd__mux2_1 _2997_ (.A0(\tms1x00.RAM[101][2] ),
    .A1(_1331_),
    .S(_1325_),
    .X(_1332_));
 sky130_fd_sc_hd__clkbuf_1 _2998_ (.A(_1332_),
    .X(_0109_));
 sky130_fd_sc_hd__clkbuf_4 _2999_ (.A(_1223_),
    .X(_1333_));
 sky130_fd_sc_hd__clkbuf_4 _3000_ (.A(_1333_),
    .X(_1334_));
 sky130_fd_sc_hd__mux2_1 _3001_ (.A0(\tms1x00.RAM[101][3] ),
    .A1(_1334_),
    .S(_1325_),
    .X(_1335_));
 sky130_fd_sc_hd__clkbuf_1 _3002_ (.A(_1335_),
    .X(_0110_));
 sky130_fd_sc_hd__or3_1 _3003_ (.A(\tms1x00.ram_addr_buff[0] ),
    .B(\tms1x00.ram_addr_buff[1] ),
    .C(_1238_),
    .X(_1336_));
 sky130_fd_sc_hd__clkbuf_8 _3004_ (.A(_1336_),
    .X(_1337_));
 sky130_fd_sc_hd__nor2_2 _3005_ (.A(_0914_),
    .B(_1337_),
    .Y(_1338_));
 sky130_fd_sc_hd__mux2_1 _3006_ (.A0(\tms1x00.RAM[100][0] ),
    .A1(_1324_),
    .S(_1338_),
    .X(_1339_));
 sky130_fd_sc_hd__clkbuf_1 _3007_ (.A(_1339_),
    .X(_0111_));
 sky130_fd_sc_hd__mux2_1 _3008_ (.A0(\tms1x00.RAM[100][1] ),
    .A1(_1328_),
    .S(_1338_),
    .X(_1340_));
 sky130_fd_sc_hd__clkbuf_1 _3009_ (.A(_1340_),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _3010_ (.A0(\tms1x00.RAM[100][2] ),
    .A1(_1331_),
    .S(_1338_),
    .X(_1341_));
 sky130_fd_sc_hd__clkbuf_1 _3011_ (.A(_1341_),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _3012_ (.A0(\tms1x00.RAM[100][3] ),
    .A1(_1334_),
    .S(_1338_),
    .X(_1342_));
 sky130_fd_sc_hd__clkbuf_1 _3013_ (.A(_1342_),
    .X(_0114_));
 sky130_fd_sc_hd__or3_4 _3014_ (.A(\tms1x00.ram_addr_buff[4] ),
    .B(\tms1x00.ram_addr_buff[5] ),
    .C(\tms1x00.ram_addr_buff[6] ),
    .X(_1343_));
 sky130_fd_sc_hd__buf_6 _3015_ (.A(_1343_),
    .X(_1344_));
 sky130_fd_sc_hd__or3_4 _3016_ (.A(_0717_),
    .B(_0728_),
    .C(_1228_),
    .X(_1345_));
 sky130_fd_sc_hd__or2_2 _3017_ (.A(_1344_),
    .B(_1345_),
    .X(_1346_));
 sky130_fd_sc_hd__mux2_1 _3018_ (.A0(_0912_),
    .A1(\tms1x00.RAM[0][0] ),
    .S(_1346_),
    .X(_1347_));
 sky130_fd_sc_hd__clkbuf_1 _3019_ (.A(_1347_),
    .X(_0115_));
 sky130_fd_sc_hd__mux2_1 _3020_ (.A0(_1035_),
    .A1(\tms1x00.RAM[0][1] ),
    .S(_1346_),
    .X(_1348_));
 sky130_fd_sc_hd__clkbuf_1 _3021_ (.A(_1348_),
    .X(_0116_));
 sky130_fd_sc_hd__mux2_1 _3022_ (.A0(_1130_),
    .A1(\tms1x00.RAM[0][2] ),
    .S(_1346_),
    .X(_1349_));
 sky130_fd_sc_hd__clkbuf_1 _3023_ (.A(_1349_),
    .X(_0117_));
 sky130_fd_sc_hd__mux2_1 _3024_ (.A0(_1225_),
    .A1(\tms1x00.RAM[0][3] ),
    .S(_1346_),
    .X(_1350_));
 sky130_fd_sc_hd__clkbuf_1 _3025_ (.A(_1350_),
    .X(_0118_));
 sky130_fd_sc_hd__or2_2 _3026_ (.A(_0913_),
    .B(_1273_),
    .X(_1351_));
 sky130_fd_sc_hd__mux2_1 _3027_ (.A0(_0912_),
    .A1(\tms1x00.RAM[98][0] ),
    .S(_1351_),
    .X(_1352_));
 sky130_fd_sc_hd__clkbuf_1 _3028_ (.A(_1352_),
    .X(_0119_));
 sky130_fd_sc_hd__mux2_1 _3029_ (.A0(_1035_),
    .A1(\tms1x00.RAM[98][1] ),
    .S(_1351_),
    .X(_1353_));
 sky130_fd_sc_hd__clkbuf_1 _3030_ (.A(_1353_),
    .X(_0120_));
 sky130_fd_sc_hd__mux2_1 _3031_ (.A0(_1130_),
    .A1(\tms1x00.RAM[98][2] ),
    .S(_1351_),
    .X(_1354_));
 sky130_fd_sc_hd__clkbuf_1 _3032_ (.A(_1354_),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _3033_ (.A0(_1225_),
    .A1(\tms1x00.RAM[98][3] ),
    .S(_1351_),
    .X(_1355_));
 sky130_fd_sc_hd__clkbuf_1 _3034_ (.A(_1355_),
    .X(_0122_));
 sky130_fd_sc_hd__or2_2 _3035_ (.A(_0913_),
    .B(_1251_),
    .X(_1356_));
 sky130_fd_sc_hd__mux2_1 _3036_ (.A0(_0912_),
    .A1(\tms1x00.RAM[97][0] ),
    .S(_1356_),
    .X(_1357_));
 sky130_fd_sc_hd__clkbuf_1 _3037_ (.A(_1357_),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _3038_ (.A0(_1035_),
    .A1(\tms1x00.RAM[97][1] ),
    .S(_1356_),
    .X(_1358_));
 sky130_fd_sc_hd__clkbuf_1 _3039_ (.A(_1358_),
    .X(_0124_));
 sky130_fd_sc_hd__mux2_1 _3040_ (.A0(_1130_),
    .A1(\tms1x00.RAM[97][2] ),
    .S(_1356_),
    .X(_1359_));
 sky130_fd_sc_hd__clkbuf_1 _3041_ (.A(_1359_),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_1 _3042_ (.A0(_1225_),
    .A1(\tms1x00.RAM[97][3] ),
    .S(_1356_),
    .X(_1360_));
 sky130_fd_sc_hd__clkbuf_1 _3043_ (.A(_1360_),
    .X(_0126_));
 sky130_fd_sc_hd__buf_2 _3044_ (.A(_0911_),
    .X(_1361_));
 sky130_fd_sc_hd__or2_2 _3045_ (.A(_0913_),
    .B(_1345_),
    .X(_1362_));
 sky130_fd_sc_hd__mux2_1 _3046_ (.A0(_1361_),
    .A1(\tms1x00.RAM[96][0] ),
    .S(_1362_),
    .X(_1363_));
 sky130_fd_sc_hd__clkbuf_1 _3047_ (.A(_1363_),
    .X(_0127_));
 sky130_fd_sc_hd__clkbuf_4 _3048_ (.A(_1034_),
    .X(_1364_));
 sky130_fd_sc_hd__mux2_1 _3049_ (.A0(_1364_),
    .A1(\tms1x00.RAM[96][1] ),
    .S(_1362_),
    .X(_1365_));
 sky130_fd_sc_hd__clkbuf_1 _3050_ (.A(_1365_),
    .X(_0128_));
 sky130_fd_sc_hd__clkbuf_4 _3051_ (.A(_1129_),
    .X(_1366_));
 sky130_fd_sc_hd__mux2_1 _3052_ (.A0(_1366_),
    .A1(\tms1x00.RAM[96][2] ),
    .S(_1362_),
    .X(_1367_));
 sky130_fd_sc_hd__clkbuf_1 _3053_ (.A(_1367_),
    .X(_0129_));
 sky130_fd_sc_hd__clkbuf_4 _3054_ (.A(_1224_),
    .X(_1368_));
 sky130_fd_sc_hd__mux2_1 _3055_ (.A0(_1368_),
    .A1(\tms1x00.RAM[96][3] ),
    .S(_1362_),
    .X(_1369_));
 sky130_fd_sc_hd__clkbuf_1 _3056_ (.A(_1369_),
    .X(_0130_));
 sky130_fd_sc_hd__or2_2 _3057_ (.A(_1258_),
    .B(_1267_),
    .X(_1370_));
 sky130_fd_sc_hd__mux2_1 _3058_ (.A0(_1361_),
    .A1(\tms1x00.RAM[95][0] ),
    .S(_1370_),
    .X(_1371_));
 sky130_fd_sc_hd__clkbuf_1 _3059_ (.A(_1371_),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_1 _3060_ (.A0(_1364_),
    .A1(\tms1x00.RAM[95][1] ),
    .S(_1370_),
    .X(_1372_));
 sky130_fd_sc_hd__clkbuf_1 _3061_ (.A(_1372_),
    .X(_0132_));
 sky130_fd_sc_hd__mux2_1 _3062_ (.A0(_1366_),
    .A1(\tms1x00.RAM[95][2] ),
    .S(_1370_),
    .X(_1373_));
 sky130_fd_sc_hd__clkbuf_1 _3063_ (.A(_1373_),
    .X(_0133_));
 sky130_fd_sc_hd__mux2_1 _3064_ (.A0(_1368_),
    .A1(\tms1x00.RAM[95][3] ),
    .S(_1370_),
    .X(_1374_));
 sky130_fd_sc_hd__clkbuf_1 _3065_ (.A(_1374_),
    .X(_0134_));
 sky130_fd_sc_hd__nand3_2 _3066_ (.A(\tms1x00.ram_addr_buff[4] ),
    .B(\tms1x00.ram_addr_buff[5] ),
    .C(\tms1x00.ram_addr_buff[6] ),
    .Y(_1375_));
 sky130_fd_sc_hd__or2_2 _3067_ (.A(_1273_),
    .B(_1375_),
    .X(_1376_));
 sky130_fd_sc_hd__mux2_1 _3068_ (.A0(_1361_),
    .A1(\tms1x00.RAM[114][0] ),
    .S(_1376_),
    .X(_1377_));
 sky130_fd_sc_hd__clkbuf_1 _3069_ (.A(_1377_),
    .X(_0135_));
 sky130_fd_sc_hd__mux2_1 _3070_ (.A0(_1364_),
    .A1(\tms1x00.RAM[114][1] ),
    .S(_1376_),
    .X(_1378_));
 sky130_fd_sc_hd__clkbuf_1 _3071_ (.A(_1378_),
    .X(_0136_));
 sky130_fd_sc_hd__mux2_1 _3072_ (.A0(_1366_),
    .A1(\tms1x00.RAM[114][2] ),
    .S(_1376_),
    .X(_1379_));
 sky130_fd_sc_hd__clkbuf_1 _3073_ (.A(_1379_),
    .X(_0137_));
 sky130_fd_sc_hd__mux2_1 _3074_ (.A0(_1368_),
    .A1(\tms1x00.RAM[114][3] ),
    .S(_1376_),
    .X(_1380_));
 sky130_fd_sc_hd__clkbuf_1 _3075_ (.A(_1380_),
    .X(_0138_));
 sky130_fd_sc_hd__or2_2 _3076_ (.A(_1251_),
    .B(_1375_),
    .X(_1381_));
 sky130_fd_sc_hd__mux2_1 _3077_ (.A0(_1361_),
    .A1(\tms1x00.RAM[113][0] ),
    .S(_1381_),
    .X(_1382_));
 sky130_fd_sc_hd__clkbuf_1 _3078_ (.A(_1382_),
    .X(_0139_));
 sky130_fd_sc_hd__mux2_1 _3079_ (.A0(_1364_),
    .A1(\tms1x00.RAM[113][1] ),
    .S(_1381_),
    .X(_1383_));
 sky130_fd_sc_hd__clkbuf_1 _3080_ (.A(_1383_),
    .X(_0140_));
 sky130_fd_sc_hd__mux2_1 _3081_ (.A0(_1366_),
    .A1(\tms1x00.RAM[113][2] ),
    .S(_1381_),
    .X(_1384_));
 sky130_fd_sc_hd__clkbuf_1 _3082_ (.A(_1384_),
    .X(_0141_));
 sky130_fd_sc_hd__mux2_1 _3083_ (.A0(_1368_),
    .A1(\tms1x00.RAM[113][3] ),
    .S(_1381_),
    .X(_1385_));
 sky130_fd_sc_hd__clkbuf_1 _3084_ (.A(_1385_),
    .X(_0142_));
 sky130_fd_sc_hd__or2_2 _3085_ (.A(_1345_),
    .B(_1375_),
    .X(_1386_));
 sky130_fd_sc_hd__mux2_1 _3086_ (.A0(_1361_),
    .A1(\tms1x00.RAM[112][0] ),
    .S(_1386_),
    .X(_1387_));
 sky130_fd_sc_hd__clkbuf_1 _3087_ (.A(_1387_),
    .X(_0143_));
 sky130_fd_sc_hd__mux2_1 _3088_ (.A0(_1364_),
    .A1(\tms1x00.RAM[112][1] ),
    .S(_1386_),
    .X(_1388_));
 sky130_fd_sc_hd__clkbuf_1 _3089_ (.A(_1388_),
    .X(_0144_));
 sky130_fd_sc_hd__mux2_1 _3090_ (.A0(_1366_),
    .A1(\tms1x00.RAM[112][2] ),
    .S(_1386_),
    .X(_1389_));
 sky130_fd_sc_hd__clkbuf_1 _3091_ (.A(_1389_),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _3092_ (.A0(_1368_),
    .A1(\tms1x00.RAM[112][3] ),
    .S(_1386_),
    .X(_1390_));
 sky130_fd_sc_hd__clkbuf_1 _3093_ (.A(_1390_),
    .X(_0146_));
 sky130_fd_sc_hd__or2_2 _3094_ (.A(_0913_),
    .B(_1267_),
    .X(_1391_));
 sky130_fd_sc_hd__mux2_1 _3095_ (.A0(_1361_),
    .A1(\tms1x00.RAM[111][0] ),
    .S(_1391_),
    .X(_1392_));
 sky130_fd_sc_hd__clkbuf_1 _3096_ (.A(_1392_),
    .X(_0147_));
 sky130_fd_sc_hd__mux2_1 _3097_ (.A0(_1364_),
    .A1(\tms1x00.RAM[111][1] ),
    .S(_1391_),
    .X(_1393_));
 sky130_fd_sc_hd__clkbuf_1 _3098_ (.A(_1393_),
    .X(_0148_));
 sky130_fd_sc_hd__mux2_1 _3099_ (.A0(_1366_),
    .A1(\tms1x00.RAM[111][2] ),
    .S(_1391_),
    .X(_1394_));
 sky130_fd_sc_hd__clkbuf_1 _3100_ (.A(_1394_),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_1 _3101_ (.A0(_1368_),
    .A1(\tms1x00.RAM[111][3] ),
    .S(_1391_),
    .X(_1395_));
 sky130_fd_sc_hd__clkbuf_1 _3102_ (.A(_1395_),
    .X(_0150_));
 sky130_fd_sc_hd__nand3b_4 _3103_ (.A_N(_0717_),
    .B(_0728_),
    .C(_0916_),
    .Y(_1396_));
 sky130_fd_sc_hd__or2_2 _3104_ (.A(_0913_),
    .B(_1396_),
    .X(_1397_));
 sky130_fd_sc_hd__mux2_1 _3105_ (.A0(_1361_),
    .A1(\tms1x00.RAM[110][0] ),
    .S(_1397_),
    .X(_1398_));
 sky130_fd_sc_hd__clkbuf_1 _3106_ (.A(_1398_),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _3107_ (.A0(_1364_),
    .A1(\tms1x00.RAM[110][1] ),
    .S(_1397_),
    .X(_1399_));
 sky130_fd_sc_hd__clkbuf_1 _3108_ (.A(_1399_),
    .X(_0152_));
 sky130_fd_sc_hd__mux2_1 _3109_ (.A0(_1366_),
    .A1(\tms1x00.RAM[110][2] ),
    .S(_1397_),
    .X(_1400_));
 sky130_fd_sc_hd__clkbuf_1 _3110_ (.A(_1400_),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _3111_ (.A0(_1368_),
    .A1(\tms1x00.RAM[110][3] ),
    .S(_1397_),
    .X(_1401_));
 sky130_fd_sc_hd__clkbuf_1 _3112_ (.A(_1401_),
    .X(_0154_));
 sky130_fd_sc_hd__or3b_1 _3113_ (.A(_1259_),
    .B(\tms1x00.ram_addr_buff[0] ),
    .C_N(\tms1x00.ram_addr_buff[1] ),
    .X(_1402_));
 sky130_fd_sc_hd__buf_6 _3114_ (.A(_1402_),
    .X(_1403_));
 sky130_fd_sc_hd__nor2_2 _3115_ (.A(_1344_),
    .B(_1403_),
    .Y(_1404_));
 sky130_fd_sc_hd__mux2_1 _3116_ (.A0(\tms1x00.RAM[10][0] ),
    .A1(_1324_),
    .S(_1404_),
    .X(_1405_));
 sky130_fd_sc_hd__clkbuf_1 _3117_ (.A(_1405_),
    .X(_0155_));
 sky130_fd_sc_hd__mux2_1 _3118_ (.A0(\tms1x00.RAM[10][1] ),
    .A1(_1328_),
    .S(_1404_),
    .X(_1406_));
 sky130_fd_sc_hd__clkbuf_1 _3119_ (.A(_1406_),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _3120_ (.A0(\tms1x00.RAM[10][2] ),
    .A1(_1331_),
    .S(_1404_),
    .X(_1407_));
 sky130_fd_sc_hd__clkbuf_1 _3121_ (.A(_1407_),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_1 _3122_ (.A0(\tms1x00.RAM[10][3] ),
    .A1(_1334_),
    .S(_1404_),
    .X(_1408_));
 sky130_fd_sc_hd__clkbuf_1 _3123_ (.A(_1408_),
    .X(_0158_));
 sky130_fd_sc_hd__or3b_4 _3124_ (.A(_0717_),
    .B(_0728_),
    .C_N(_0916_),
    .X(_1409_));
 sky130_fd_sc_hd__or2_2 _3125_ (.A(_0913_),
    .B(_1409_),
    .X(_1410_));
 sky130_fd_sc_hd__mux2_1 _3126_ (.A0(_1361_),
    .A1(\tms1x00.RAM[108][0] ),
    .S(_1410_),
    .X(_1411_));
 sky130_fd_sc_hd__clkbuf_1 _3127_ (.A(_1411_),
    .X(_0159_));
 sky130_fd_sc_hd__mux2_1 _3128_ (.A0(_1364_),
    .A1(\tms1x00.RAM[108][1] ),
    .S(_1410_),
    .X(_1412_));
 sky130_fd_sc_hd__clkbuf_1 _3129_ (.A(_1412_),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _3130_ (.A0(_1366_),
    .A1(\tms1x00.RAM[108][2] ),
    .S(_1410_),
    .X(_1413_));
 sky130_fd_sc_hd__clkbuf_1 _3131_ (.A(_1413_),
    .X(_0161_));
 sky130_fd_sc_hd__mux2_1 _3132_ (.A0(_1368_),
    .A1(\tms1x00.RAM[108][3] ),
    .S(_1410_),
    .X(_1414_));
 sky130_fd_sc_hd__clkbuf_1 _3133_ (.A(_1414_),
    .X(_0162_));
 sky130_fd_sc_hd__nor2_2 _3134_ (.A(_0914_),
    .B(_1286_),
    .Y(_1415_));
 sky130_fd_sc_hd__mux2_1 _3135_ (.A0(\tms1x00.RAM[107][0] ),
    .A1(_1324_),
    .S(_1415_),
    .X(_1416_));
 sky130_fd_sc_hd__clkbuf_1 _3136_ (.A(_1416_),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _3137_ (.A0(\tms1x00.RAM[107][1] ),
    .A1(_1328_),
    .S(_1415_),
    .X(_1417_));
 sky130_fd_sc_hd__clkbuf_1 _3138_ (.A(_1417_),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_1 _3139_ (.A0(\tms1x00.RAM[107][2] ),
    .A1(_1331_),
    .S(_1415_),
    .X(_1418_));
 sky130_fd_sc_hd__clkbuf_1 _3140_ (.A(_1418_),
    .X(_0165_));
 sky130_fd_sc_hd__mux2_1 _3141_ (.A0(\tms1x00.RAM[107][3] ),
    .A1(_1334_),
    .S(_1415_),
    .X(_1419_));
 sky130_fd_sc_hd__clkbuf_1 _3142_ (.A(_1419_),
    .X(_0166_));
 sky130_fd_sc_hd__nor2_2 _3143_ (.A(_0914_),
    .B(_1403_),
    .Y(_1420_));
 sky130_fd_sc_hd__mux2_1 _3144_ (.A0(\tms1x00.RAM[106][0] ),
    .A1(_1324_),
    .S(_1420_),
    .X(_1421_));
 sky130_fd_sc_hd__clkbuf_1 _3145_ (.A(_1421_),
    .X(_0167_));
 sky130_fd_sc_hd__mux2_1 _3146_ (.A0(\tms1x00.RAM[106][1] ),
    .A1(_1328_),
    .S(_1420_),
    .X(_1422_));
 sky130_fd_sc_hd__clkbuf_1 _3147_ (.A(_1422_),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _3148_ (.A0(\tms1x00.RAM[106][2] ),
    .A1(_1331_),
    .S(_1420_),
    .X(_1423_));
 sky130_fd_sc_hd__clkbuf_1 _3149_ (.A(_1423_),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_1 _3150_ (.A0(\tms1x00.RAM[106][3] ),
    .A1(_1334_),
    .S(_1420_),
    .X(_1424_));
 sky130_fd_sc_hd__clkbuf_1 _3151_ (.A(_1424_),
    .X(_0170_));
 sky130_fd_sc_hd__nor2_2 _3152_ (.A(_0914_),
    .B(_1261_),
    .Y(_1425_));
 sky130_fd_sc_hd__mux2_1 _3153_ (.A0(\tms1x00.RAM[105][0] ),
    .A1(_1324_),
    .S(_1425_),
    .X(_1426_));
 sky130_fd_sc_hd__clkbuf_1 _3154_ (.A(_1426_),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _3155_ (.A0(\tms1x00.RAM[105][1] ),
    .A1(_1328_),
    .S(_1425_),
    .X(_1427_));
 sky130_fd_sc_hd__clkbuf_1 _3156_ (.A(_1427_),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_1 _3157_ (.A0(\tms1x00.RAM[105][2] ),
    .A1(_1331_),
    .S(_1425_),
    .X(_1428_));
 sky130_fd_sc_hd__clkbuf_1 _3158_ (.A(_1428_),
    .X(_0173_));
 sky130_fd_sc_hd__mux2_1 _3159_ (.A0(\tms1x00.RAM[105][3] ),
    .A1(_1334_),
    .S(_1425_),
    .X(_1429_));
 sky130_fd_sc_hd__clkbuf_1 _3160_ (.A(_1429_),
    .X(_0174_));
 sky130_fd_sc_hd__clkbuf_8 _3161_ (.A(_1375_),
    .X(_1430_));
 sky130_fd_sc_hd__or2_2 _3162_ (.A(_1430_),
    .B(_1409_),
    .X(_1431_));
 sky130_fd_sc_hd__mux2_1 _3163_ (.A0(_1361_),
    .A1(\tms1x00.RAM[124][0] ),
    .S(_1431_),
    .X(_1432_));
 sky130_fd_sc_hd__clkbuf_1 _3164_ (.A(_1432_),
    .X(_0175_));
 sky130_fd_sc_hd__mux2_1 _3165_ (.A0(_1364_),
    .A1(\tms1x00.RAM[124][1] ),
    .S(_1431_),
    .X(_1433_));
 sky130_fd_sc_hd__clkbuf_1 _3166_ (.A(_1433_),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _3167_ (.A0(_1366_),
    .A1(\tms1x00.RAM[124][2] ),
    .S(_1431_),
    .X(_1434_));
 sky130_fd_sc_hd__clkbuf_1 _3168_ (.A(_1434_),
    .X(_0177_));
 sky130_fd_sc_hd__mux2_1 _3169_ (.A0(_1368_),
    .A1(\tms1x00.RAM[124][3] ),
    .S(_1431_),
    .X(_1435_));
 sky130_fd_sc_hd__clkbuf_1 _3170_ (.A(_1435_),
    .X(_0178_));
 sky130_fd_sc_hd__nor2_2 _3171_ (.A(_1286_),
    .B(_1430_),
    .Y(_1436_));
 sky130_fd_sc_hd__mux2_1 _3172_ (.A0(\tms1x00.RAM[123][0] ),
    .A1(_1324_),
    .S(_1436_),
    .X(_1437_));
 sky130_fd_sc_hd__clkbuf_1 _3173_ (.A(_1437_),
    .X(_0179_));
 sky130_fd_sc_hd__mux2_1 _3174_ (.A0(\tms1x00.RAM[123][1] ),
    .A1(_1328_),
    .S(_1436_),
    .X(_1438_));
 sky130_fd_sc_hd__clkbuf_1 _3175_ (.A(_1438_),
    .X(_0180_));
 sky130_fd_sc_hd__mux2_1 _3176_ (.A0(\tms1x00.RAM[123][2] ),
    .A1(_1331_),
    .S(_1436_),
    .X(_1439_));
 sky130_fd_sc_hd__clkbuf_1 _3177_ (.A(_1439_),
    .X(_0181_));
 sky130_fd_sc_hd__mux2_1 _3178_ (.A0(\tms1x00.RAM[123][3] ),
    .A1(_1334_),
    .S(_1436_),
    .X(_1440_));
 sky130_fd_sc_hd__clkbuf_1 _3179_ (.A(_1440_),
    .X(_0182_));
 sky130_fd_sc_hd__nor2_2 _3180_ (.A(_1430_),
    .B(_1403_),
    .Y(_1441_));
 sky130_fd_sc_hd__mux2_1 _3181_ (.A0(\tms1x00.RAM[122][0] ),
    .A1(_1324_),
    .S(_1441_),
    .X(_1442_));
 sky130_fd_sc_hd__clkbuf_1 _3182_ (.A(_1442_),
    .X(_0183_));
 sky130_fd_sc_hd__mux2_1 _3183_ (.A0(\tms1x00.RAM[122][1] ),
    .A1(_1328_),
    .S(_1441_),
    .X(_1443_));
 sky130_fd_sc_hd__clkbuf_1 _3184_ (.A(_1443_),
    .X(_0184_));
 sky130_fd_sc_hd__mux2_1 _3185_ (.A0(\tms1x00.RAM[122][2] ),
    .A1(_1331_),
    .S(_1441_),
    .X(_1444_));
 sky130_fd_sc_hd__clkbuf_1 _3186_ (.A(_1444_),
    .X(_0185_));
 sky130_fd_sc_hd__mux2_1 _3187_ (.A0(\tms1x00.RAM[122][3] ),
    .A1(_1334_),
    .S(_1441_),
    .X(_1445_));
 sky130_fd_sc_hd__clkbuf_1 _3188_ (.A(_1445_),
    .X(_0186_));
 sky130_fd_sc_hd__nor2_2 _3189_ (.A(_1261_),
    .B(_1430_),
    .Y(_1446_));
 sky130_fd_sc_hd__mux2_1 _3190_ (.A0(\tms1x00.RAM[121][0] ),
    .A1(_1324_),
    .S(_1446_),
    .X(_1447_));
 sky130_fd_sc_hd__clkbuf_1 _3191_ (.A(_1447_),
    .X(_0187_));
 sky130_fd_sc_hd__mux2_1 _3192_ (.A0(\tms1x00.RAM[121][1] ),
    .A1(_1328_),
    .S(_1446_),
    .X(_1448_));
 sky130_fd_sc_hd__clkbuf_1 _3193_ (.A(_1448_),
    .X(_0188_));
 sky130_fd_sc_hd__mux2_1 _3194_ (.A0(\tms1x00.RAM[121][2] ),
    .A1(_1331_),
    .S(_1446_),
    .X(_1449_));
 sky130_fd_sc_hd__clkbuf_1 _3195_ (.A(_1449_),
    .X(_0189_));
 sky130_fd_sc_hd__mux2_1 _3196_ (.A0(\tms1x00.RAM[121][3] ),
    .A1(_1334_),
    .S(_1446_),
    .X(_1450_));
 sky130_fd_sc_hd__clkbuf_1 _3197_ (.A(_1450_),
    .X(_0190_));
 sky130_fd_sc_hd__nor2_2 _3198_ (.A(_1303_),
    .B(_1430_),
    .Y(_1451_));
 sky130_fd_sc_hd__mux2_1 _3199_ (.A0(\tms1x00.RAM[120][0] ),
    .A1(_1324_),
    .S(_1451_),
    .X(_1452_));
 sky130_fd_sc_hd__clkbuf_1 _3200_ (.A(_1452_),
    .X(_0191_));
 sky130_fd_sc_hd__mux2_1 _3201_ (.A0(\tms1x00.RAM[120][1] ),
    .A1(_1328_),
    .S(_1451_),
    .X(_1453_));
 sky130_fd_sc_hd__clkbuf_1 _3202_ (.A(_1453_),
    .X(_0192_));
 sky130_fd_sc_hd__mux2_1 _3203_ (.A0(\tms1x00.RAM[120][2] ),
    .A1(_1331_),
    .S(_1451_),
    .X(_1454_));
 sky130_fd_sc_hd__clkbuf_1 _3204_ (.A(_1454_),
    .X(_0193_));
 sky130_fd_sc_hd__mux2_1 _3205_ (.A0(\tms1x00.RAM[120][3] ),
    .A1(_1334_),
    .S(_1451_),
    .X(_1455_));
 sky130_fd_sc_hd__clkbuf_1 _3206_ (.A(_1455_),
    .X(_0194_));
 sky130_fd_sc_hd__clkbuf_4 _3207_ (.A(_1323_),
    .X(_1456_));
 sky130_fd_sc_hd__nor2_2 _3208_ (.A(_1286_),
    .B(_1344_),
    .Y(_1457_));
 sky130_fd_sc_hd__mux2_1 _3209_ (.A0(\tms1x00.RAM[11][0] ),
    .A1(_1456_),
    .S(_1457_),
    .X(_1458_));
 sky130_fd_sc_hd__clkbuf_1 _3210_ (.A(_1458_),
    .X(_0195_));
 sky130_fd_sc_hd__buf_2 _3211_ (.A(_1327_),
    .X(_1459_));
 sky130_fd_sc_hd__mux2_1 _3212_ (.A0(\tms1x00.RAM[11][1] ),
    .A1(_1459_),
    .S(_1457_),
    .X(_1460_));
 sky130_fd_sc_hd__clkbuf_1 _3213_ (.A(_1460_),
    .X(_0196_));
 sky130_fd_sc_hd__clkbuf_4 _3214_ (.A(_1330_),
    .X(_1461_));
 sky130_fd_sc_hd__mux2_1 _3215_ (.A0(\tms1x00.RAM[11][2] ),
    .A1(_1461_),
    .S(_1457_),
    .X(_1462_));
 sky130_fd_sc_hd__clkbuf_1 _3216_ (.A(_1462_),
    .X(_0197_));
 sky130_fd_sc_hd__buf_2 _3217_ (.A(_1333_),
    .X(_1463_));
 sky130_fd_sc_hd__mux2_1 _3218_ (.A0(\tms1x00.RAM[11][3] ),
    .A1(_1463_),
    .S(_1457_),
    .X(_1464_));
 sky130_fd_sc_hd__clkbuf_1 _3219_ (.A(_1464_),
    .X(_0198_));
 sky130_fd_sc_hd__nor2_2 _3220_ (.A(_1317_),
    .B(_1430_),
    .Y(_1465_));
 sky130_fd_sc_hd__mux2_1 _3221_ (.A0(\tms1x00.RAM[118][0] ),
    .A1(_1456_),
    .S(_1465_),
    .X(_1466_));
 sky130_fd_sc_hd__clkbuf_1 _3222_ (.A(_1466_),
    .X(_0199_));
 sky130_fd_sc_hd__mux2_1 _3223_ (.A0(\tms1x00.RAM[118][1] ),
    .A1(_1459_),
    .S(_1465_),
    .X(_1467_));
 sky130_fd_sc_hd__clkbuf_1 _3224_ (.A(_1467_),
    .X(_0200_));
 sky130_fd_sc_hd__mux2_1 _3225_ (.A0(\tms1x00.RAM[118][2] ),
    .A1(_1461_),
    .S(_1465_),
    .X(_1468_));
 sky130_fd_sc_hd__clkbuf_1 _3226_ (.A(_1468_),
    .X(_0201_));
 sky130_fd_sc_hd__mux2_1 _3227_ (.A0(\tms1x00.RAM[118][3] ),
    .A1(_1463_),
    .S(_1465_),
    .X(_1469_));
 sky130_fd_sc_hd__clkbuf_1 _3228_ (.A(_1469_),
    .X(_0202_));
 sky130_fd_sc_hd__nor2_2 _3229_ (.A(_1240_),
    .B(_1430_),
    .Y(_1470_));
 sky130_fd_sc_hd__mux2_1 _3230_ (.A0(\tms1x00.RAM[117][0] ),
    .A1(_1456_),
    .S(_1470_),
    .X(_1471_));
 sky130_fd_sc_hd__clkbuf_1 _3231_ (.A(_1471_),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_1 _3232_ (.A0(\tms1x00.RAM[117][1] ),
    .A1(_1459_),
    .S(_1470_),
    .X(_1472_));
 sky130_fd_sc_hd__clkbuf_1 _3233_ (.A(_1472_),
    .X(_0204_));
 sky130_fd_sc_hd__mux2_1 _3234_ (.A0(\tms1x00.RAM[117][2] ),
    .A1(_1461_),
    .S(_1470_),
    .X(_1473_));
 sky130_fd_sc_hd__clkbuf_1 _3235_ (.A(_1473_),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _3236_ (.A0(\tms1x00.RAM[117][3] ),
    .A1(_1463_),
    .S(_1470_),
    .X(_1474_));
 sky130_fd_sc_hd__clkbuf_1 _3237_ (.A(_1474_),
    .X(_0206_));
 sky130_fd_sc_hd__nor2_2 _3238_ (.A(_1337_),
    .B(_1430_),
    .Y(_1475_));
 sky130_fd_sc_hd__mux2_1 _3239_ (.A0(\tms1x00.RAM[116][0] ),
    .A1(_1456_),
    .S(_1475_),
    .X(_1476_));
 sky130_fd_sc_hd__clkbuf_1 _3240_ (.A(_1476_),
    .X(_0207_));
 sky130_fd_sc_hd__mux2_1 _3241_ (.A0(\tms1x00.RAM[116][1] ),
    .A1(_1459_),
    .S(_1475_),
    .X(_1477_));
 sky130_fd_sc_hd__clkbuf_1 _3242_ (.A(_1477_),
    .X(_0208_));
 sky130_fd_sc_hd__mux2_1 _3243_ (.A0(\tms1x00.RAM[116][2] ),
    .A1(_1461_),
    .S(_1475_),
    .X(_1478_));
 sky130_fd_sc_hd__clkbuf_1 _3244_ (.A(_1478_),
    .X(_0209_));
 sky130_fd_sc_hd__mux2_1 _3245_ (.A0(\tms1x00.RAM[116][3] ),
    .A1(_1463_),
    .S(_1475_),
    .X(_1479_));
 sky130_fd_sc_hd__clkbuf_1 _3246_ (.A(_1479_),
    .X(_0210_));
 sky130_fd_sc_hd__or2_2 _3247_ (.A(_1229_),
    .B(_1375_),
    .X(_1480_));
 sky130_fd_sc_hd__mux2_1 _3248_ (.A0(_1361_),
    .A1(\tms1x00.RAM[115][0] ),
    .S(_1480_),
    .X(_1481_));
 sky130_fd_sc_hd__clkbuf_1 _3249_ (.A(_1481_),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_1 _3250_ (.A0(_1364_),
    .A1(\tms1x00.RAM[115][1] ),
    .S(_1480_),
    .X(_1482_));
 sky130_fd_sc_hd__clkbuf_1 _3251_ (.A(_1482_),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_1 _3252_ (.A0(_1366_),
    .A1(\tms1x00.RAM[115][2] ),
    .S(_1480_),
    .X(_1483_));
 sky130_fd_sc_hd__clkbuf_1 _3253_ (.A(_1483_),
    .X(_0213_));
 sky130_fd_sc_hd__mux2_1 _3254_ (.A0(_1368_),
    .A1(\tms1x00.RAM[115][3] ),
    .S(_1480_),
    .X(_1484_));
 sky130_fd_sc_hd__clkbuf_1 _3255_ (.A(_1484_),
    .X(_0214_));
 sky130_fd_sc_hd__clkbuf_4 _3256_ (.A(_0911_),
    .X(_1485_));
 sky130_fd_sc_hd__or2_2 _3257_ (.A(_1430_),
    .B(_1396_),
    .X(_1486_));
 sky130_fd_sc_hd__mux2_1 _3258_ (.A0(_1485_),
    .A1(\tms1x00.RAM[126][0] ),
    .S(_1486_),
    .X(_1487_));
 sky130_fd_sc_hd__clkbuf_1 _3259_ (.A(_1487_),
    .X(_0215_));
 sky130_fd_sc_hd__buf_2 _3260_ (.A(_1034_),
    .X(_1488_));
 sky130_fd_sc_hd__mux2_1 _3261_ (.A0(_1488_),
    .A1(\tms1x00.RAM[126][1] ),
    .S(_1486_),
    .X(_1489_));
 sky130_fd_sc_hd__clkbuf_1 _3262_ (.A(_1489_),
    .X(_0216_));
 sky130_fd_sc_hd__buf_2 _3263_ (.A(_1129_),
    .X(_1490_));
 sky130_fd_sc_hd__mux2_1 _3264_ (.A0(_1490_),
    .A1(\tms1x00.RAM[126][2] ),
    .S(_1486_),
    .X(_1491_));
 sky130_fd_sc_hd__clkbuf_1 _3265_ (.A(_1491_),
    .X(_0217_));
 sky130_fd_sc_hd__buf_2 _3266_ (.A(_1224_),
    .X(_1492_));
 sky130_fd_sc_hd__mux2_1 _3267_ (.A0(_1492_),
    .A1(\tms1x00.RAM[126][3] ),
    .S(_1486_),
    .X(_1493_));
 sky130_fd_sc_hd__clkbuf_1 _3268_ (.A(_1493_),
    .X(_0218_));
 sky130_fd_sc_hd__or2_1 _3269_ (.A(_0917_),
    .B(_1375_),
    .X(_1494_));
 sky130_fd_sc_hd__mux2_1 _3270_ (.A0(_1485_),
    .A1(\tms1x00.RAM[125][0] ),
    .S(_1494_),
    .X(_1495_));
 sky130_fd_sc_hd__clkbuf_1 _3271_ (.A(_1495_),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _3272_ (.A0(_1488_),
    .A1(\tms1x00.RAM[125][1] ),
    .S(_1494_),
    .X(_1496_));
 sky130_fd_sc_hd__clkbuf_1 _3273_ (.A(_1496_),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _3274_ (.A0(_1490_),
    .A1(\tms1x00.RAM[125][2] ),
    .S(_1494_),
    .X(_1497_));
 sky130_fd_sc_hd__clkbuf_1 _3275_ (.A(_1497_),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _3276_ (.A0(_1492_),
    .A1(\tms1x00.RAM[125][3] ),
    .S(_1494_),
    .X(_1498_));
 sky130_fd_sc_hd__clkbuf_1 _3277_ (.A(_1498_),
    .X(_0222_));
 sky130_fd_sc_hd__nor2_2 _3278_ (.A(_1250_),
    .B(_1261_),
    .Y(_1499_));
 sky130_fd_sc_hd__mux2_1 _3279_ (.A0(\tms1x00.RAM[25][0] ),
    .A1(_1456_),
    .S(_1499_),
    .X(_1500_));
 sky130_fd_sc_hd__clkbuf_1 _3280_ (.A(_1500_),
    .X(_0223_));
 sky130_fd_sc_hd__mux2_1 _3281_ (.A0(\tms1x00.RAM[25][1] ),
    .A1(_1459_),
    .S(_1499_),
    .X(_1501_));
 sky130_fd_sc_hd__clkbuf_1 _3282_ (.A(_1501_),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_1 _3283_ (.A0(\tms1x00.RAM[25][2] ),
    .A1(_1461_),
    .S(_1499_),
    .X(_1502_));
 sky130_fd_sc_hd__clkbuf_1 _3284_ (.A(_1502_),
    .X(_0225_));
 sky130_fd_sc_hd__mux2_1 _3285_ (.A0(\tms1x00.RAM[25][3] ),
    .A1(_1463_),
    .S(_1499_),
    .X(_1503_));
 sky130_fd_sc_hd__clkbuf_1 _3286_ (.A(_1503_),
    .X(_0226_));
 sky130_fd_sc_hd__nor2_2 _3287_ (.A(_1250_),
    .B(_1303_),
    .Y(_1504_));
 sky130_fd_sc_hd__mux2_1 _3288_ (.A0(\tms1x00.RAM[24][0] ),
    .A1(_1456_),
    .S(_1504_),
    .X(_1505_));
 sky130_fd_sc_hd__clkbuf_1 _3289_ (.A(_1505_),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_1 _3290_ (.A0(\tms1x00.RAM[24][1] ),
    .A1(_1459_),
    .S(_1504_),
    .X(_1506_));
 sky130_fd_sc_hd__clkbuf_1 _3291_ (.A(_1506_),
    .X(_0228_));
 sky130_fd_sc_hd__mux2_1 _3292_ (.A0(\tms1x00.RAM[24][2] ),
    .A1(_1461_),
    .S(_1504_),
    .X(_1507_));
 sky130_fd_sc_hd__clkbuf_1 _3293_ (.A(_1507_),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_1 _3294_ (.A0(\tms1x00.RAM[24][3] ),
    .A1(_1463_),
    .S(_1504_),
    .X(_1508_));
 sky130_fd_sc_hd__clkbuf_1 _3295_ (.A(_1508_),
    .X(_0230_));
 sky130_fd_sc_hd__or2_2 _3296_ (.A(_1249_),
    .B(_1409_),
    .X(_1509_));
 sky130_fd_sc_hd__mux2_1 _3297_ (.A0(_1485_),
    .A1(\tms1x00.RAM[28][0] ),
    .S(_1509_),
    .X(_1510_));
 sky130_fd_sc_hd__clkbuf_1 _3298_ (.A(_1510_),
    .X(_0231_));
 sky130_fd_sc_hd__mux2_1 _3299_ (.A0(_1488_),
    .A1(\tms1x00.RAM[28][1] ),
    .S(_1509_),
    .X(_1511_));
 sky130_fd_sc_hd__clkbuf_1 _3300_ (.A(_1511_),
    .X(_0232_));
 sky130_fd_sc_hd__mux2_1 _3301_ (.A0(_1490_),
    .A1(\tms1x00.RAM[28][2] ),
    .S(_1509_),
    .X(_1512_));
 sky130_fd_sc_hd__clkbuf_1 _3302_ (.A(_1512_),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_1 _3303_ (.A0(_1492_),
    .A1(\tms1x00.RAM[28][3] ),
    .S(_1509_),
    .X(_1513_));
 sky130_fd_sc_hd__clkbuf_1 _3304_ (.A(_1513_),
    .X(_0234_));
 sky130_fd_sc_hd__nor2_2 _3305_ (.A(_1250_),
    .B(_1286_),
    .Y(_1514_));
 sky130_fd_sc_hd__mux2_1 _3306_ (.A0(\tms1x00.RAM[27][0] ),
    .A1(_1456_),
    .S(_1514_),
    .X(_1515_));
 sky130_fd_sc_hd__clkbuf_1 _3307_ (.A(_1515_),
    .X(_0235_));
 sky130_fd_sc_hd__mux2_1 _3308_ (.A0(\tms1x00.RAM[27][1] ),
    .A1(_1459_),
    .S(_1514_),
    .X(_1516_));
 sky130_fd_sc_hd__clkbuf_1 _3309_ (.A(_1516_),
    .X(_0236_));
 sky130_fd_sc_hd__mux2_1 _3310_ (.A0(\tms1x00.RAM[27][2] ),
    .A1(_1461_),
    .S(_1514_),
    .X(_1517_));
 sky130_fd_sc_hd__clkbuf_1 _3311_ (.A(_1517_),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _3312_ (.A0(\tms1x00.RAM[27][3] ),
    .A1(_1463_),
    .S(_1514_),
    .X(_1518_));
 sky130_fd_sc_hd__clkbuf_1 _3313_ (.A(_1518_),
    .X(_0238_));
 sky130_fd_sc_hd__nor2_2 _3314_ (.A(_1250_),
    .B(_1403_),
    .Y(_1519_));
 sky130_fd_sc_hd__mux2_1 _3315_ (.A0(\tms1x00.RAM[26][0] ),
    .A1(_1456_),
    .S(_1519_),
    .X(_1520_));
 sky130_fd_sc_hd__clkbuf_1 _3316_ (.A(_1520_),
    .X(_0239_));
 sky130_fd_sc_hd__mux2_1 _3317_ (.A0(\tms1x00.RAM[26][1] ),
    .A1(_1459_),
    .S(_1519_),
    .X(_1521_));
 sky130_fd_sc_hd__clkbuf_1 _3318_ (.A(_1521_),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _3319_ (.A0(\tms1x00.RAM[26][2] ),
    .A1(_1461_),
    .S(_1519_),
    .X(_1522_));
 sky130_fd_sc_hd__clkbuf_1 _3320_ (.A(_1522_),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_1 _3321_ (.A0(\tms1x00.RAM[26][3] ),
    .A1(_1463_),
    .S(_1519_),
    .X(_1523_));
 sky130_fd_sc_hd__clkbuf_1 _3322_ (.A(_1523_),
    .X(_0242_));
 sky130_fd_sc_hd__or3b_2 _3323_ (.A(\tms1x00.ram_addr_buff[4] ),
    .B(\tms1x00.ram_addr_buff[6] ),
    .C_N(\tms1x00.ram_addr_buff[5] ),
    .X(_1524_));
 sky130_fd_sc_hd__buf_4 _3324_ (.A(_1524_),
    .X(_1525_));
 sky130_fd_sc_hd__or2_2 _3325_ (.A(_1345_),
    .B(_1525_),
    .X(_1526_));
 sky130_fd_sc_hd__mux2_1 _3326_ (.A0(_1485_),
    .A1(\tms1x00.RAM[32][0] ),
    .S(_1526_),
    .X(_1527_));
 sky130_fd_sc_hd__clkbuf_1 _3327_ (.A(_1527_),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _3328_ (.A0(_1488_),
    .A1(\tms1x00.RAM[32][1] ),
    .S(_1526_),
    .X(_1528_));
 sky130_fd_sc_hd__clkbuf_1 _3329_ (.A(_1528_),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _3330_ (.A0(_1490_),
    .A1(\tms1x00.RAM[32][2] ),
    .S(_1526_),
    .X(_1529_));
 sky130_fd_sc_hd__clkbuf_1 _3331_ (.A(_1529_),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _3332_ (.A0(_1492_),
    .A1(\tms1x00.RAM[32][3] ),
    .S(_1526_),
    .X(_1530_));
 sky130_fd_sc_hd__clkbuf_1 _3333_ (.A(_1530_),
    .X(_0246_));
 sky130_fd_sc_hd__or2_2 _3334_ (.A(_1249_),
    .B(_1267_),
    .X(_1531_));
 sky130_fd_sc_hd__mux2_1 _3335_ (.A0(_1485_),
    .A1(\tms1x00.RAM[31][0] ),
    .S(_1531_),
    .X(_1532_));
 sky130_fd_sc_hd__clkbuf_1 _3336_ (.A(_1532_),
    .X(_0247_));
 sky130_fd_sc_hd__mux2_1 _3337_ (.A0(_1488_),
    .A1(\tms1x00.RAM[31][1] ),
    .S(_1531_),
    .X(_1533_));
 sky130_fd_sc_hd__clkbuf_1 _3338_ (.A(_1533_),
    .X(_0248_));
 sky130_fd_sc_hd__mux2_1 _3339_ (.A0(_1490_),
    .A1(\tms1x00.RAM[31][2] ),
    .S(_1531_),
    .X(_1534_));
 sky130_fd_sc_hd__clkbuf_1 _3340_ (.A(_1534_),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _3341_ (.A0(_1492_),
    .A1(\tms1x00.RAM[31][3] ),
    .S(_1531_),
    .X(_1535_));
 sky130_fd_sc_hd__clkbuf_1 _3342_ (.A(_1535_),
    .X(_0250_));
 sky130_fd_sc_hd__or2_2 _3343_ (.A(_1249_),
    .B(_1396_),
    .X(_1536_));
 sky130_fd_sc_hd__mux2_1 _3344_ (.A0(_1485_),
    .A1(\tms1x00.RAM[30][0] ),
    .S(_1536_),
    .X(_1537_));
 sky130_fd_sc_hd__clkbuf_1 _3345_ (.A(_1537_),
    .X(_0251_));
 sky130_fd_sc_hd__mux2_1 _3346_ (.A0(_1488_),
    .A1(\tms1x00.RAM[30][1] ),
    .S(_1536_),
    .X(_1538_));
 sky130_fd_sc_hd__clkbuf_1 _3347_ (.A(_1538_),
    .X(_0252_));
 sky130_fd_sc_hd__mux2_1 _3348_ (.A0(_1490_),
    .A1(\tms1x00.RAM[30][2] ),
    .S(_1536_),
    .X(_1539_));
 sky130_fd_sc_hd__clkbuf_1 _3349_ (.A(_1539_),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _3350_ (.A0(_1492_),
    .A1(\tms1x00.RAM[30][3] ),
    .S(_1536_),
    .X(_1540_));
 sky130_fd_sc_hd__clkbuf_1 _3351_ (.A(_1540_),
    .X(_0254_));
 sky130_fd_sc_hd__or2_2 _3352_ (.A(_1273_),
    .B(_1343_),
    .X(_1541_));
 sky130_fd_sc_hd__mux2_1 _3353_ (.A0(_1485_),
    .A1(\tms1x00.RAM[2][0] ),
    .S(_1541_),
    .X(_1542_));
 sky130_fd_sc_hd__clkbuf_1 _3354_ (.A(_1542_),
    .X(_0255_));
 sky130_fd_sc_hd__mux2_1 _3355_ (.A0(_1488_),
    .A1(\tms1x00.RAM[2][1] ),
    .S(_1541_),
    .X(_1543_));
 sky130_fd_sc_hd__clkbuf_1 _3356_ (.A(_1543_),
    .X(_0256_));
 sky130_fd_sc_hd__mux2_1 _3357_ (.A0(_1490_),
    .A1(\tms1x00.RAM[2][2] ),
    .S(_1541_),
    .X(_1544_));
 sky130_fd_sc_hd__clkbuf_1 _3358_ (.A(_1544_),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _3359_ (.A0(_1492_),
    .A1(\tms1x00.RAM[2][3] ),
    .S(_1541_),
    .X(_1545_));
 sky130_fd_sc_hd__clkbuf_1 _3360_ (.A(_1545_),
    .X(_0258_));
 sky130_fd_sc_hd__nor2_2 _3361_ (.A(_1240_),
    .B(_1525_),
    .Y(_1546_));
 sky130_fd_sc_hd__mux2_1 _3362_ (.A0(\tms1x00.RAM[37][0] ),
    .A1(_1456_),
    .S(_1546_),
    .X(_1547_));
 sky130_fd_sc_hd__clkbuf_1 _3363_ (.A(_1547_),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _3364_ (.A0(\tms1x00.RAM[37][1] ),
    .A1(_1459_),
    .S(_1546_),
    .X(_1548_));
 sky130_fd_sc_hd__clkbuf_1 _3365_ (.A(_1548_),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_1 _3366_ (.A0(\tms1x00.RAM[37][2] ),
    .A1(_1461_),
    .S(_1546_),
    .X(_1549_));
 sky130_fd_sc_hd__clkbuf_1 _3367_ (.A(_1549_),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _3368_ (.A0(\tms1x00.RAM[37][3] ),
    .A1(_1463_),
    .S(_1546_),
    .X(_1550_));
 sky130_fd_sc_hd__clkbuf_1 _3369_ (.A(_1550_),
    .X(_0262_));
 sky130_fd_sc_hd__nor2_2 _3370_ (.A(_1337_),
    .B(_1525_),
    .Y(_1551_));
 sky130_fd_sc_hd__mux2_1 _3371_ (.A0(\tms1x00.RAM[36][0] ),
    .A1(_1456_),
    .S(_1551_),
    .X(_1552_));
 sky130_fd_sc_hd__clkbuf_1 _3372_ (.A(_1552_),
    .X(_0263_));
 sky130_fd_sc_hd__mux2_1 _3373_ (.A0(\tms1x00.RAM[36][1] ),
    .A1(_1459_),
    .S(_1551_),
    .X(_1553_));
 sky130_fd_sc_hd__clkbuf_1 _3374_ (.A(_1553_),
    .X(_0264_));
 sky130_fd_sc_hd__mux2_1 _3375_ (.A0(\tms1x00.RAM[36][2] ),
    .A1(_1461_),
    .S(_1551_),
    .X(_1554_));
 sky130_fd_sc_hd__clkbuf_1 _3376_ (.A(_1554_),
    .X(_0265_));
 sky130_fd_sc_hd__mux2_1 _3377_ (.A0(\tms1x00.RAM[36][3] ),
    .A1(_1463_),
    .S(_1551_),
    .X(_1555_));
 sky130_fd_sc_hd__clkbuf_1 _3378_ (.A(_1555_),
    .X(_0266_));
 sky130_fd_sc_hd__or2_2 _3379_ (.A(_1229_),
    .B(_1525_),
    .X(_1556_));
 sky130_fd_sc_hd__mux2_1 _3380_ (.A0(_1485_),
    .A1(\tms1x00.RAM[35][0] ),
    .S(_1556_),
    .X(_1557_));
 sky130_fd_sc_hd__clkbuf_1 _3381_ (.A(_1557_),
    .X(_0267_));
 sky130_fd_sc_hd__mux2_1 _3382_ (.A0(_1488_),
    .A1(\tms1x00.RAM[35][1] ),
    .S(_1556_),
    .X(_1558_));
 sky130_fd_sc_hd__clkbuf_1 _3383_ (.A(_1558_),
    .X(_0268_));
 sky130_fd_sc_hd__mux2_1 _3384_ (.A0(_1490_),
    .A1(\tms1x00.RAM[35][2] ),
    .S(_1556_),
    .X(_1559_));
 sky130_fd_sc_hd__clkbuf_1 _3385_ (.A(_1559_),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _3386_ (.A0(_1492_),
    .A1(\tms1x00.RAM[35][3] ),
    .S(_1556_),
    .X(_1560_));
 sky130_fd_sc_hd__clkbuf_1 _3387_ (.A(_1560_),
    .X(_0270_));
 sky130_fd_sc_hd__or2_2 _3388_ (.A(_1273_),
    .B(_1524_),
    .X(_1561_));
 sky130_fd_sc_hd__mux2_1 _3389_ (.A0(_1485_),
    .A1(\tms1x00.RAM[34][0] ),
    .S(_1561_),
    .X(_1562_));
 sky130_fd_sc_hd__clkbuf_1 _3390_ (.A(_1562_),
    .X(_0271_));
 sky130_fd_sc_hd__mux2_1 _3391_ (.A0(_1488_),
    .A1(\tms1x00.RAM[34][1] ),
    .S(_1561_),
    .X(_1563_));
 sky130_fd_sc_hd__clkbuf_1 _3392_ (.A(_1563_),
    .X(_0272_));
 sky130_fd_sc_hd__mux2_1 _3393_ (.A0(_1490_),
    .A1(\tms1x00.RAM[34][2] ),
    .S(_1561_),
    .X(_1564_));
 sky130_fd_sc_hd__clkbuf_1 _3394_ (.A(_1564_),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _3395_ (.A0(_1492_),
    .A1(\tms1x00.RAM[34][3] ),
    .S(_1561_),
    .X(_1565_));
 sky130_fd_sc_hd__clkbuf_1 _3396_ (.A(_1565_),
    .X(_0274_));
 sky130_fd_sc_hd__or2_2 _3397_ (.A(_1251_),
    .B(_1524_),
    .X(_1566_));
 sky130_fd_sc_hd__mux2_1 _3398_ (.A0(_1485_),
    .A1(\tms1x00.RAM[33][0] ),
    .S(_1566_),
    .X(_1567_));
 sky130_fd_sc_hd__clkbuf_1 _3399_ (.A(_1567_),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_1 _3400_ (.A0(_1488_),
    .A1(\tms1x00.RAM[33][1] ),
    .S(_1566_),
    .X(_1568_));
 sky130_fd_sc_hd__clkbuf_1 _3401_ (.A(_1568_),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_1 _3402_ (.A0(_1490_),
    .A1(\tms1x00.RAM[33][2] ),
    .S(_1566_),
    .X(_1569_));
 sky130_fd_sc_hd__clkbuf_1 _3403_ (.A(_1569_),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_1 _3404_ (.A0(_1492_),
    .A1(\tms1x00.RAM[33][3] ),
    .S(_1566_),
    .X(_1570_));
 sky130_fd_sc_hd__clkbuf_1 _3405_ (.A(_1570_),
    .X(_0278_));
 sky130_fd_sc_hd__clkbuf_4 _3406_ (.A(_0911_),
    .X(_1571_));
 sky130_fd_sc_hd__nor2_2 _3407_ (.A(_1261_),
    .B(_1525_),
    .Y(_1572_));
 sky130_fd_sc_hd__mux2_1 _3408_ (.A0(\tms1x00.RAM[41][0] ),
    .A1(_1571_),
    .S(_1572_),
    .X(_1573_));
 sky130_fd_sc_hd__clkbuf_1 _3409_ (.A(_1573_),
    .X(_0279_));
 sky130_fd_sc_hd__clkbuf_4 _3410_ (.A(_1034_),
    .X(_1574_));
 sky130_fd_sc_hd__mux2_1 _3411_ (.A0(\tms1x00.RAM[41][1] ),
    .A1(_1574_),
    .S(_1572_),
    .X(_1575_));
 sky130_fd_sc_hd__clkbuf_1 _3412_ (.A(_1575_),
    .X(_0280_));
 sky130_fd_sc_hd__clkbuf_4 _3413_ (.A(_1129_),
    .X(_1576_));
 sky130_fd_sc_hd__mux2_1 _3414_ (.A0(\tms1x00.RAM[41][2] ),
    .A1(_1576_),
    .S(_1572_),
    .X(_1577_));
 sky130_fd_sc_hd__clkbuf_1 _3415_ (.A(_1577_),
    .X(_0281_));
 sky130_fd_sc_hd__clkbuf_4 _3416_ (.A(_1224_),
    .X(_1578_));
 sky130_fd_sc_hd__mux2_1 _3417_ (.A0(\tms1x00.RAM[41][3] ),
    .A1(_1578_),
    .S(_1572_),
    .X(_1579_));
 sky130_fd_sc_hd__clkbuf_1 _3418_ (.A(_1579_),
    .X(_0282_));
 sky130_fd_sc_hd__nor2_2 _3419_ (.A(_1303_),
    .B(_1525_),
    .Y(_1580_));
 sky130_fd_sc_hd__mux2_1 _3420_ (.A0(\tms1x00.RAM[40][0] ),
    .A1(_1571_),
    .S(_1580_),
    .X(_1581_));
 sky130_fd_sc_hd__clkbuf_1 _3421_ (.A(_1581_),
    .X(_0283_));
 sky130_fd_sc_hd__mux2_1 _3422_ (.A0(\tms1x00.RAM[40][1] ),
    .A1(_1574_),
    .S(_1580_),
    .X(_1582_));
 sky130_fd_sc_hd__clkbuf_1 _3423_ (.A(_1582_),
    .X(_0284_));
 sky130_fd_sc_hd__mux2_1 _3424_ (.A0(\tms1x00.RAM[40][2] ),
    .A1(_1576_),
    .S(_1580_),
    .X(_1583_));
 sky130_fd_sc_hd__clkbuf_1 _3425_ (.A(_1583_),
    .X(_0285_));
 sky130_fd_sc_hd__mux2_1 _3426_ (.A0(\tms1x00.RAM[40][3] ),
    .A1(_1578_),
    .S(_1580_),
    .X(_1584_));
 sky130_fd_sc_hd__clkbuf_1 _3427_ (.A(_1584_),
    .X(_0286_));
 sky130_fd_sc_hd__buf_2 _3428_ (.A(_0911_),
    .X(_1585_));
 sky130_fd_sc_hd__or2_2 _3429_ (.A(_1229_),
    .B(_1343_),
    .X(_1586_));
 sky130_fd_sc_hd__mux2_1 _3430_ (.A0(_1585_),
    .A1(\tms1x00.RAM[3][0] ),
    .S(_1586_),
    .X(_1587_));
 sky130_fd_sc_hd__clkbuf_1 _3431_ (.A(_1587_),
    .X(_0287_));
 sky130_fd_sc_hd__buf_2 _3432_ (.A(_1034_),
    .X(_1588_));
 sky130_fd_sc_hd__mux2_1 _3433_ (.A0(_1588_),
    .A1(\tms1x00.RAM[3][1] ),
    .S(_1586_),
    .X(_1589_));
 sky130_fd_sc_hd__clkbuf_1 _3434_ (.A(_1589_),
    .X(_0288_));
 sky130_fd_sc_hd__buf_2 _3435_ (.A(_1129_),
    .X(_1590_));
 sky130_fd_sc_hd__mux2_1 _3436_ (.A0(_1590_),
    .A1(\tms1x00.RAM[3][2] ),
    .S(_1586_),
    .X(_1591_));
 sky130_fd_sc_hd__clkbuf_1 _3437_ (.A(_1591_),
    .X(_0289_));
 sky130_fd_sc_hd__buf_2 _3438_ (.A(_1224_),
    .X(_1592_));
 sky130_fd_sc_hd__mux2_1 _3439_ (.A0(_1592_),
    .A1(\tms1x00.RAM[3][3] ),
    .S(_1586_),
    .X(_1593_));
 sky130_fd_sc_hd__clkbuf_1 _3440_ (.A(_1593_),
    .X(_0290_));
 sky130_fd_sc_hd__nor2_2 _3441_ (.A(_1317_),
    .B(_1525_),
    .Y(_1594_));
 sky130_fd_sc_hd__mux2_1 _3442_ (.A0(\tms1x00.RAM[38][0] ),
    .A1(_1571_),
    .S(_1594_),
    .X(_1595_));
 sky130_fd_sc_hd__clkbuf_1 _3443_ (.A(_1595_),
    .X(_0291_));
 sky130_fd_sc_hd__mux2_1 _3444_ (.A0(\tms1x00.RAM[38][1] ),
    .A1(_1574_),
    .S(_1594_),
    .X(_1596_));
 sky130_fd_sc_hd__clkbuf_1 _3445_ (.A(_1596_),
    .X(_0292_));
 sky130_fd_sc_hd__mux2_1 _3446_ (.A0(\tms1x00.RAM[38][2] ),
    .A1(_1576_),
    .S(_1594_),
    .X(_1597_));
 sky130_fd_sc_hd__clkbuf_1 _3447_ (.A(_1597_),
    .X(_0293_));
 sky130_fd_sc_hd__mux2_1 _3448_ (.A0(\tms1x00.RAM[38][3] ),
    .A1(_1578_),
    .S(_1594_),
    .X(_1598_));
 sky130_fd_sc_hd__clkbuf_1 _3449_ (.A(_1598_),
    .X(_0294_));
 sky130_fd_sc_hd__or2_2 _3450_ (.A(_0917_),
    .B(_1524_),
    .X(_1599_));
 sky130_fd_sc_hd__mux2_1 _3451_ (.A0(_1585_),
    .A1(\tms1x00.RAM[45][0] ),
    .S(_1599_),
    .X(_1600_));
 sky130_fd_sc_hd__clkbuf_1 _3452_ (.A(_1600_),
    .X(_0295_));
 sky130_fd_sc_hd__mux2_1 _3453_ (.A0(_1588_),
    .A1(\tms1x00.RAM[45][1] ),
    .S(_1599_),
    .X(_1601_));
 sky130_fd_sc_hd__clkbuf_1 _3454_ (.A(_1601_),
    .X(_0296_));
 sky130_fd_sc_hd__mux2_1 _3455_ (.A0(_1590_),
    .A1(\tms1x00.RAM[45][2] ),
    .S(_1599_),
    .X(_1602_));
 sky130_fd_sc_hd__clkbuf_1 _3456_ (.A(_1602_),
    .X(_0297_));
 sky130_fd_sc_hd__mux2_1 _3457_ (.A0(_1592_),
    .A1(\tms1x00.RAM[45][3] ),
    .S(_1599_),
    .X(_1603_));
 sky130_fd_sc_hd__clkbuf_1 _3458_ (.A(_1603_),
    .X(_0298_));
 sky130_fd_sc_hd__or2_2 _3459_ (.A(_1409_),
    .B(_1524_),
    .X(_1604_));
 sky130_fd_sc_hd__mux2_1 _3460_ (.A0(_1585_),
    .A1(\tms1x00.RAM[44][0] ),
    .S(_1604_),
    .X(_1605_));
 sky130_fd_sc_hd__clkbuf_1 _3461_ (.A(_1605_),
    .X(_0299_));
 sky130_fd_sc_hd__mux2_1 _3462_ (.A0(_1588_),
    .A1(\tms1x00.RAM[44][1] ),
    .S(_1604_),
    .X(_1606_));
 sky130_fd_sc_hd__clkbuf_1 _3463_ (.A(_1606_),
    .X(_0300_));
 sky130_fd_sc_hd__mux2_1 _3464_ (.A0(_1590_),
    .A1(\tms1x00.RAM[44][2] ),
    .S(_1604_),
    .X(_1607_));
 sky130_fd_sc_hd__clkbuf_1 _3465_ (.A(_1607_),
    .X(_0301_));
 sky130_fd_sc_hd__mux2_1 _3466_ (.A0(_1592_),
    .A1(\tms1x00.RAM[44][3] ),
    .S(_1604_),
    .X(_1608_));
 sky130_fd_sc_hd__clkbuf_1 _3467_ (.A(_1608_),
    .X(_0302_));
 sky130_fd_sc_hd__nor2_2 _3468_ (.A(_1286_),
    .B(_1525_),
    .Y(_1609_));
 sky130_fd_sc_hd__mux2_1 _3469_ (.A0(\tms1x00.RAM[43][0] ),
    .A1(_1571_),
    .S(_1609_),
    .X(_1610_));
 sky130_fd_sc_hd__clkbuf_1 _3470_ (.A(_1610_),
    .X(_0303_));
 sky130_fd_sc_hd__mux2_1 _3471_ (.A0(\tms1x00.RAM[43][1] ),
    .A1(_1574_),
    .S(_1609_),
    .X(_1611_));
 sky130_fd_sc_hd__clkbuf_1 _3472_ (.A(_1611_),
    .X(_0304_));
 sky130_fd_sc_hd__mux2_1 _3473_ (.A0(\tms1x00.RAM[43][2] ),
    .A1(_1576_),
    .S(_1609_),
    .X(_1612_));
 sky130_fd_sc_hd__clkbuf_1 _3474_ (.A(_1612_),
    .X(_0305_));
 sky130_fd_sc_hd__mux2_1 _3475_ (.A0(\tms1x00.RAM[43][3] ),
    .A1(_1578_),
    .S(_1609_),
    .X(_1613_));
 sky130_fd_sc_hd__clkbuf_1 _3476_ (.A(_1613_),
    .X(_0306_));
 sky130_fd_sc_hd__nor2_2 _3477_ (.A(_1403_),
    .B(_1525_),
    .Y(_1614_));
 sky130_fd_sc_hd__mux2_1 _3478_ (.A0(\tms1x00.RAM[42][0] ),
    .A1(_1571_),
    .S(_1614_),
    .X(_1615_));
 sky130_fd_sc_hd__clkbuf_1 _3479_ (.A(_1615_),
    .X(_0307_));
 sky130_fd_sc_hd__mux2_1 _3480_ (.A0(\tms1x00.RAM[42][1] ),
    .A1(_1574_),
    .S(_1614_),
    .X(_1616_));
 sky130_fd_sc_hd__clkbuf_1 _3481_ (.A(_1616_),
    .X(_0308_));
 sky130_fd_sc_hd__mux2_1 _3482_ (.A0(\tms1x00.RAM[42][2] ),
    .A1(_1576_),
    .S(_1614_),
    .X(_1617_));
 sky130_fd_sc_hd__clkbuf_1 _3483_ (.A(_1617_),
    .X(_0309_));
 sky130_fd_sc_hd__mux2_1 _3484_ (.A0(\tms1x00.RAM[42][3] ),
    .A1(_1578_),
    .S(_1614_),
    .X(_1618_));
 sky130_fd_sc_hd__clkbuf_1 _3485_ (.A(_1618_),
    .X(_0310_));
 sky130_fd_sc_hd__or2_2 _3486_ (.A(_1273_),
    .B(_1283_),
    .X(_1619_));
 sky130_fd_sc_hd__mux2_1 _3487_ (.A0(_1585_),
    .A1(\tms1x00.RAM[50][0] ),
    .S(_1619_),
    .X(_1620_));
 sky130_fd_sc_hd__clkbuf_1 _3488_ (.A(_1620_),
    .X(_0311_));
 sky130_fd_sc_hd__mux2_1 _3489_ (.A0(_1588_),
    .A1(\tms1x00.RAM[50][1] ),
    .S(_1619_),
    .X(_1621_));
 sky130_fd_sc_hd__clkbuf_1 _3490_ (.A(_1621_),
    .X(_0312_));
 sky130_fd_sc_hd__mux2_1 _3491_ (.A0(_1590_),
    .A1(\tms1x00.RAM[50][2] ),
    .S(_1619_),
    .X(_1622_));
 sky130_fd_sc_hd__clkbuf_1 _3492_ (.A(_1622_),
    .X(_0313_));
 sky130_fd_sc_hd__mux2_1 _3493_ (.A0(_1592_),
    .A1(\tms1x00.RAM[50][3] ),
    .S(_1619_),
    .X(_1623_));
 sky130_fd_sc_hd__clkbuf_1 _3494_ (.A(_1623_),
    .X(_0314_));
 sky130_fd_sc_hd__nor2_2 _3495_ (.A(_1337_),
    .B(_1344_),
    .Y(_1624_));
 sky130_fd_sc_hd__mux2_1 _3496_ (.A0(\tms1x00.RAM[4][0] ),
    .A1(_1571_),
    .S(_1624_),
    .X(_1625_));
 sky130_fd_sc_hd__clkbuf_1 _3497_ (.A(_1625_),
    .X(_0315_));
 sky130_fd_sc_hd__mux2_1 _3498_ (.A0(\tms1x00.RAM[4][1] ),
    .A1(_1574_),
    .S(_1624_),
    .X(_1626_));
 sky130_fd_sc_hd__clkbuf_1 _3499_ (.A(_1626_),
    .X(_0316_));
 sky130_fd_sc_hd__mux2_1 _3500_ (.A0(\tms1x00.RAM[4][2] ),
    .A1(_1576_),
    .S(_1624_),
    .X(_1627_));
 sky130_fd_sc_hd__clkbuf_1 _3501_ (.A(_1627_),
    .X(_0317_));
 sky130_fd_sc_hd__mux2_1 _3502_ (.A0(\tms1x00.RAM[4][3] ),
    .A1(_1578_),
    .S(_1624_),
    .X(_1628_));
 sky130_fd_sc_hd__clkbuf_1 _3503_ (.A(_1628_),
    .X(_0318_));
 sky130_fd_sc_hd__or2_2 _3504_ (.A(_1284_),
    .B(_1345_),
    .X(_1629_));
 sky130_fd_sc_hd__mux2_1 _3505_ (.A0(_1585_),
    .A1(\tms1x00.RAM[48][0] ),
    .S(_1629_),
    .X(_1630_));
 sky130_fd_sc_hd__clkbuf_1 _3506_ (.A(_1630_),
    .X(_0319_));
 sky130_fd_sc_hd__mux2_1 _3507_ (.A0(_1588_),
    .A1(\tms1x00.RAM[48][1] ),
    .S(_1629_),
    .X(_1631_));
 sky130_fd_sc_hd__clkbuf_1 _3508_ (.A(_1631_),
    .X(_0320_));
 sky130_fd_sc_hd__mux2_1 _3509_ (.A0(_1590_),
    .A1(\tms1x00.RAM[48][2] ),
    .S(_1629_),
    .X(_1632_));
 sky130_fd_sc_hd__clkbuf_1 _3510_ (.A(_1632_),
    .X(_0321_));
 sky130_fd_sc_hd__mux2_1 _3511_ (.A0(_1592_),
    .A1(\tms1x00.RAM[48][3] ),
    .S(_1629_),
    .X(_1633_));
 sky130_fd_sc_hd__clkbuf_1 _3512_ (.A(_1633_),
    .X(_0322_));
 sky130_fd_sc_hd__or2_2 _3513_ (.A(_1267_),
    .B(_1524_),
    .X(_1634_));
 sky130_fd_sc_hd__mux2_1 _3514_ (.A0(_1585_),
    .A1(\tms1x00.RAM[47][0] ),
    .S(_1634_),
    .X(_1635_));
 sky130_fd_sc_hd__clkbuf_1 _3515_ (.A(_1635_),
    .X(_0323_));
 sky130_fd_sc_hd__mux2_1 _3516_ (.A0(_1588_),
    .A1(\tms1x00.RAM[47][1] ),
    .S(_1634_),
    .X(_1636_));
 sky130_fd_sc_hd__clkbuf_1 _3517_ (.A(_1636_),
    .X(_0324_));
 sky130_fd_sc_hd__mux2_1 _3518_ (.A0(_1590_),
    .A1(\tms1x00.RAM[47][2] ),
    .S(_1634_),
    .X(_1637_));
 sky130_fd_sc_hd__clkbuf_1 _3519_ (.A(_1637_),
    .X(_0325_));
 sky130_fd_sc_hd__mux2_1 _3520_ (.A0(_1592_),
    .A1(\tms1x00.RAM[47][3] ),
    .S(_1634_),
    .X(_1638_));
 sky130_fd_sc_hd__clkbuf_1 _3521_ (.A(_1638_),
    .X(_0326_));
 sky130_fd_sc_hd__or2_2 _3522_ (.A(_1396_),
    .B(_1524_),
    .X(_1639_));
 sky130_fd_sc_hd__mux2_1 _3523_ (.A0(_1585_),
    .A1(\tms1x00.RAM[46][0] ),
    .S(_1639_),
    .X(_1640_));
 sky130_fd_sc_hd__clkbuf_1 _3524_ (.A(_1640_),
    .X(_0327_));
 sky130_fd_sc_hd__mux2_1 _3525_ (.A0(_1588_),
    .A1(\tms1x00.RAM[46][1] ),
    .S(_1639_),
    .X(_1641_));
 sky130_fd_sc_hd__clkbuf_1 _3526_ (.A(_1641_),
    .X(_0328_));
 sky130_fd_sc_hd__mux2_1 _3527_ (.A0(_1590_),
    .A1(\tms1x00.RAM[46][2] ),
    .S(_1639_),
    .X(_1642_));
 sky130_fd_sc_hd__clkbuf_1 _3528_ (.A(_1642_),
    .X(_0329_));
 sky130_fd_sc_hd__mux2_1 _3529_ (.A0(_1592_),
    .A1(\tms1x00.RAM[46][3] ),
    .S(_1639_),
    .X(_1643_));
 sky130_fd_sc_hd__clkbuf_1 _3530_ (.A(_1643_),
    .X(_0330_));
 sky130_fd_sc_hd__nor2_2 _3531_ (.A(_1284_),
    .B(_1317_),
    .Y(_1644_));
 sky130_fd_sc_hd__mux2_1 _3532_ (.A0(\tms1x00.RAM[54][0] ),
    .A1(_1571_),
    .S(_1644_),
    .X(_1645_));
 sky130_fd_sc_hd__clkbuf_1 _3533_ (.A(_1645_),
    .X(_0331_));
 sky130_fd_sc_hd__mux2_1 _3534_ (.A0(\tms1x00.RAM[54][1] ),
    .A1(_1574_),
    .S(_1644_),
    .X(_1646_));
 sky130_fd_sc_hd__clkbuf_1 _3535_ (.A(_1646_),
    .X(_0332_));
 sky130_fd_sc_hd__mux2_1 _3536_ (.A0(\tms1x00.RAM[54][2] ),
    .A1(_1576_),
    .S(_1644_),
    .X(_1647_));
 sky130_fd_sc_hd__clkbuf_1 _3537_ (.A(_1647_),
    .X(_0333_));
 sky130_fd_sc_hd__mux2_1 _3538_ (.A0(\tms1x00.RAM[54][3] ),
    .A1(_1578_),
    .S(_1644_),
    .X(_1648_));
 sky130_fd_sc_hd__clkbuf_1 _3539_ (.A(_1648_),
    .X(_0334_));
 sky130_fd_sc_hd__nor2_2 _3540_ (.A(_1240_),
    .B(_1284_),
    .Y(_1649_));
 sky130_fd_sc_hd__mux2_1 _3541_ (.A0(\tms1x00.RAM[53][0] ),
    .A1(_1571_),
    .S(_1649_),
    .X(_1650_));
 sky130_fd_sc_hd__clkbuf_1 _3542_ (.A(_1650_),
    .X(_0335_));
 sky130_fd_sc_hd__mux2_1 _3543_ (.A0(\tms1x00.RAM[53][1] ),
    .A1(_1574_),
    .S(_1649_),
    .X(_1651_));
 sky130_fd_sc_hd__clkbuf_1 _3544_ (.A(_1651_),
    .X(_0336_));
 sky130_fd_sc_hd__mux2_1 _3545_ (.A0(\tms1x00.RAM[53][2] ),
    .A1(_1576_),
    .S(_1649_),
    .X(_1652_));
 sky130_fd_sc_hd__clkbuf_1 _3546_ (.A(_1652_),
    .X(_0337_));
 sky130_fd_sc_hd__mux2_1 _3547_ (.A0(\tms1x00.RAM[53][3] ),
    .A1(_1578_),
    .S(_1649_),
    .X(_1653_));
 sky130_fd_sc_hd__clkbuf_1 _3548_ (.A(_1653_),
    .X(_0338_));
 sky130_fd_sc_hd__nor2_2 _3549_ (.A(_1284_),
    .B(_1337_),
    .Y(_1654_));
 sky130_fd_sc_hd__mux2_1 _3550_ (.A0(\tms1x00.RAM[52][0] ),
    .A1(_1571_),
    .S(_1654_),
    .X(_1655_));
 sky130_fd_sc_hd__clkbuf_1 _3551_ (.A(_1655_),
    .X(_0339_));
 sky130_fd_sc_hd__mux2_1 _3552_ (.A0(\tms1x00.RAM[52][1] ),
    .A1(_1574_),
    .S(_1654_),
    .X(_1656_));
 sky130_fd_sc_hd__clkbuf_1 _3553_ (.A(_1656_),
    .X(_0340_));
 sky130_fd_sc_hd__mux2_1 _3554_ (.A0(\tms1x00.RAM[52][2] ),
    .A1(_1576_),
    .S(_1654_),
    .X(_1657_));
 sky130_fd_sc_hd__clkbuf_1 _3555_ (.A(_1657_),
    .X(_0341_));
 sky130_fd_sc_hd__mux2_1 _3556_ (.A0(\tms1x00.RAM[52][3] ),
    .A1(_1578_),
    .S(_1654_),
    .X(_1658_));
 sky130_fd_sc_hd__clkbuf_1 _3557_ (.A(_1658_),
    .X(_0342_));
 sky130_fd_sc_hd__or2_2 _3558_ (.A(_1229_),
    .B(_1283_),
    .X(_1659_));
 sky130_fd_sc_hd__mux2_1 _3559_ (.A0(_1585_),
    .A1(\tms1x00.RAM[51][0] ),
    .S(_1659_),
    .X(_1660_));
 sky130_fd_sc_hd__clkbuf_1 _3560_ (.A(_1660_),
    .X(_0343_));
 sky130_fd_sc_hd__mux2_1 _3561_ (.A0(_1588_),
    .A1(\tms1x00.RAM[51][1] ),
    .S(_1659_),
    .X(_1661_));
 sky130_fd_sc_hd__clkbuf_1 _3562_ (.A(_1661_),
    .X(_0344_));
 sky130_fd_sc_hd__mux2_1 _3563_ (.A0(_1590_),
    .A1(\tms1x00.RAM[51][2] ),
    .S(_1659_),
    .X(_1662_));
 sky130_fd_sc_hd__clkbuf_1 _3564_ (.A(_1662_),
    .X(_0345_));
 sky130_fd_sc_hd__mux2_1 _3565_ (.A0(_1592_),
    .A1(\tms1x00.RAM[51][3] ),
    .S(_1659_),
    .X(_1663_));
 sky130_fd_sc_hd__clkbuf_1 _3566_ (.A(_1663_),
    .X(_0346_));
 sky130_fd_sc_hd__nor2_2 _3567_ (.A(_1240_),
    .B(_1344_),
    .Y(_1664_));
 sky130_fd_sc_hd__mux2_1 _3568_ (.A0(\tms1x00.RAM[5][0] ),
    .A1(_1571_),
    .S(_1664_),
    .X(_1665_));
 sky130_fd_sc_hd__clkbuf_1 _3569_ (.A(_1665_),
    .X(_0347_));
 sky130_fd_sc_hd__mux2_1 _3570_ (.A0(\tms1x00.RAM[5][1] ),
    .A1(_1574_),
    .S(_1664_),
    .X(_1666_));
 sky130_fd_sc_hd__clkbuf_1 _3571_ (.A(_1666_),
    .X(_0348_));
 sky130_fd_sc_hd__mux2_1 _3572_ (.A0(\tms1x00.RAM[5][2] ),
    .A1(_1576_),
    .S(_1664_),
    .X(_1667_));
 sky130_fd_sc_hd__clkbuf_1 _3573_ (.A(_1667_),
    .X(_0349_));
 sky130_fd_sc_hd__mux2_1 _3574_ (.A0(\tms1x00.RAM[5][3] ),
    .A1(_1578_),
    .S(_1664_),
    .X(_1668_));
 sky130_fd_sc_hd__clkbuf_1 _3575_ (.A(_1668_),
    .X(_0350_));
 sky130_fd_sc_hd__clkbuf_4 _3576_ (.A(_0911_),
    .X(_1669_));
 sky130_fd_sc_hd__nor2_2 _3577_ (.A(_1284_),
    .B(_1403_),
    .Y(_1670_));
 sky130_fd_sc_hd__mux2_1 _3578_ (.A0(\tms1x00.RAM[58][0] ),
    .A1(_1669_),
    .S(_1670_),
    .X(_1671_));
 sky130_fd_sc_hd__clkbuf_1 _3579_ (.A(_1671_),
    .X(_0351_));
 sky130_fd_sc_hd__clkbuf_4 _3580_ (.A(_1034_),
    .X(_1672_));
 sky130_fd_sc_hd__mux2_1 _3581_ (.A0(\tms1x00.RAM[58][1] ),
    .A1(_1672_),
    .S(_1670_),
    .X(_1673_));
 sky130_fd_sc_hd__clkbuf_1 _3582_ (.A(_1673_),
    .X(_0352_));
 sky130_fd_sc_hd__buf_2 _3583_ (.A(_1129_),
    .X(_1674_));
 sky130_fd_sc_hd__mux2_1 _3584_ (.A0(\tms1x00.RAM[58][2] ),
    .A1(_1674_),
    .S(_1670_),
    .X(_1675_));
 sky130_fd_sc_hd__clkbuf_1 _3585_ (.A(_1675_),
    .X(_0353_));
 sky130_fd_sc_hd__clkbuf_4 _3586_ (.A(_1224_),
    .X(_1676_));
 sky130_fd_sc_hd__mux2_1 _3587_ (.A0(\tms1x00.RAM[58][3] ),
    .A1(_1676_),
    .S(_1670_),
    .X(_1677_));
 sky130_fd_sc_hd__clkbuf_1 _3588_ (.A(_1677_),
    .X(_0354_));
 sky130_fd_sc_hd__nor2_2 _3589_ (.A(_1261_),
    .B(_1284_),
    .Y(_1678_));
 sky130_fd_sc_hd__mux2_1 _3590_ (.A0(\tms1x00.RAM[57][0] ),
    .A1(_1669_),
    .S(_1678_),
    .X(_1679_));
 sky130_fd_sc_hd__clkbuf_1 _3591_ (.A(_1679_),
    .X(_0355_));
 sky130_fd_sc_hd__mux2_1 _3592_ (.A0(\tms1x00.RAM[57][1] ),
    .A1(_1672_),
    .S(_1678_),
    .X(_1680_));
 sky130_fd_sc_hd__clkbuf_1 _3593_ (.A(_1680_),
    .X(_0356_));
 sky130_fd_sc_hd__mux2_1 _3594_ (.A0(\tms1x00.RAM[57][2] ),
    .A1(_1674_),
    .S(_1678_),
    .X(_1681_));
 sky130_fd_sc_hd__clkbuf_1 _3595_ (.A(_1681_),
    .X(_0357_));
 sky130_fd_sc_hd__mux2_1 _3596_ (.A0(\tms1x00.RAM[57][3] ),
    .A1(_1676_),
    .S(_1678_),
    .X(_1682_));
 sky130_fd_sc_hd__clkbuf_1 _3597_ (.A(_1682_),
    .X(_0358_));
 sky130_fd_sc_hd__nor2_2 _3598_ (.A(_1284_),
    .B(_1303_),
    .Y(_1683_));
 sky130_fd_sc_hd__mux2_1 _3599_ (.A0(\tms1x00.RAM[56][0] ),
    .A1(_1669_),
    .S(_1683_),
    .X(_1684_));
 sky130_fd_sc_hd__clkbuf_1 _3600_ (.A(_1684_),
    .X(_0359_));
 sky130_fd_sc_hd__mux2_1 _3601_ (.A0(\tms1x00.RAM[56][1] ),
    .A1(_1672_),
    .S(_1683_),
    .X(_1685_));
 sky130_fd_sc_hd__clkbuf_1 _3602_ (.A(_1685_),
    .X(_0360_));
 sky130_fd_sc_hd__mux2_1 _3603_ (.A0(\tms1x00.RAM[56][2] ),
    .A1(_1674_),
    .S(_1683_),
    .X(_1686_));
 sky130_fd_sc_hd__clkbuf_1 _3604_ (.A(_1686_),
    .X(_0361_));
 sky130_fd_sc_hd__mux2_1 _3605_ (.A0(\tms1x00.RAM[56][3] ),
    .A1(_1676_),
    .S(_1683_),
    .X(_1687_));
 sky130_fd_sc_hd__clkbuf_1 _3606_ (.A(_1687_),
    .X(_0362_));
 sky130_fd_sc_hd__nor2_2 _3607_ (.A(_1284_),
    .B(_1310_),
    .Y(_1688_));
 sky130_fd_sc_hd__mux2_1 _3608_ (.A0(\tms1x00.RAM[55][0] ),
    .A1(_1669_),
    .S(_1688_),
    .X(_1689_));
 sky130_fd_sc_hd__clkbuf_1 _3609_ (.A(_1689_),
    .X(_0363_));
 sky130_fd_sc_hd__mux2_1 _3610_ (.A0(\tms1x00.RAM[55][1] ),
    .A1(_1672_),
    .S(_1688_),
    .X(_1690_));
 sky130_fd_sc_hd__clkbuf_1 _3611_ (.A(_1690_),
    .X(_0364_));
 sky130_fd_sc_hd__mux2_1 _3612_ (.A0(\tms1x00.RAM[55][2] ),
    .A1(_1674_),
    .S(_1688_),
    .X(_1691_));
 sky130_fd_sc_hd__clkbuf_1 _3613_ (.A(_1691_),
    .X(_0365_));
 sky130_fd_sc_hd__mux2_1 _3614_ (.A0(\tms1x00.RAM[55][3] ),
    .A1(_1676_),
    .S(_1688_),
    .X(_1692_));
 sky130_fd_sc_hd__clkbuf_1 _3615_ (.A(_1692_),
    .X(_0366_));
 sky130_fd_sc_hd__or2_2 _3616_ (.A(_1267_),
    .B(_1283_),
    .X(_1693_));
 sky130_fd_sc_hd__mux2_1 _3617_ (.A0(_1585_),
    .A1(\tms1x00.RAM[63][0] ),
    .S(_1693_),
    .X(_1694_));
 sky130_fd_sc_hd__clkbuf_1 _3618_ (.A(_1694_),
    .X(_0367_));
 sky130_fd_sc_hd__mux2_1 _3619_ (.A0(_1588_),
    .A1(\tms1x00.RAM[63][1] ),
    .S(_1693_),
    .X(_1695_));
 sky130_fd_sc_hd__clkbuf_1 _3620_ (.A(_1695_),
    .X(_0368_));
 sky130_fd_sc_hd__mux2_1 _3621_ (.A0(_1590_),
    .A1(\tms1x00.RAM[63][2] ),
    .S(_1693_),
    .X(_1696_));
 sky130_fd_sc_hd__clkbuf_1 _3622_ (.A(_1696_),
    .X(_0369_));
 sky130_fd_sc_hd__mux2_1 _3623_ (.A0(_1592_),
    .A1(\tms1x00.RAM[63][3] ),
    .S(_1693_),
    .X(_1697_));
 sky130_fd_sc_hd__clkbuf_1 _3624_ (.A(_1697_),
    .X(_0370_));
 sky130_fd_sc_hd__or2_2 _3625_ (.A(_1284_),
    .B(_1396_),
    .X(_1698_));
 sky130_fd_sc_hd__mux2_1 _3626_ (.A0(_1585_),
    .A1(\tms1x00.RAM[62][0] ),
    .S(_1698_),
    .X(_1699_));
 sky130_fd_sc_hd__clkbuf_1 _3627_ (.A(_1699_),
    .X(_0371_));
 sky130_fd_sc_hd__mux2_1 _3628_ (.A0(_1588_),
    .A1(\tms1x00.RAM[62][1] ),
    .S(_1698_),
    .X(_1700_));
 sky130_fd_sc_hd__clkbuf_1 _3629_ (.A(_1700_),
    .X(_0372_));
 sky130_fd_sc_hd__mux2_1 _3630_ (.A0(_1590_),
    .A1(\tms1x00.RAM[62][2] ),
    .S(_1698_),
    .X(_1701_));
 sky130_fd_sc_hd__clkbuf_1 _3631_ (.A(_1701_),
    .X(_0373_));
 sky130_fd_sc_hd__mux2_1 _3632_ (.A0(_1592_),
    .A1(\tms1x00.RAM[62][3] ),
    .S(_1698_),
    .X(_1702_));
 sky130_fd_sc_hd__clkbuf_1 _3633_ (.A(_1702_),
    .X(_0374_));
 sky130_fd_sc_hd__clkbuf_4 _3634_ (.A(_0911_),
    .X(_1703_));
 sky130_fd_sc_hd__or2_2 _3635_ (.A(_0917_),
    .B(_1283_),
    .X(_1704_));
 sky130_fd_sc_hd__mux2_1 _3636_ (.A0(_1703_),
    .A1(\tms1x00.RAM[61][0] ),
    .S(_1704_),
    .X(_1705_));
 sky130_fd_sc_hd__clkbuf_1 _3637_ (.A(_1705_),
    .X(_0375_));
 sky130_fd_sc_hd__buf_2 _3638_ (.A(_1034_),
    .X(_1706_));
 sky130_fd_sc_hd__mux2_1 _3639_ (.A0(_1706_),
    .A1(\tms1x00.RAM[61][1] ),
    .S(_1704_),
    .X(_1707_));
 sky130_fd_sc_hd__clkbuf_1 _3640_ (.A(_1707_),
    .X(_0376_));
 sky130_fd_sc_hd__buf_2 _3641_ (.A(_1129_),
    .X(_1708_));
 sky130_fd_sc_hd__mux2_1 _3642_ (.A0(_1708_),
    .A1(\tms1x00.RAM[61][2] ),
    .S(_1704_),
    .X(_1709_));
 sky130_fd_sc_hd__clkbuf_1 _3643_ (.A(_1709_),
    .X(_0377_));
 sky130_fd_sc_hd__clkbuf_4 _3644_ (.A(_1224_),
    .X(_1710_));
 sky130_fd_sc_hd__mux2_1 _3645_ (.A0(_1710_),
    .A1(\tms1x00.RAM[61][3] ),
    .S(_1704_),
    .X(_1711_));
 sky130_fd_sc_hd__clkbuf_1 _3646_ (.A(_1711_),
    .X(_0378_));
 sky130_fd_sc_hd__or2_2 _3647_ (.A(_1283_),
    .B(_1409_),
    .X(_1712_));
 sky130_fd_sc_hd__mux2_1 _3648_ (.A0(_1703_),
    .A1(\tms1x00.RAM[60][0] ),
    .S(_1712_),
    .X(_1713_));
 sky130_fd_sc_hd__clkbuf_1 _3649_ (.A(_1713_),
    .X(_0379_));
 sky130_fd_sc_hd__mux2_1 _3650_ (.A0(_1706_),
    .A1(\tms1x00.RAM[60][1] ),
    .S(_1712_),
    .X(_1714_));
 sky130_fd_sc_hd__clkbuf_1 _3651_ (.A(_1714_),
    .X(_0380_));
 sky130_fd_sc_hd__mux2_1 _3652_ (.A0(_1708_),
    .A1(\tms1x00.RAM[60][2] ),
    .S(_1712_),
    .X(_1715_));
 sky130_fd_sc_hd__clkbuf_1 _3653_ (.A(_1715_),
    .X(_0381_));
 sky130_fd_sc_hd__mux2_1 _3654_ (.A0(_1710_),
    .A1(\tms1x00.RAM[60][3] ),
    .S(_1712_),
    .X(_1716_));
 sky130_fd_sc_hd__clkbuf_1 _3655_ (.A(_1716_),
    .X(_0382_));
 sky130_fd_sc_hd__or2_2 _3656_ (.A(_1229_),
    .B(_1236_),
    .X(_1717_));
 sky130_fd_sc_hd__mux2_1 _3657_ (.A0(_1703_),
    .A1(\tms1x00.RAM[67][0] ),
    .S(_1717_),
    .X(_1718_));
 sky130_fd_sc_hd__clkbuf_1 _3658_ (.A(_1718_),
    .X(_0383_));
 sky130_fd_sc_hd__mux2_1 _3659_ (.A0(_1706_),
    .A1(\tms1x00.RAM[67][1] ),
    .S(_1717_),
    .X(_1719_));
 sky130_fd_sc_hd__clkbuf_1 _3660_ (.A(_1719_),
    .X(_0384_));
 sky130_fd_sc_hd__mux2_1 _3661_ (.A0(_1708_),
    .A1(\tms1x00.RAM[67][2] ),
    .S(_1717_),
    .X(_1720_));
 sky130_fd_sc_hd__clkbuf_1 _3662_ (.A(_1720_),
    .X(_0385_));
 sky130_fd_sc_hd__mux2_1 _3663_ (.A0(_1710_),
    .A1(\tms1x00.RAM[67][3] ),
    .S(_1717_),
    .X(_1721_));
 sky130_fd_sc_hd__clkbuf_1 _3664_ (.A(_1721_),
    .X(_0386_));
 sky130_fd_sc_hd__or2_2 _3665_ (.A(_1237_),
    .B(_1273_),
    .X(_1722_));
 sky130_fd_sc_hd__mux2_1 _3666_ (.A0(_1703_),
    .A1(\tms1x00.RAM[66][0] ),
    .S(_1722_),
    .X(_1723_));
 sky130_fd_sc_hd__clkbuf_1 _3667_ (.A(_1723_),
    .X(_0387_));
 sky130_fd_sc_hd__mux2_1 _3668_ (.A0(_1706_),
    .A1(\tms1x00.RAM[66][1] ),
    .S(_1722_),
    .X(_1724_));
 sky130_fd_sc_hd__clkbuf_1 _3669_ (.A(_1724_),
    .X(_0388_));
 sky130_fd_sc_hd__mux2_1 _3670_ (.A0(_1708_),
    .A1(\tms1x00.RAM[66][2] ),
    .S(_1722_),
    .X(_1725_));
 sky130_fd_sc_hd__clkbuf_1 _3671_ (.A(_1725_),
    .X(_0389_));
 sky130_fd_sc_hd__mux2_1 _3672_ (.A0(_1710_),
    .A1(\tms1x00.RAM[66][3] ),
    .S(_1722_),
    .X(_1726_));
 sky130_fd_sc_hd__clkbuf_1 _3673_ (.A(_1726_),
    .X(_0390_));
 sky130_fd_sc_hd__or2_2 _3674_ (.A(_1236_),
    .B(_1251_),
    .X(_1727_));
 sky130_fd_sc_hd__mux2_1 _3675_ (.A0(_1703_),
    .A1(\tms1x00.RAM[65][0] ),
    .S(_1727_),
    .X(_1728_));
 sky130_fd_sc_hd__clkbuf_1 _3676_ (.A(_1728_),
    .X(_0391_));
 sky130_fd_sc_hd__mux2_1 _3677_ (.A0(_1706_),
    .A1(\tms1x00.RAM[65][1] ),
    .S(_1727_),
    .X(_1729_));
 sky130_fd_sc_hd__clkbuf_1 _3678_ (.A(_1729_),
    .X(_0392_));
 sky130_fd_sc_hd__mux2_1 _3679_ (.A0(_1708_),
    .A1(\tms1x00.RAM[65][2] ),
    .S(_1727_),
    .X(_1730_));
 sky130_fd_sc_hd__clkbuf_1 _3680_ (.A(_1730_),
    .X(_0393_));
 sky130_fd_sc_hd__mux2_1 _3681_ (.A0(_1710_),
    .A1(\tms1x00.RAM[65][3] ),
    .S(_1727_),
    .X(_1731_));
 sky130_fd_sc_hd__clkbuf_1 _3682_ (.A(_1731_),
    .X(_0394_));
 sky130_fd_sc_hd__or2_2 _3683_ (.A(_1236_),
    .B(_1345_),
    .X(_1732_));
 sky130_fd_sc_hd__mux2_1 _3684_ (.A0(_1703_),
    .A1(\tms1x00.RAM[64][0] ),
    .S(_1732_),
    .X(_1733_));
 sky130_fd_sc_hd__clkbuf_1 _3685_ (.A(_1733_),
    .X(_0395_));
 sky130_fd_sc_hd__mux2_1 _3686_ (.A0(_1706_),
    .A1(\tms1x00.RAM[64][1] ),
    .S(_1732_),
    .X(_1734_));
 sky130_fd_sc_hd__clkbuf_1 _3687_ (.A(_1734_),
    .X(_0396_));
 sky130_fd_sc_hd__mux2_1 _3688_ (.A0(_1708_),
    .A1(\tms1x00.RAM[64][2] ),
    .S(_1732_),
    .X(_1735_));
 sky130_fd_sc_hd__clkbuf_1 _3689_ (.A(_1735_),
    .X(_0397_));
 sky130_fd_sc_hd__mux2_1 _3690_ (.A0(_1710_),
    .A1(\tms1x00.RAM[64][3] ),
    .S(_1732_),
    .X(_1736_));
 sky130_fd_sc_hd__clkbuf_1 _3691_ (.A(_1736_),
    .X(_0398_));
 sky130_fd_sc_hd__nor2_2 _3692_ (.A(_1237_),
    .B(_1303_),
    .Y(_1737_));
 sky130_fd_sc_hd__mux2_1 _3693_ (.A0(\tms1x00.RAM[72][0] ),
    .A1(_1669_),
    .S(_1737_),
    .X(_1738_));
 sky130_fd_sc_hd__clkbuf_1 _3694_ (.A(_1738_),
    .X(_0399_));
 sky130_fd_sc_hd__mux2_1 _3695_ (.A0(\tms1x00.RAM[72][1] ),
    .A1(_1672_),
    .S(_1737_),
    .X(_1739_));
 sky130_fd_sc_hd__clkbuf_1 _3696_ (.A(_1739_),
    .X(_0400_));
 sky130_fd_sc_hd__mux2_1 _3697_ (.A0(\tms1x00.RAM[72][2] ),
    .A1(_1674_),
    .S(_1737_),
    .X(_1740_));
 sky130_fd_sc_hd__clkbuf_1 _3698_ (.A(_1740_),
    .X(_0401_));
 sky130_fd_sc_hd__mux2_1 _3699_ (.A0(\tms1x00.RAM[72][3] ),
    .A1(_1676_),
    .S(_1737_),
    .X(_1741_));
 sky130_fd_sc_hd__clkbuf_1 _3700_ (.A(_1741_),
    .X(_0402_));
 sky130_fd_sc_hd__nor2_2 _3701_ (.A(_1237_),
    .B(_1310_),
    .Y(_1742_));
 sky130_fd_sc_hd__mux2_1 _3702_ (.A0(\tms1x00.RAM[71][0] ),
    .A1(_1669_),
    .S(_1742_),
    .X(_1743_));
 sky130_fd_sc_hd__clkbuf_1 _3703_ (.A(_1743_),
    .X(_0403_));
 sky130_fd_sc_hd__mux2_1 _3704_ (.A0(\tms1x00.RAM[71][1] ),
    .A1(_1672_),
    .S(_1742_),
    .X(_1744_));
 sky130_fd_sc_hd__clkbuf_1 _3705_ (.A(_1744_),
    .X(_0404_));
 sky130_fd_sc_hd__mux2_1 _3706_ (.A0(\tms1x00.RAM[71][2] ),
    .A1(_1674_),
    .S(_1742_),
    .X(_1745_));
 sky130_fd_sc_hd__clkbuf_1 _3707_ (.A(_1745_),
    .X(_0405_));
 sky130_fd_sc_hd__mux2_1 _3708_ (.A0(\tms1x00.RAM[71][3] ),
    .A1(_1676_),
    .S(_1742_),
    .X(_1746_));
 sky130_fd_sc_hd__clkbuf_1 _3709_ (.A(_1746_),
    .X(_0406_));
 sky130_fd_sc_hd__nor2_2 _3710_ (.A(_1237_),
    .B(_1317_),
    .Y(_1747_));
 sky130_fd_sc_hd__mux2_1 _3711_ (.A0(\tms1x00.RAM[70][0] ),
    .A1(_1669_),
    .S(_1747_),
    .X(_1748_));
 sky130_fd_sc_hd__clkbuf_1 _3712_ (.A(_1748_),
    .X(_0407_));
 sky130_fd_sc_hd__mux2_1 _3713_ (.A0(\tms1x00.RAM[70][1] ),
    .A1(_1672_),
    .S(_1747_),
    .X(_1749_));
 sky130_fd_sc_hd__clkbuf_1 _3714_ (.A(_1749_),
    .X(_0408_));
 sky130_fd_sc_hd__mux2_1 _3715_ (.A0(\tms1x00.RAM[70][2] ),
    .A1(_1674_),
    .S(_1747_),
    .X(_1750_));
 sky130_fd_sc_hd__clkbuf_1 _3716_ (.A(_1750_),
    .X(_0409_));
 sky130_fd_sc_hd__mux2_1 _3717_ (.A0(\tms1x00.RAM[70][3] ),
    .A1(_1676_),
    .S(_1747_),
    .X(_1751_));
 sky130_fd_sc_hd__clkbuf_1 _3718_ (.A(_1751_),
    .X(_0410_));
 sky130_fd_sc_hd__nor2_2 _3719_ (.A(_1317_),
    .B(_1344_),
    .Y(_1752_));
 sky130_fd_sc_hd__mux2_1 _3720_ (.A0(\tms1x00.RAM[6][0] ),
    .A1(_1669_),
    .S(_1752_),
    .X(_1753_));
 sky130_fd_sc_hd__clkbuf_1 _3721_ (.A(_1753_),
    .X(_0411_));
 sky130_fd_sc_hd__mux2_1 _3722_ (.A0(\tms1x00.RAM[6][1] ),
    .A1(_1672_),
    .S(_1752_),
    .X(_1754_));
 sky130_fd_sc_hd__clkbuf_1 _3723_ (.A(_1754_),
    .X(_0412_));
 sky130_fd_sc_hd__mux2_1 _3724_ (.A0(\tms1x00.RAM[6][2] ),
    .A1(_1674_),
    .S(_1752_),
    .X(_1755_));
 sky130_fd_sc_hd__clkbuf_1 _3725_ (.A(_1755_),
    .X(_0413_));
 sky130_fd_sc_hd__mux2_1 _3726_ (.A0(\tms1x00.RAM[6][3] ),
    .A1(_1676_),
    .S(_1752_),
    .X(_1756_));
 sky130_fd_sc_hd__clkbuf_1 _3727_ (.A(_1756_),
    .X(_0414_));
 sky130_fd_sc_hd__nor2_2 _3728_ (.A(_1237_),
    .B(_1337_),
    .Y(_1757_));
 sky130_fd_sc_hd__mux2_1 _3729_ (.A0(\tms1x00.RAM[68][0] ),
    .A1(_1669_),
    .S(_1757_),
    .X(_1758_));
 sky130_fd_sc_hd__clkbuf_1 _3730_ (.A(_1758_),
    .X(_0415_));
 sky130_fd_sc_hd__mux2_1 _3731_ (.A0(\tms1x00.RAM[68][1] ),
    .A1(_1672_),
    .S(_1757_),
    .X(_1759_));
 sky130_fd_sc_hd__clkbuf_1 _3732_ (.A(_1759_),
    .X(_0416_));
 sky130_fd_sc_hd__mux2_1 _3733_ (.A0(\tms1x00.RAM[68][2] ),
    .A1(_1674_),
    .S(_1757_),
    .X(_1760_));
 sky130_fd_sc_hd__clkbuf_1 _3734_ (.A(_1760_),
    .X(_0417_));
 sky130_fd_sc_hd__mux2_1 _3735_ (.A0(\tms1x00.RAM[68][3] ),
    .A1(_1676_),
    .S(_1757_),
    .X(_1761_));
 sky130_fd_sc_hd__clkbuf_1 _3736_ (.A(_1761_),
    .X(_0418_));
 sky130_fd_sc_hd__or2_2 _3737_ (.A(_1236_),
    .B(_1409_),
    .X(_1762_));
 sky130_fd_sc_hd__mux2_1 _3738_ (.A0(_1703_),
    .A1(\tms1x00.RAM[76][0] ),
    .S(_1762_),
    .X(_1763_));
 sky130_fd_sc_hd__clkbuf_1 _3739_ (.A(_1763_),
    .X(_0419_));
 sky130_fd_sc_hd__mux2_1 _3740_ (.A0(_1706_),
    .A1(\tms1x00.RAM[76][1] ),
    .S(_1762_),
    .X(_1764_));
 sky130_fd_sc_hd__clkbuf_1 _3741_ (.A(_1764_),
    .X(_0420_));
 sky130_fd_sc_hd__mux2_1 _3742_ (.A0(_1708_),
    .A1(\tms1x00.RAM[76][2] ),
    .S(_1762_),
    .X(_1765_));
 sky130_fd_sc_hd__clkbuf_1 _3743_ (.A(_1765_),
    .X(_0421_));
 sky130_fd_sc_hd__mux2_1 _3744_ (.A0(_1710_),
    .A1(\tms1x00.RAM[76][3] ),
    .S(_1762_),
    .X(_1766_));
 sky130_fd_sc_hd__clkbuf_1 _3745_ (.A(_1766_),
    .X(_0422_));
 sky130_fd_sc_hd__nor2_2 _3746_ (.A(_1237_),
    .B(_1286_),
    .Y(_1767_));
 sky130_fd_sc_hd__mux2_1 _3747_ (.A0(\tms1x00.RAM[75][0] ),
    .A1(_1669_),
    .S(_1767_),
    .X(_1768_));
 sky130_fd_sc_hd__clkbuf_1 _3748_ (.A(_1768_),
    .X(_0423_));
 sky130_fd_sc_hd__mux2_1 _3749_ (.A0(\tms1x00.RAM[75][1] ),
    .A1(_1672_),
    .S(_1767_),
    .X(_1769_));
 sky130_fd_sc_hd__clkbuf_1 _3750_ (.A(_1769_),
    .X(_0424_));
 sky130_fd_sc_hd__mux2_1 _3751_ (.A0(\tms1x00.RAM[75][2] ),
    .A1(_1674_),
    .S(_1767_),
    .X(_1770_));
 sky130_fd_sc_hd__clkbuf_1 _3752_ (.A(_1770_),
    .X(_0425_));
 sky130_fd_sc_hd__mux2_1 _3753_ (.A0(\tms1x00.RAM[75][3] ),
    .A1(_1676_),
    .S(_1767_),
    .X(_1771_));
 sky130_fd_sc_hd__clkbuf_1 _3754_ (.A(_1771_),
    .X(_0426_));
 sky130_fd_sc_hd__clkbuf_4 _3755_ (.A(_0911_),
    .X(_1772_));
 sky130_fd_sc_hd__nor2_2 _3756_ (.A(_1237_),
    .B(_1403_),
    .Y(_1773_));
 sky130_fd_sc_hd__mux2_1 _3757_ (.A0(\tms1x00.RAM[74][0] ),
    .A1(_1772_),
    .S(_1773_),
    .X(_1774_));
 sky130_fd_sc_hd__clkbuf_1 _3758_ (.A(_1774_),
    .X(_0427_));
 sky130_fd_sc_hd__clkbuf_4 _3759_ (.A(_1034_),
    .X(_1775_));
 sky130_fd_sc_hd__mux2_1 _3760_ (.A0(\tms1x00.RAM[74][1] ),
    .A1(_1775_),
    .S(_1773_),
    .X(_1776_));
 sky130_fd_sc_hd__clkbuf_1 _3761_ (.A(_1776_),
    .X(_0428_));
 sky130_fd_sc_hd__clkbuf_4 _3762_ (.A(_1129_),
    .X(_1777_));
 sky130_fd_sc_hd__mux2_1 _3763_ (.A0(\tms1x00.RAM[74][2] ),
    .A1(_1777_),
    .S(_1773_),
    .X(_1778_));
 sky130_fd_sc_hd__clkbuf_1 _3764_ (.A(_1778_),
    .X(_0429_));
 sky130_fd_sc_hd__clkbuf_4 _3765_ (.A(_1224_),
    .X(_1779_));
 sky130_fd_sc_hd__mux2_1 _3766_ (.A0(\tms1x00.RAM[74][3] ),
    .A1(_1779_),
    .S(_1773_),
    .X(_1780_));
 sky130_fd_sc_hd__clkbuf_1 _3767_ (.A(_1780_),
    .X(_0430_));
 sky130_fd_sc_hd__nor2_2 _3768_ (.A(_1237_),
    .B(_1261_),
    .Y(_1781_));
 sky130_fd_sc_hd__mux2_1 _3769_ (.A0(\tms1x00.RAM[73][0] ),
    .A1(_1772_),
    .S(_1781_),
    .X(_1782_));
 sky130_fd_sc_hd__clkbuf_1 _3770_ (.A(_1782_),
    .X(_0431_));
 sky130_fd_sc_hd__mux2_1 _3771_ (.A0(\tms1x00.RAM[73][1] ),
    .A1(_1775_),
    .S(_1781_),
    .X(_1783_));
 sky130_fd_sc_hd__clkbuf_1 _3772_ (.A(_1783_),
    .X(_0432_));
 sky130_fd_sc_hd__mux2_1 _3773_ (.A0(\tms1x00.RAM[73][2] ),
    .A1(_1777_),
    .S(_1781_),
    .X(_1784_));
 sky130_fd_sc_hd__clkbuf_1 _3774_ (.A(_1784_),
    .X(_0433_));
 sky130_fd_sc_hd__mux2_1 _3775_ (.A0(\tms1x00.RAM[73][3] ),
    .A1(_1779_),
    .S(_1781_),
    .X(_1785_));
 sky130_fd_sc_hd__clkbuf_1 _3776_ (.A(_1785_),
    .X(_0434_));
 sky130_fd_sc_hd__or2_2 _3777_ (.A(_1258_),
    .B(_1345_),
    .X(_1786_));
 sky130_fd_sc_hd__mux2_1 _3778_ (.A0(_1703_),
    .A1(\tms1x00.RAM[80][0] ),
    .S(_1786_),
    .X(_1787_));
 sky130_fd_sc_hd__clkbuf_1 _3779_ (.A(_1787_),
    .X(_0435_));
 sky130_fd_sc_hd__mux2_1 _3780_ (.A0(_1706_),
    .A1(\tms1x00.RAM[80][1] ),
    .S(_1786_),
    .X(_1788_));
 sky130_fd_sc_hd__clkbuf_1 _3781_ (.A(_1788_),
    .X(_0436_));
 sky130_fd_sc_hd__mux2_1 _3782_ (.A0(_1708_),
    .A1(\tms1x00.RAM[80][2] ),
    .S(_1786_),
    .X(_1789_));
 sky130_fd_sc_hd__clkbuf_1 _3783_ (.A(_1789_),
    .X(_0437_));
 sky130_fd_sc_hd__mux2_1 _3784_ (.A0(_1710_),
    .A1(\tms1x00.RAM[80][3] ),
    .S(_1786_),
    .X(_1790_));
 sky130_fd_sc_hd__clkbuf_1 _3785_ (.A(_1790_),
    .X(_0438_));
 sky130_fd_sc_hd__nor2_2 _3786_ (.A(_1310_),
    .B(_1344_),
    .Y(_1791_));
 sky130_fd_sc_hd__mux2_1 _3787_ (.A0(\tms1x00.RAM[7][0] ),
    .A1(_1772_),
    .S(_1791_),
    .X(_1792_));
 sky130_fd_sc_hd__clkbuf_1 _3788_ (.A(_1792_),
    .X(_0439_));
 sky130_fd_sc_hd__mux2_1 _3789_ (.A0(\tms1x00.RAM[7][1] ),
    .A1(_1775_),
    .S(_1791_),
    .X(_1793_));
 sky130_fd_sc_hd__clkbuf_1 _3790_ (.A(_1793_),
    .X(_0440_));
 sky130_fd_sc_hd__mux2_1 _3791_ (.A0(\tms1x00.RAM[7][2] ),
    .A1(_1777_),
    .S(_1791_),
    .X(_1794_));
 sky130_fd_sc_hd__clkbuf_1 _3792_ (.A(_1794_),
    .X(_0441_));
 sky130_fd_sc_hd__mux2_1 _3793_ (.A0(\tms1x00.RAM[7][3] ),
    .A1(_1779_),
    .S(_1791_),
    .X(_1795_));
 sky130_fd_sc_hd__clkbuf_1 _3794_ (.A(_1795_),
    .X(_0442_));
 sky130_fd_sc_hd__or2_2 _3795_ (.A(_1236_),
    .B(_1396_),
    .X(_1796_));
 sky130_fd_sc_hd__mux2_1 _3796_ (.A0(_1703_),
    .A1(\tms1x00.RAM[78][0] ),
    .S(_1796_),
    .X(_1797_));
 sky130_fd_sc_hd__clkbuf_1 _3797_ (.A(_1797_),
    .X(_0443_));
 sky130_fd_sc_hd__mux2_1 _3798_ (.A0(_1706_),
    .A1(\tms1x00.RAM[78][1] ),
    .S(_1796_),
    .X(_1798_));
 sky130_fd_sc_hd__clkbuf_1 _3799_ (.A(_1798_),
    .X(_0444_));
 sky130_fd_sc_hd__mux2_1 _3800_ (.A0(_1708_),
    .A1(\tms1x00.RAM[78][2] ),
    .S(_1796_),
    .X(_1799_));
 sky130_fd_sc_hd__clkbuf_1 _3801_ (.A(_1799_),
    .X(_0445_));
 sky130_fd_sc_hd__mux2_1 _3802_ (.A0(_1710_),
    .A1(\tms1x00.RAM[78][3] ),
    .S(_1796_),
    .X(_1800_));
 sky130_fd_sc_hd__clkbuf_1 _3803_ (.A(_1800_),
    .X(_0446_));
 sky130_fd_sc_hd__or2_2 _3804_ (.A(_0917_),
    .B(_1236_),
    .X(_1801_));
 sky130_fd_sc_hd__mux2_1 _3805_ (.A0(_1703_),
    .A1(\tms1x00.RAM[77][0] ),
    .S(_1801_),
    .X(_1802_));
 sky130_fd_sc_hd__clkbuf_1 _3806_ (.A(_1802_),
    .X(_0447_));
 sky130_fd_sc_hd__mux2_1 _3807_ (.A0(_1706_),
    .A1(\tms1x00.RAM[77][1] ),
    .S(_1801_),
    .X(_1803_));
 sky130_fd_sc_hd__clkbuf_1 _3808_ (.A(_1803_),
    .X(_0448_));
 sky130_fd_sc_hd__mux2_1 _3809_ (.A0(_1708_),
    .A1(\tms1x00.RAM[77][2] ),
    .S(_1801_),
    .X(_1804_));
 sky130_fd_sc_hd__clkbuf_1 _3810_ (.A(_1804_),
    .X(_0449_));
 sky130_fd_sc_hd__mux2_1 _3811_ (.A0(_1710_),
    .A1(\tms1x00.RAM[77][3] ),
    .S(_1801_),
    .X(_1805_));
 sky130_fd_sc_hd__clkbuf_1 _3812_ (.A(_1805_),
    .X(_0450_));
 sky130_fd_sc_hd__nor2_2 _3813_ (.A(_1240_),
    .B(_1258_),
    .Y(_1806_));
 sky130_fd_sc_hd__mux2_1 _3814_ (.A0(\tms1x00.RAM[85][0] ),
    .A1(_1772_),
    .S(_1806_),
    .X(_1807_));
 sky130_fd_sc_hd__clkbuf_1 _3815_ (.A(_1807_),
    .X(_0451_));
 sky130_fd_sc_hd__mux2_1 _3816_ (.A0(\tms1x00.RAM[85][1] ),
    .A1(_1775_),
    .S(_1806_),
    .X(_1808_));
 sky130_fd_sc_hd__clkbuf_1 _3817_ (.A(_1808_),
    .X(_0452_));
 sky130_fd_sc_hd__mux2_1 _3818_ (.A0(\tms1x00.RAM[85][2] ),
    .A1(_1777_),
    .S(_1806_),
    .X(_1809_));
 sky130_fd_sc_hd__clkbuf_1 _3819_ (.A(_1809_),
    .X(_0453_));
 sky130_fd_sc_hd__mux2_1 _3820_ (.A0(\tms1x00.RAM[85][3] ),
    .A1(_1779_),
    .S(_1806_),
    .X(_1810_));
 sky130_fd_sc_hd__clkbuf_1 _3821_ (.A(_1810_),
    .X(_0454_));
 sky130_fd_sc_hd__nor2_2 _3822_ (.A(_1258_),
    .B(_1337_),
    .Y(_1811_));
 sky130_fd_sc_hd__mux2_1 _3823_ (.A0(\tms1x00.RAM[84][0] ),
    .A1(_1772_),
    .S(_1811_),
    .X(_1812_));
 sky130_fd_sc_hd__clkbuf_1 _3824_ (.A(_1812_),
    .X(_0455_));
 sky130_fd_sc_hd__mux2_1 _3825_ (.A0(\tms1x00.RAM[84][1] ),
    .A1(_1775_),
    .S(_1811_),
    .X(_1813_));
 sky130_fd_sc_hd__clkbuf_1 _3826_ (.A(_1813_),
    .X(_0456_));
 sky130_fd_sc_hd__mux2_1 _3827_ (.A0(\tms1x00.RAM[84][2] ),
    .A1(_1777_),
    .S(_1811_),
    .X(_1814_));
 sky130_fd_sc_hd__clkbuf_1 _3828_ (.A(_1814_),
    .X(_0457_));
 sky130_fd_sc_hd__mux2_1 _3829_ (.A0(\tms1x00.RAM[84][3] ),
    .A1(_1779_),
    .S(_1811_),
    .X(_1815_));
 sky130_fd_sc_hd__clkbuf_1 _3830_ (.A(_1815_),
    .X(_0458_));
 sky130_fd_sc_hd__clkbuf_4 _3831_ (.A(_0911_),
    .X(_1816_));
 sky130_fd_sc_hd__or2_2 _3832_ (.A(_1229_),
    .B(_1257_),
    .X(_1817_));
 sky130_fd_sc_hd__mux2_1 _3833_ (.A0(_1816_),
    .A1(\tms1x00.RAM[83][0] ),
    .S(_1817_),
    .X(_1818_));
 sky130_fd_sc_hd__clkbuf_1 _3834_ (.A(_1818_),
    .X(_0459_));
 sky130_fd_sc_hd__clkbuf_4 _3835_ (.A(_1034_),
    .X(_1819_));
 sky130_fd_sc_hd__mux2_1 _3836_ (.A0(_1819_),
    .A1(\tms1x00.RAM[83][1] ),
    .S(_1817_),
    .X(_1820_));
 sky130_fd_sc_hd__clkbuf_1 _3837_ (.A(_1820_),
    .X(_0460_));
 sky130_fd_sc_hd__clkbuf_4 _3838_ (.A(_1129_),
    .X(_1821_));
 sky130_fd_sc_hd__mux2_1 _3839_ (.A0(_1821_),
    .A1(\tms1x00.RAM[83][2] ),
    .S(_1817_),
    .X(_1822_));
 sky130_fd_sc_hd__clkbuf_1 _3840_ (.A(_1822_),
    .X(_0461_));
 sky130_fd_sc_hd__clkbuf_4 _3841_ (.A(_1224_),
    .X(_1823_));
 sky130_fd_sc_hd__mux2_1 _3842_ (.A0(_1823_),
    .A1(\tms1x00.RAM[83][3] ),
    .S(_1817_),
    .X(_1824_));
 sky130_fd_sc_hd__clkbuf_1 _3843_ (.A(_1824_),
    .X(_0462_));
 sky130_fd_sc_hd__or2_2 _3844_ (.A(_1257_),
    .B(_1273_),
    .X(_1825_));
 sky130_fd_sc_hd__mux2_1 _3845_ (.A0(_1816_),
    .A1(\tms1x00.RAM[82][0] ),
    .S(_1825_),
    .X(_1826_));
 sky130_fd_sc_hd__clkbuf_1 _3846_ (.A(_1826_),
    .X(_0463_));
 sky130_fd_sc_hd__mux2_1 _3847_ (.A0(_1819_),
    .A1(\tms1x00.RAM[82][1] ),
    .S(_1825_),
    .X(_1827_));
 sky130_fd_sc_hd__clkbuf_1 _3848_ (.A(_1827_),
    .X(_0464_));
 sky130_fd_sc_hd__mux2_1 _3849_ (.A0(_1821_),
    .A1(\tms1x00.RAM[82][2] ),
    .S(_1825_),
    .X(_1828_));
 sky130_fd_sc_hd__clkbuf_1 _3850_ (.A(_1828_),
    .X(_0465_));
 sky130_fd_sc_hd__mux2_1 _3851_ (.A0(_1823_),
    .A1(\tms1x00.RAM[82][3] ),
    .S(_1825_),
    .X(_1829_));
 sky130_fd_sc_hd__clkbuf_1 _3852_ (.A(_1829_),
    .X(_0466_));
 sky130_fd_sc_hd__or2_2 _3853_ (.A(_1251_),
    .B(_1257_),
    .X(_1830_));
 sky130_fd_sc_hd__mux2_1 _3854_ (.A0(_1816_),
    .A1(\tms1x00.RAM[81][0] ),
    .S(_1830_),
    .X(_1831_));
 sky130_fd_sc_hd__clkbuf_1 _3855_ (.A(_1831_),
    .X(_0467_));
 sky130_fd_sc_hd__mux2_1 _3856_ (.A0(_1819_),
    .A1(\tms1x00.RAM[81][1] ),
    .S(_1830_),
    .X(_1832_));
 sky130_fd_sc_hd__clkbuf_1 _3857_ (.A(_1832_),
    .X(_0468_));
 sky130_fd_sc_hd__mux2_1 _3858_ (.A0(_1821_),
    .A1(\tms1x00.RAM[81][2] ),
    .S(_1830_),
    .X(_1833_));
 sky130_fd_sc_hd__clkbuf_1 _3859_ (.A(_1833_),
    .X(_0469_));
 sky130_fd_sc_hd__mux2_1 _3860_ (.A0(_1823_),
    .A1(\tms1x00.RAM[81][3] ),
    .S(_1830_),
    .X(_1834_));
 sky130_fd_sc_hd__clkbuf_1 _3861_ (.A(_1834_),
    .X(_0470_));
 sky130_fd_sc_hd__nor2_2 _3862_ (.A(_1258_),
    .B(_1317_),
    .Y(_1835_));
 sky130_fd_sc_hd__mux2_1 _3863_ (.A0(\tms1x00.RAM[86][0] ),
    .A1(_1772_),
    .S(_1835_),
    .X(_1836_));
 sky130_fd_sc_hd__clkbuf_1 _3864_ (.A(_1836_),
    .X(_0471_));
 sky130_fd_sc_hd__mux2_1 _3865_ (.A0(\tms1x00.RAM[86][1] ),
    .A1(_1775_),
    .S(_1835_),
    .X(_1837_));
 sky130_fd_sc_hd__clkbuf_1 _3866_ (.A(_1837_),
    .X(_0472_));
 sky130_fd_sc_hd__mux2_1 _3867_ (.A0(\tms1x00.RAM[86][2] ),
    .A1(_1777_),
    .S(_1835_),
    .X(_1838_));
 sky130_fd_sc_hd__clkbuf_1 _3868_ (.A(_1838_),
    .X(_0473_));
 sky130_fd_sc_hd__mux2_1 _3869_ (.A0(\tms1x00.RAM[86][3] ),
    .A1(_1779_),
    .S(_1835_),
    .X(_1839_));
 sky130_fd_sc_hd__clkbuf_1 _3870_ (.A(_1839_),
    .X(_0474_));
 sky130_fd_sc_hd__nor2_2 _3871_ (.A(_1303_),
    .B(_1344_),
    .Y(_1840_));
 sky130_fd_sc_hd__mux2_1 _3872_ (.A0(\tms1x00.RAM[8][0] ),
    .A1(_1772_),
    .S(_1840_),
    .X(_1841_));
 sky130_fd_sc_hd__clkbuf_1 _3873_ (.A(_1841_),
    .X(_0475_));
 sky130_fd_sc_hd__mux2_1 _3874_ (.A0(\tms1x00.RAM[8][1] ),
    .A1(_1775_),
    .S(_1840_),
    .X(_1842_));
 sky130_fd_sc_hd__clkbuf_1 _3875_ (.A(_1842_),
    .X(_0476_));
 sky130_fd_sc_hd__mux2_1 _3876_ (.A0(\tms1x00.RAM[8][2] ),
    .A1(_1777_),
    .S(_1840_),
    .X(_1843_));
 sky130_fd_sc_hd__clkbuf_1 _3877_ (.A(_1843_),
    .X(_0477_));
 sky130_fd_sc_hd__mux2_1 _3878_ (.A0(\tms1x00.RAM[8][3] ),
    .A1(_1779_),
    .S(_1840_),
    .X(_1844_));
 sky130_fd_sc_hd__clkbuf_1 _3879_ (.A(_1844_),
    .X(_0478_));
 sky130_fd_sc_hd__nor2_2 _3880_ (.A(_1258_),
    .B(_1303_),
    .Y(_1845_));
 sky130_fd_sc_hd__mux2_1 _3881_ (.A0(\tms1x00.RAM[88][0] ),
    .A1(_1772_),
    .S(_1845_),
    .X(_1846_));
 sky130_fd_sc_hd__clkbuf_1 _3882_ (.A(_1846_),
    .X(_0479_));
 sky130_fd_sc_hd__mux2_1 _3883_ (.A0(\tms1x00.RAM[88][1] ),
    .A1(_1775_),
    .S(_1845_),
    .X(_1847_));
 sky130_fd_sc_hd__clkbuf_1 _3884_ (.A(_1847_),
    .X(_0480_));
 sky130_fd_sc_hd__mux2_1 _3885_ (.A0(\tms1x00.RAM[88][2] ),
    .A1(_1777_),
    .S(_1845_),
    .X(_1848_));
 sky130_fd_sc_hd__clkbuf_1 _3886_ (.A(_1848_),
    .X(_0481_));
 sky130_fd_sc_hd__mux2_1 _3887_ (.A0(\tms1x00.RAM[88][3] ),
    .A1(_1779_),
    .S(_1845_),
    .X(_1849_));
 sky130_fd_sc_hd__clkbuf_1 _3888_ (.A(_1849_),
    .X(_0482_));
 sky130_fd_sc_hd__nor2_2 _3889_ (.A(_1258_),
    .B(_1310_),
    .Y(_1850_));
 sky130_fd_sc_hd__mux2_1 _3890_ (.A0(\tms1x00.RAM[87][0] ),
    .A1(_1772_),
    .S(_1850_),
    .X(_1851_));
 sky130_fd_sc_hd__clkbuf_1 _3891_ (.A(_1851_),
    .X(_0483_));
 sky130_fd_sc_hd__mux2_1 _3892_ (.A0(\tms1x00.RAM[87][1] ),
    .A1(_1775_),
    .S(_1850_),
    .X(_1852_));
 sky130_fd_sc_hd__clkbuf_1 _3893_ (.A(_1852_),
    .X(_0484_));
 sky130_fd_sc_hd__mux2_1 _3894_ (.A0(\tms1x00.RAM[87][2] ),
    .A1(_1777_),
    .S(_1850_),
    .X(_1853_));
 sky130_fd_sc_hd__clkbuf_1 _3895_ (.A(_1853_),
    .X(_0485_));
 sky130_fd_sc_hd__mux2_1 _3896_ (.A0(\tms1x00.RAM[87][3] ),
    .A1(_1779_),
    .S(_1850_),
    .X(_1854_));
 sky130_fd_sc_hd__clkbuf_1 _3897_ (.A(_1854_),
    .X(_0486_));
 sky130_fd_sc_hd__or2_2 _3898_ (.A(_1257_),
    .B(_1396_),
    .X(_1855_));
 sky130_fd_sc_hd__mux2_1 _3899_ (.A0(_1816_),
    .A1(\tms1x00.RAM[94][0] ),
    .S(_1855_),
    .X(_1856_));
 sky130_fd_sc_hd__clkbuf_1 _3900_ (.A(_1856_),
    .X(_0487_));
 sky130_fd_sc_hd__mux2_1 _3901_ (.A0(_1819_),
    .A1(\tms1x00.RAM[94][1] ),
    .S(_1855_),
    .X(_1857_));
 sky130_fd_sc_hd__clkbuf_1 _3902_ (.A(_1857_),
    .X(_0488_));
 sky130_fd_sc_hd__mux2_1 _3903_ (.A0(_1821_),
    .A1(\tms1x00.RAM[94][2] ),
    .S(_1855_),
    .X(_1858_));
 sky130_fd_sc_hd__clkbuf_1 _3904_ (.A(_1858_),
    .X(_0489_));
 sky130_fd_sc_hd__mux2_1 _3905_ (.A0(_1823_),
    .A1(\tms1x00.RAM[94][3] ),
    .S(_1855_),
    .X(_1859_));
 sky130_fd_sc_hd__clkbuf_1 _3906_ (.A(_1859_),
    .X(_0490_));
 sky130_fd_sc_hd__or2_2 _3907_ (.A(_0917_),
    .B(_1257_),
    .X(_1860_));
 sky130_fd_sc_hd__mux2_1 _3908_ (.A0(_1816_),
    .A1(\tms1x00.RAM[93][0] ),
    .S(_1860_),
    .X(_1861_));
 sky130_fd_sc_hd__clkbuf_1 _3909_ (.A(_1861_),
    .X(_0491_));
 sky130_fd_sc_hd__mux2_1 _3910_ (.A0(_1819_),
    .A1(\tms1x00.RAM[93][1] ),
    .S(_1860_),
    .X(_1862_));
 sky130_fd_sc_hd__clkbuf_1 _3911_ (.A(_1862_),
    .X(_0492_));
 sky130_fd_sc_hd__mux2_1 _3912_ (.A0(_1821_),
    .A1(\tms1x00.RAM[93][2] ),
    .S(_1860_),
    .X(_1863_));
 sky130_fd_sc_hd__clkbuf_1 _3913_ (.A(_1863_),
    .X(_0493_));
 sky130_fd_sc_hd__mux2_1 _3914_ (.A0(_1823_),
    .A1(\tms1x00.RAM[93][3] ),
    .S(_1860_),
    .X(_1864_));
 sky130_fd_sc_hd__clkbuf_1 _3915_ (.A(_1864_),
    .X(_0494_));
 sky130_fd_sc_hd__or2_2 _3916_ (.A(_1257_),
    .B(_1409_),
    .X(_1865_));
 sky130_fd_sc_hd__mux2_1 _3917_ (.A0(_1816_),
    .A1(\tms1x00.RAM[92][0] ),
    .S(_1865_),
    .X(_1866_));
 sky130_fd_sc_hd__clkbuf_1 _3918_ (.A(_1866_),
    .X(_0495_));
 sky130_fd_sc_hd__mux2_1 _3919_ (.A0(_1819_),
    .A1(\tms1x00.RAM[92][1] ),
    .S(_1865_),
    .X(_1867_));
 sky130_fd_sc_hd__clkbuf_1 _3920_ (.A(_1867_),
    .X(_0496_));
 sky130_fd_sc_hd__mux2_1 _3921_ (.A0(_1821_),
    .A1(\tms1x00.RAM[92][2] ),
    .S(_1865_),
    .X(_1868_));
 sky130_fd_sc_hd__clkbuf_1 _3922_ (.A(_1868_),
    .X(_0497_));
 sky130_fd_sc_hd__mux2_1 _3923_ (.A0(_1823_),
    .A1(\tms1x00.RAM[92][3] ),
    .S(_1865_),
    .X(_1869_));
 sky130_fd_sc_hd__clkbuf_1 _3924_ (.A(_1869_),
    .X(_0498_));
 sky130_fd_sc_hd__nor2_2 _3925_ (.A(_1258_),
    .B(_1286_),
    .Y(_1870_));
 sky130_fd_sc_hd__mux2_1 _3926_ (.A0(\tms1x00.RAM[91][0] ),
    .A1(_1772_),
    .S(_1870_),
    .X(_1871_));
 sky130_fd_sc_hd__clkbuf_1 _3927_ (.A(_1871_),
    .X(_0499_));
 sky130_fd_sc_hd__mux2_1 _3928_ (.A0(\tms1x00.RAM[91][1] ),
    .A1(_1775_),
    .S(_1870_),
    .X(_1872_));
 sky130_fd_sc_hd__clkbuf_1 _3929_ (.A(_1872_),
    .X(_0500_));
 sky130_fd_sc_hd__mux2_1 _3930_ (.A0(\tms1x00.RAM[91][2] ),
    .A1(_1777_),
    .S(_1870_),
    .X(_1873_));
 sky130_fd_sc_hd__clkbuf_1 _3931_ (.A(_1873_),
    .X(_0501_));
 sky130_fd_sc_hd__mux2_1 _3932_ (.A0(\tms1x00.RAM[91][3] ),
    .A1(_1779_),
    .S(_1870_),
    .X(_1874_));
 sky130_fd_sc_hd__clkbuf_1 _3933_ (.A(_1874_),
    .X(_0502_));
 sky130_fd_sc_hd__nor2_2 _3934_ (.A(_1258_),
    .B(_1403_),
    .Y(_1875_));
 sky130_fd_sc_hd__mux2_1 _3935_ (.A0(\tms1x00.RAM[90][0] ),
    .A1(_1323_),
    .S(_1875_),
    .X(_1876_));
 sky130_fd_sc_hd__clkbuf_1 _3936_ (.A(_1876_),
    .X(_0503_));
 sky130_fd_sc_hd__mux2_1 _3937_ (.A0(\tms1x00.RAM[90][1] ),
    .A1(_1327_),
    .S(_1875_),
    .X(_1877_));
 sky130_fd_sc_hd__clkbuf_1 _3938_ (.A(_1877_),
    .X(_0504_));
 sky130_fd_sc_hd__mux2_1 _3939_ (.A0(\tms1x00.RAM[90][2] ),
    .A1(_1330_),
    .S(_1875_),
    .X(_1878_));
 sky130_fd_sc_hd__clkbuf_1 _3940_ (.A(_1878_),
    .X(_0505_));
 sky130_fd_sc_hd__mux2_1 _3941_ (.A0(\tms1x00.RAM[90][3] ),
    .A1(_1333_),
    .S(_1875_),
    .X(_1879_));
 sky130_fd_sc_hd__clkbuf_1 _3942_ (.A(_1879_),
    .X(_0506_));
 sky130_fd_sc_hd__nor2_2 _3943_ (.A(_1250_),
    .B(_1310_),
    .Y(_1880_));
 sky130_fd_sc_hd__mux2_1 _3944_ (.A0(\tms1x00.RAM[23][0] ),
    .A1(_1323_),
    .S(_1880_),
    .X(_1881_));
 sky130_fd_sc_hd__clkbuf_1 _3945_ (.A(_1881_),
    .X(_0507_));
 sky130_fd_sc_hd__mux2_1 _3946_ (.A0(\tms1x00.RAM[23][1] ),
    .A1(_1327_),
    .S(_1880_),
    .X(_1882_));
 sky130_fd_sc_hd__clkbuf_1 _3947_ (.A(_1882_),
    .X(_0508_));
 sky130_fd_sc_hd__mux2_1 _3948_ (.A0(\tms1x00.RAM[23][2] ),
    .A1(_1330_),
    .S(_1880_),
    .X(_1883_));
 sky130_fd_sc_hd__clkbuf_1 _3949_ (.A(_1883_),
    .X(_0509_));
 sky130_fd_sc_hd__mux2_1 _3950_ (.A0(\tms1x00.RAM[23][3] ),
    .A1(_1333_),
    .S(_1880_),
    .X(_1884_));
 sky130_fd_sc_hd__clkbuf_1 _3951_ (.A(_1884_),
    .X(_0510_));
 sky130_fd_sc_hd__mux2_1 _3952_ (.A0(\tms1x00.Y[0] ),
    .A1(_0717_),
    .S(_0726_),
    .X(_1885_));
 sky130_fd_sc_hd__clkbuf_1 _3953_ (.A(_1885_),
    .X(_0511_));
 sky130_fd_sc_hd__mux2_1 _3954_ (.A0(\tms1x00.Y[1] ),
    .A1(_0728_),
    .S(_0726_),
    .X(_1886_));
 sky130_fd_sc_hd__clkbuf_1 _3955_ (.A(_1886_),
    .X(_0512_));
 sky130_fd_sc_hd__mux2_1 _3956_ (.A0(_0730_),
    .A1(\tms1x00.ram_addr_buff[2] ),
    .S(_0726_),
    .X(_1887_));
 sky130_fd_sc_hd__clkbuf_1 _3957_ (.A(_1887_),
    .X(_0513_));
 sky130_fd_sc_hd__mux2_1 _3958_ (.A0(_0733_),
    .A1(\tms1x00.ram_addr_buff[3] ),
    .S(_0725_),
    .X(_1888_));
 sky130_fd_sc_hd__clkbuf_1 _3959_ (.A(_1888_),
    .X(_0514_));
 sky130_fd_sc_hd__mux2_1 _3960_ (.A0(\tms1x00.X[2] ),
    .A1(\tms1x00.ram_addr_buff[4] ),
    .S(_0725_),
    .X(_1889_));
 sky130_fd_sc_hd__clkbuf_1 _3961_ (.A(_1889_),
    .X(_0515_));
 sky130_fd_sc_hd__mux2_1 _3962_ (.A0(\tms1x00.X[0] ),
    .A1(\tms1x00.ram_addr_buff[5] ),
    .S(_0725_),
    .X(_1890_));
 sky130_fd_sc_hd__clkbuf_1 _3963_ (.A(_1890_),
    .X(_0516_));
 sky130_fd_sc_hd__mux2_1 _3964_ (.A0(\tms1x00.X[1] ),
    .A1(\tms1x00.ram_addr_buff[6] ),
    .S(_0725_),
    .X(_1891_));
 sky130_fd_sc_hd__clkbuf_1 _3965_ (.A(_1891_),
    .X(_0517_));
 sky130_fd_sc_hd__and2_1 _3966_ (.A(\tms1x00.wb_step ),
    .B(_0766_),
    .X(_1892_));
 sky130_fd_sc_hd__clkbuf_1 _3967_ (.A(_1892_),
    .X(_0518_));
 sky130_fd_sc_hd__mux2_1 _3968_ (.A0(net1),
    .A1(chip_sel_override),
    .S(net148),
    .X(_1893_));
 sky130_fd_sc_hd__mux2_1 _3969_ (.A0(net93),
    .A1(_1893_),
    .S(_0738_),
    .X(_1894_));
 sky130_fd_sc_hd__clkbuf_1 _3970_ (.A(_1894_),
    .X(_0519_));
 sky130_fd_sc_hd__mux2_1 _3971_ (.A0(_0742_),
    .A1(net6),
    .S(_0724_),
    .X(_1895_));
 sky130_fd_sc_hd__or2_1 _3972_ (.A(net103),
    .B(_1895_),
    .X(_1896_));
 sky130_fd_sc_hd__clkbuf_1 _3973_ (.A(_1896_),
    .X(_0520_));
 sky130_fd_sc_hd__mux2_1 _3974_ (.A0(\tms1x00.ins_in[1] ),
    .A1(net7),
    .S(_0724_),
    .X(_1897_));
 sky130_fd_sc_hd__or2_1 _3975_ (.A(net103),
    .B(_1897_),
    .X(_1898_));
 sky130_fd_sc_hd__clkbuf_1 _3976_ (.A(_1898_),
    .X(_0521_));
 sky130_fd_sc_hd__or3b_1 _3977_ (.A(_0701_),
    .B(_0760_),
    .C_N(_0720_),
    .X(_1899_));
 sky130_fd_sc_hd__or2_1 _3978_ (.A(net8),
    .B(_1899_),
    .X(_1900_));
 sky130_fd_sc_hd__buf_4 _3979_ (.A(_0718_),
    .X(_1901_));
 sky130_fd_sc_hd__o211a_1 _3980_ (.A1(\tms1x00.ins_in[2] ),
    .A2(_0724_),
    .B1(_1900_),
    .C1(_1901_),
    .X(_0522_));
 sky130_fd_sc_hd__or2_1 _3981_ (.A(net9),
    .B(_1899_),
    .X(_1902_));
 sky130_fd_sc_hd__o211a_1 _3982_ (.A1(_0743_),
    .A2(_0724_),
    .B1(_1902_),
    .C1(_1901_),
    .X(_0523_));
 sky130_fd_sc_hd__or2_1 _3983_ (.A(net10),
    .B(_1899_),
    .X(_1903_));
 sky130_fd_sc_hd__o211a_1 _3984_ (.A1(\tms1x00.ins_in[4] ),
    .A2(_0724_),
    .B1(_1903_),
    .C1(_1901_),
    .X(_0524_));
 sky130_fd_sc_hd__mux2_1 _3985_ (.A0(\tms1x00.ins_in[5] ),
    .A1(net11),
    .S(_0724_),
    .X(_1904_));
 sky130_fd_sc_hd__or2_1 _3986_ (.A(net103),
    .B(_1904_),
    .X(_1905_));
 sky130_fd_sc_hd__clkbuf_1 _3987_ (.A(_1905_),
    .X(_0525_));
 sky130_fd_sc_hd__or2_1 _3988_ (.A(net12),
    .B(_1899_),
    .X(_1906_));
 sky130_fd_sc_hd__o211a_1 _3989_ (.A1(_0748_),
    .A2(_0724_),
    .B1(_1906_),
    .C1(_1901_),
    .X(_0526_));
 sky130_fd_sc_hd__or2_1 _3990_ (.A(net13),
    .B(_1899_),
    .X(_1907_));
 sky130_fd_sc_hd__o211a_1 _3991_ (.A1(_0747_),
    .A2(_0724_),
    .B1(_1907_),
    .C1(_1901_),
    .X(_0527_));
 sky130_fd_sc_hd__buf_2 _3992_ (.A(_0722_),
    .X(_1908_));
 sky130_fd_sc_hd__nand2_1 _3993_ (.A(_0701_),
    .B(_1908_),
    .Y(_1909_));
 sky130_fd_sc_hd__or2_1 _3994_ (.A(_0701_),
    .B(_1908_),
    .X(_1910_));
 sky130_fd_sc_hd__and3_1 _3995_ (.A(_0718_),
    .B(_1909_),
    .C(_1910_),
    .X(_1911_));
 sky130_fd_sc_hd__clkbuf_1 _3996_ (.A(_1911_),
    .X(_0528_));
 sky130_fd_sc_hd__nor2_1 _3997_ (.A(net76),
    .B(net75),
    .Y(_1912_));
 sky130_fd_sc_hd__a21o_1 _3998_ (.A1(_0701_),
    .A2(_1908_),
    .B1(net75),
    .X(_1913_));
 sky130_fd_sc_hd__o211a_1 _3999_ (.A1(_1909_),
    .A2(_1912_),
    .B1(_1913_),
    .C1(_1901_),
    .X(_0529_));
 sky130_fd_sc_hd__a21oi_1 _4000_ (.A1(net76),
    .A2(_1909_),
    .B1(_0761_),
    .Y(_1914_));
 sky130_fd_sc_hd__nor2_1 _4001_ (.A(net103),
    .B(_1914_),
    .Y(_0530_));
 sky130_fd_sc_hd__and2b_1 _4002_ (.A_N(\tms1x00.Y[1] ),
    .B(\tms1x00.Y[0] ),
    .X(_1915_));
 sky130_fd_sc_hd__and4_1 _4003_ (.A(_0755_),
    .B(_0739_),
    .C(_0764_),
    .D(_1915_),
    .X(_1916_));
 sky130_fd_sc_hd__or4b_1 _4004_ (.A(_0732_),
    .B(_0730_),
    .C(_0752_),
    .D_N(_1915_),
    .X(_1917_));
 sky130_fd_sc_hd__o211a_1 _4005_ (.A1(net78),
    .A2(_1916_),
    .B1(_1917_),
    .C1(_1901_),
    .X(_0531_));
 sky130_fd_sc_hd__and2b_1 _4006_ (.A_N(\tms1x00.Y[0] ),
    .B(\tms1x00.Y[1] ),
    .X(_1918_));
 sky130_fd_sc_hd__and4_1 _4007_ (.A(_0755_),
    .B(_0739_),
    .C(_0763_),
    .D(_1918_),
    .X(_1919_));
 sky130_fd_sc_hd__or4b_1 _4008_ (.A(_0732_),
    .B(_0730_),
    .C(_0752_),
    .D_N(_1918_),
    .X(_1920_));
 sky130_fd_sc_hd__o211a_1 _4009_ (.A1(net79),
    .A2(_1919_),
    .B1(_1920_),
    .C1(_1901_),
    .X(_0532_));
 sky130_fd_sc_hd__nand2_1 _4010_ (.A(\tms1x00.Y[1] ),
    .B(\tms1x00.Y[0] ),
    .Y(_1921_));
 sky130_fd_sc_hd__nor2_1 _4011_ (.A(\tms1x00.Y[2] ),
    .B(_1921_),
    .Y(_1922_));
 sky130_fd_sc_hd__nand3_1 _4012_ (.A(_0754_),
    .B(_0763_),
    .C(_1922_),
    .Y(_1923_));
 sky130_fd_sc_hd__inv_2 _4013_ (.A(_1923_),
    .Y(_1924_));
 sky130_fd_sc_hd__or3b_1 _4014_ (.A(_0732_),
    .B(_0753_),
    .C_N(_1922_),
    .X(_1925_));
 sky130_fd_sc_hd__o211a_1 _4015_ (.A1(net80),
    .A2(_1924_),
    .B1(_1925_),
    .C1(_1901_),
    .X(_0533_));
 sky130_fd_sc_hd__or3b_1 _4016_ (.A(_0732_),
    .B(_0739_),
    .C_N(_0740_),
    .X(_1926_));
 sky130_fd_sc_hd__a41o_1 _4017_ (.A1(_0755_),
    .A2(_0730_),
    .A3(_0740_),
    .A4(_0764_),
    .B1(net81),
    .X(_1927_));
 sky130_fd_sc_hd__o211a_1 _4018_ (.A1(_0753_),
    .A2(_1926_),
    .B1(_1927_),
    .C1(_1901_),
    .X(_0534_));
 sky130_fd_sc_hd__nand2_1 _4019_ (.A(\tms1x00.Y[2] ),
    .B(_1915_),
    .Y(_1928_));
 sky130_fd_sc_hd__and3b_1 _4020_ (.A_N(_1928_),
    .B(_0755_),
    .C(_0764_),
    .X(_1929_));
 sky130_fd_sc_hd__or3_1 _4021_ (.A(_0732_),
    .B(_0753_),
    .C(_1928_),
    .X(_1930_));
 sky130_fd_sc_hd__clkbuf_4 _4022_ (.A(_0718_),
    .X(_1931_));
 sky130_fd_sc_hd__o211a_1 _4023_ (.A1(net82),
    .A2(_1929_),
    .B1(_1930_),
    .C1(_1931_),
    .X(_0535_));
 sky130_fd_sc_hd__nand2_1 _4024_ (.A(\tms1x00.Y[2] ),
    .B(_1918_),
    .Y(_1932_));
 sky130_fd_sc_hd__and3b_1 _4025_ (.A_N(_1932_),
    .B(_0755_),
    .C(_0764_),
    .X(_1933_));
 sky130_fd_sc_hd__or3_1 _4026_ (.A(_0732_),
    .B(_0753_),
    .C(_1932_),
    .X(_1934_));
 sky130_fd_sc_hd__o211a_1 _4027_ (.A1(net83),
    .A2(_1933_),
    .B1(_1934_),
    .C1(_1931_),
    .X(_0536_));
 sky130_fd_sc_hd__nor2_1 _4028_ (.A(_0739_),
    .B(_1921_),
    .Y(_1935_));
 sky130_fd_sc_hd__a31o_1 _4029_ (.A1(_0754_),
    .A2(_0763_),
    .A3(_1935_),
    .B1(net84),
    .X(_1936_));
 sky130_fd_sc_hd__or3b_1 _4030_ (.A(\tms1x00.Y[3] ),
    .B(_0752_),
    .C_N(_1935_),
    .X(_1937_));
 sky130_fd_sc_hd__and3_1 _4031_ (.A(_0718_),
    .B(_1936_),
    .C(_1937_),
    .X(_1938_));
 sky130_fd_sc_hd__clkbuf_1 _4032_ (.A(_1938_),
    .X(_0537_));
 sky130_fd_sc_hd__a31o_1 _4033_ (.A1(_0733_),
    .A2(_0756_),
    .A3(_0764_),
    .B1(net85),
    .X(_1939_));
 sky130_fd_sc_hd__o311a_1 _4034_ (.A1(_0755_),
    .A2(_0741_),
    .A3(_0753_),
    .B1(_1939_),
    .C1(_0766_),
    .X(_0538_));
 sky130_fd_sc_hd__or3b_1 _4035_ (.A(_0755_),
    .B(_0730_),
    .C_N(_1915_),
    .X(_1940_));
 sky130_fd_sc_hd__a41o_1 _4036_ (.A1(_0733_),
    .A2(_0739_),
    .A3(_0764_),
    .A4(_1915_),
    .B1(net86),
    .X(_1941_));
 sky130_fd_sc_hd__o211a_1 _4037_ (.A1(_0753_),
    .A2(_1940_),
    .B1(_1941_),
    .C1(_1931_),
    .X(_0539_));
 sky130_fd_sc_hd__or3b_1 _4038_ (.A(_0754_),
    .B(_0730_),
    .C_N(_1918_),
    .X(_1942_));
 sky130_fd_sc_hd__a41o_1 _4039_ (.A1(_0733_),
    .A2(_0739_),
    .A3(_0764_),
    .A4(_1918_),
    .B1(net87),
    .X(_1943_));
 sky130_fd_sc_hd__o211a_1 _4040_ (.A1(_0753_),
    .A2(_1942_),
    .B1(_1943_),
    .C1(_1931_),
    .X(_0540_));
 sky130_fd_sc_hd__a31o_1 _4041_ (.A1(_0732_),
    .A2(_0763_),
    .A3(_1922_),
    .B1(net88),
    .X(_1944_));
 sky130_fd_sc_hd__or3b_1 _4042_ (.A(_0754_),
    .B(_0752_),
    .C_N(_1922_),
    .X(_1945_));
 sky130_fd_sc_hd__and3_1 _4043_ (.A(_0718_),
    .B(_1944_),
    .C(_1945_),
    .X(_1946_));
 sky130_fd_sc_hd__clkbuf_1 _4044_ (.A(_1946_),
    .X(_0541_));
 sky130_fd_sc_hd__and3_1 _4045_ (.A(\tms1x00.Y[3] ),
    .B(\tms1x00.Y[2] ),
    .C(_0740_),
    .X(_1947_));
 sky130_fd_sc_hd__inv_2 _4046_ (.A(_1947_),
    .Y(_1948_));
 sky130_fd_sc_hd__a21o_1 _4047_ (.A1(_0764_),
    .A2(_1947_),
    .B1(net89),
    .X(_1949_));
 sky130_fd_sc_hd__o211a_1 _4048_ (.A1(_0753_),
    .A2(_1948_),
    .B1(_1949_),
    .C1(_1931_),
    .X(_0542_));
 sky130_fd_sc_hd__and4_1 _4049_ (.A(_0733_),
    .B(_0730_),
    .C(_0763_),
    .D(_1915_),
    .X(_1950_));
 sky130_fd_sc_hd__or3_1 _4050_ (.A(_0755_),
    .B(_0752_),
    .C(_1928_),
    .X(_1951_));
 sky130_fd_sc_hd__o211a_1 _4051_ (.A1(net90),
    .A2(_1950_),
    .B1(_1951_),
    .C1(_1931_),
    .X(_0543_));
 sky130_fd_sc_hd__and4_1 _4052_ (.A(_0733_),
    .B(_0730_),
    .C(_0763_),
    .D(_1918_),
    .X(_1952_));
 sky130_fd_sc_hd__or3_1 _4053_ (.A(_0755_),
    .B(_0752_),
    .C(_1932_),
    .X(_1953_));
 sky130_fd_sc_hd__o211a_1 _4054_ (.A1(net91),
    .A2(_1952_),
    .B1(_1953_),
    .C1(_1931_),
    .X(_0544_));
 sky130_fd_sc_hd__nand2_1 _4055_ (.A(_0733_),
    .B(_1935_),
    .Y(_1954_));
 sky130_fd_sc_hd__a31o_1 _4056_ (.A1(_0733_),
    .A2(_0764_),
    .A3(_1935_),
    .B1(net92),
    .X(_1955_));
 sky130_fd_sc_hd__o211a_1 _4057_ (.A1(_0753_),
    .A2(_1954_),
    .B1(_1955_),
    .C1(_1931_),
    .X(_0545_));
 sky130_fd_sc_hd__nor2_2 _4058_ (.A(\tms1x00.ins_in[4] ),
    .B(_0749_),
    .Y(_1956_));
 sky130_fd_sc_hd__and4_1 _4059_ (.A(_0743_),
    .B(_0768_),
    .C(\tms1x00.ins_in[1] ),
    .D(_1956_),
    .X(_1957_));
 sky130_fd_sc_hd__nand2_1 _4060_ (.A(_0761_),
    .B(_1957_),
    .Y(_1958_));
 sky130_fd_sc_hd__and2b_1 _4061_ (.A_N(_0742_),
    .B(\tms1x00.A[0] ),
    .X(_1959_));
 sky130_fd_sc_hd__and2_1 _4062_ (.A(_0761_),
    .B(_1957_),
    .X(_1960_));
 sky130_fd_sc_hd__or2_1 _4063_ (.A(net69),
    .B(_1960_),
    .X(_1961_));
 sky130_fd_sc_hd__o211a_1 _4064_ (.A1(_1958_),
    .A2(_1959_),
    .B1(_1961_),
    .C1(_1931_),
    .X(_0546_));
 sky130_fd_sc_hd__and2b_1 _4065_ (.A_N(_0742_),
    .B(\tms1x00.A[1] ),
    .X(_1962_));
 sky130_fd_sc_hd__or2_1 _4066_ (.A(net70),
    .B(_1960_),
    .X(_1963_));
 sky130_fd_sc_hd__o211a_1 _4067_ (.A1(_1958_),
    .A2(_1962_),
    .B1(_1963_),
    .C1(_1931_),
    .X(_0547_));
 sky130_fd_sc_hd__and2b_1 _4068_ (.A_N(_0742_),
    .B(\tms1x00.A[2] ),
    .X(_1964_));
 sky130_fd_sc_hd__or2_1 _4069_ (.A(net71),
    .B(_1960_),
    .X(_1965_));
 sky130_fd_sc_hd__clkbuf_4 _4070_ (.A(_0718_),
    .X(_1966_));
 sky130_fd_sc_hd__o211a_1 _4071_ (.A1(_1958_),
    .A2(_1964_),
    .B1(_1965_),
    .C1(_1966_),
    .X(_0548_));
 sky130_fd_sc_hd__and2b_1 _4072_ (.A_N(_0742_),
    .B(\tms1x00.A[3] ),
    .X(_1967_));
 sky130_fd_sc_hd__or2_1 _4073_ (.A(net72),
    .B(_1960_),
    .X(_1968_));
 sky130_fd_sc_hd__o211a_1 _4074_ (.A1(_1958_),
    .A2(_1967_),
    .B1(_1968_),
    .C1(_1966_),
    .X(_0549_));
 sky130_fd_sc_hd__and2b_1 _4075_ (.A_N(_0742_),
    .B(\tms1x00.status ),
    .X(_1969_));
 sky130_fd_sc_hd__or2_1 _4076_ (.A(net73),
    .B(_1960_),
    .X(_1970_));
 sky130_fd_sc_hd__o211a_1 _4077_ (.A1(_1958_),
    .A2(_1969_),
    .B1(_1970_),
    .C1(_1966_),
    .X(_0550_));
 sky130_fd_sc_hd__nand2_4 _4078_ (.A(net74),
    .B(_0720_),
    .Y(_1971_));
 sky130_fd_sc_hd__nor2_1 _4079_ (.A(_0760_),
    .B(_1971_),
    .Y(_1972_));
 sky130_fd_sc_hd__and4_2 _4080_ (.A(\tms1x00.status ),
    .B(_0747_),
    .C(_0748_),
    .D(_1972_),
    .X(_1973_));
 sky130_fd_sc_hd__or2_1 _4081_ (.A(_0760_),
    .B(_1971_),
    .X(_1974_));
 sky130_fd_sc_hd__nand2_1 _4082_ (.A(\tms1x00.ins_in[1] ),
    .B(\tms1x00.ins_in[0] ),
    .Y(_1975_));
 sky130_fd_sc_hd__or4_1 _4083_ (.A(_0744_),
    .B(_0750_),
    .C(_1974_),
    .D(_1975_),
    .X(_1976_));
 sky130_fd_sc_hd__o211a_1 _4084_ (.A1(\tms1x00.CL ),
    .A2(_1973_),
    .B1(_1976_),
    .C1(_1966_),
    .X(_0551_));
 sky130_fd_sc_hd__or3_1 _4085_ (.A(\tms1x00.status ),
    .B(_0738_),
    .C(_1972_),
    .X(_1977_));
 sky130_fd_sc_hd__clkbuf_1 _4086_ (.A(_1977_),
    .X(_0552_));
 sky130_fd_sc_hd__nand2_1 _4087_ (.A(_0718_),
    .B(_1973_),
    .Y(_1978_));
 sky130_fd_sc_hd__nor2_4 _4088_ (.A(\tms1x00.CL ),
    .B(_1978_),
    .Y(_1979_));
 sky130_fd_sc_hd__mux2_1 _4089_ (.A0(\tms1x00.SR[0] ),
    .A1(\tms1x00.PC[0] ),
    .S(_1979_),
    .X(_1980_));
 sky130_fd_sc_hd__clkbuf_1 _4090_ (.A(_1980_),
    .X(_0553_));
 sky130_fd_sc_hd__mux2_1 _4091_ (.A0(\tms1x00.SR[1] ),
    .A1(\tms1x00.PC[1] ),
    .S(_1979_),
    .X(_1981_));
 sky130_fd_sc_hd__clkbuf_1 _4092_ (.A(_1981_),
    .X(_0554_));
 sky130_fd_sc_hd__mux2_1 _4093_ (.A0(\tms1x00.SR[2] ),
    .A1(\tms1x00.PC[2] ),
    .S(_1979_),
    .X(_1982_));
 sky130_fd_sc_hd__clkbuf_1 _4094_ (.A(_1982_),
    .X(_0555_));
 sky130_fd_sc_hd__mux2_1 _4095_ (.A0(\tms1x00.SR[3] ),
    .A1(\tms1x00.PC[3] ),
    .S(_1979_),
    .X(_1983_));
 sky130_fd_sc_hd__clkbuf_1 _4096_ (.A(_1983_),
    .X(_0556_));
 sky130_fd_sc_hd__mux2_1 _4097_ (.A0(\tms1x00.SR[4] ),
    .A1(\tms1x00.PC[4] ),
    .S(_1979_),
    .X(_1984_));
 sky130_fd_sc_hd__clkbuf_1 _4098_ (.A(_1984_),
    .X(_0557_));
 sky130_fd_sc_hd__mux2_1 _4099_ (.A0(\tms1x00.SR[5] ),
    .A1(\tms1x00.PC[5] ),
    .S(_1979_),
    .X(_1985_));
 sky130_fd_sc_hd__clkbuf_1 _4100_ (.A(_1985_),
    .X(_0558_));
 sky130_fd_sc_hd__nor2_1 _4101_ (.A(_0762_),
    .B(_0745_),
    .Y(_1986_));
 sky130_fd_sc_hd__a31oi_4 _4102_ (.A1(_0722_),
    .A2(_0758_),
    .A3(_1986_),
    .B1(_1973_),
    .Y(_1987_));
 sky130_fd_sc_hd__or3b_1 _4103_ (.A(\tms1x00.PB[0] ),
    .B(_0738_),
    .C_N(_1987_),
    .X(_1988_));
 sky130_fd_sc_hd__o21a_1 _4104_ (.A1(\tms1x00.PA[0] ),
    .A2(_1978_),
    .B1(_1988_),
    .X(_0559_));
 sky130_fd_sc_hd__a22o_1 _4105_ (.A1(\tms1x00.PA[1] ),
    .A2(_1973_),
    .B1(_1987_),
    .B2(\tms1x00.PB[1] ),
    .X(_1989_));
 sky130_fd_sc_hd__or2_1 _4106_ (.A(net103),
    .B(_1989_),
    .X(_1990_));
 sky130_fd_sc_hd__clkbuf_1 _4107_ (.A(_1990_),
    .X(_0560_));
 sky130_fd_sc_hd__a22o_1 _4108_ (.A1(\tms1x00.PA[2] ),
    .A2(_1973_),
    .B1(_1987_),
    .B2(\tms1x00.PB[2] ),
    .X(_1991_));
 sky130_fd_sc_hd__or2_1 _4109_ (.A(net103),
    .B(_1991_),
    .X(_1992_));
 sky130_fd_sc_hd__clkbuf_1 _4110_ (.A(_1992_),
    .X(_0561_));
 sky130_fd_sc_hd__a22o_1 _4111_ (.A1(\tms1x00.PA[3] ),
    .A2(_1973_),
    .B1(_1987_),
    .B2(\tms1x00.PB[3] ),
    .X(_1993_));
 sky130_fd_sc_hd__or2_1 _4112_ (.A(net103),
    .B(_1993_),
    .X(_1994_));
 sky130_fd_sc_hd__clkbuf_1 _4113_ (.A(_1994_),
    .X(_0562_));
 sky130_fd_sc_hd__nand2_4 _4114_ (.A(\tms1x00.status ),
    .B(_0747_),
    .Y(_1995_));
 sky130_fd_sc_hd__o31a_2 _4115_ (.A1(\tms1x00.CL ),
    .A2(_1974_),
    .A3(_1995_),
    .B1(_1976_),
    .X(_1996_));
 sky130_fd_sc_hd__mux2_1 _4116_ (.A0(\tms1x00.PB[0] ),
    .A1(\tms1x00.PA[0] ),
    .S(_1996_),
    .X(_1997_));
 sky130_fd_sc_hd__or2_1 _4117_ (.A(net103),
    .B(_1997_),
    .X(_1998_));
 sky130_fd_sc_hd__clkbuf_1 _4118_ (.A(_1998_),
    .X(_0563_));
 sky130_fd_sc_hd__mux2_1 _4119_ (.A0(\tms1x00.PB[1] ),
    .A1(\tms1x00.PA[1] ),
    .S(_1996_),
    .X(_1999_));
 sky130_fd_sc_hd__or2_1 _4120_ (.A(net103),
    .B(_1999_),
    .X(_2000_));
 sky130_fd_sc_hd__clkbuf_1 _4121_ (.A(_2000_),
    .X(_0564_));
 sky130_fd_sc_hd__mux2_1 _4122_ (.A0(\tms1x00.PB[2] ),
    .A1(\tms1x00.PA[2] ),
    .S(_1996_),
    .X(_2001_));
 sky130_fd_sc_hd__or2_1 _4123_ (.A(_0738_),
    .B(_2001_),
    .X(_2002_));
 sky130_fd_sc_hd__clkbuf_1 _4124_ (.A(_2002_),
    .X(_0565_));
 sky130_fd_sc_hd__mux2_1 _4125_ (.A0(\tms1x00.PB[3] ),
    .A1(\tms1x00.PA[3] ),
    .S(_1996_),
    .X(_2003_));
 sky130_fd_sc_hd__or2_1 _4126_ (.A(_0738_),
    .B(_2003_),
    .X(_2004_));
 sky130_fd_sc_hd__clkbuf_1 _4127_ (.A(_2004_),
    .X(_0566_));
 sky130_fd_sc_hd__or3b_1 _4128_ (.A(_0738_),
    .B(_0760_),
    .C_N(_1912_),
    .X(_2005_));
 sky130_fd_sc_hd__buf_4 _4129_ (.A(_2005_),
    .X(_2006_));
 sky130_fd_sc_hd__nor2_2 _4130_ (.A(_0701_),
    .B(_2006_),
    .Y(_2007_));
 sky130_fd_sc_hd__nand2_1 _4131_ (.A(_0858_),
    .B(_0903_),
    .Y(_2008_));
 sky130_fd_sc_hd__and4_1 _4132_ (.A(_0743_),
    .B(_0768_),
    .C(_0769_),
    .D(_0908_),
    .X(_2009_));
 sky130_fd_sc_hd__nor2_1 _4133_ (.A(_2008_),
    .B(_2009_),
    .Y(_2010_));
 sky130_fd_sc_hd__or2_1 _4134_ (.A(_0701_),
    .B(_2006_),
    .X(_2011_));
 sky130_fd_sc_hd__or2_1 _4135_ (.A(_0770_),
    .B(_1975_),
    .X(_2012_));
 sky130_fd_sc_hd__a32o_1 _4136_ (.A1(_0743_),
    .A2(\tms1x00.K_latch[0] ),
    .A3(_1956_),
    .B1(_2012_),
    .B2(\tms1x00.Y[0] ),
    .X(_2013_));
 sky130_fd_sc_hd__a211o_1 _4137_ (.A1(\tms1x00.ins_in[4] ),
    .A2(_1031_),
    .B1(_2011_),
    .C1(_2013_),
    .X(_2014_));
 sky130_fd_sc_hd__o22a_1 _4138_ (.A1(\tms1x00.P[0] ),
    .A2(_2007_),
    .B1(_2010_),
    .B2(_2014_),
    .X(_0567_));
 sky130_fd_sc_hd__and2b_1 _4139_ (.A_N(_2009_),
    .B(_1030_),
    .X(_2015_));
 sky130_fd_sc_hd__a32o_1 _4140_ (.A1(_0743_),
    .A2(\tms1x00.K_latch[1] ),
    .A3(_1956_),
    .B1(_2012_),
    .B2(\tms1x00.Y[1] ),
    .X(_2016_));
 sky130_fd_sc_hd__a211o_1 _4141_ (.A1(\tms1x00.ins_in[5] ),
    .A2(_1031_),
    .B1(_2011_),
    .C1(_2016_),
    .X(_2017_));
 sky130_fd_sc_hd__o22a_1 _4142_ (.A1(\tms1x00.P[1] ),
    .A2(_2007_),
    .B1(_2015_),
    .B2(_2017_),
    .X(_0568_));
 sky130_fd_sc_hd__and2b_1 _4143_ (.A_N(_2009_),
    .B(_1126_),
    .X(_2018_));
 sky130_fd_sc_hd__a31o_1 _4144_ (.A1(_0743_),
    .A2(\tms1x00.K_latch[2] ),
    .A3(_1956_),
    .B1(_1031_),
    .X(_2019_));
 sky130_fd_sc_hd__a211o_1 _4145_ (.A1(_0730_),
    .A2(_2012_),
    .B1(_2019_),
    .C1(_2011_),
    .X(_2020_));
 sky130_fd_sc_hd__o22a_1 _4146_ (.A1(\tms1x00.P[2] ),
    .A2(_2007_),
    .B1(_2018_),
    .B2(_2020_),
    .X(_0569_));
 sky130_fd_sc_hd__and2b_1 _4147_ (.A_N(_2009_),
    .B(_1221_),
    .X(_2021_));
 sky130_fd_sc_hd__a32o_1 _4148_ (.A1(_0743_),
    .A2(\tms1x00.K_latch[3] ),
    .A3(_1956_),
    .B1(_2012_),
    .B2(_0732_),
    .X(_2022_));
 sky130_fd_sc_hd__or2_1 _4149_ (.A(_2011_),
    .B(_2022_),
    .X(_2023_));
 sky130_fd_sc_hd__o22a_1 _4150_ (.A1(\tms1x00.P[3] ),
    .A2(_2007_),
    .B1(_2021_),
    .B2(_2023_),
    .X(_0570_));
 sky130_fd_sc_hd__and3b_1 _4151_ (.A_N(_0701_),
    .B(_0720_),
    .C(\tms1x00.PC[0] ),
    .X(_2024_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _4152_ (.A(_2024_),
    .X(_2025_));
 sky130_fd_sc_hd__inv_2 _4153_ (.A(\tms1x00.CL ),
    .Y(_2026_));
 sky130_fd_sc_hd__or4_4 _4154_ (.A(_2026_),
    .B(_0744_),
    .C(_0750_),
    .D(_1975_),
    .X(_2027_));
 sky130_fd_sc_hd__inv_2 _4155_ (.A(\tms1x00.SR[0] ),
    .Y(_2028_));
 sky130_fd_sc_hd__o221a_1 _4156_ (.A1(_0768_),
    .A2(_1995_),
    .B1(_2027_),
    .B2(_2028_),
    .C1(_0701_),
    .X(_2029_));
 sky130_fd_sc_hd__a21oi_4 _4157_ (.A1(_1995_),
    .A2(_2027_),
    .B1(_1971_),
    .Y(_2030_));
 sky130_fd_sc_hd__inv_2 _4158_ (.A(\tms1x00.PC[0] ),
    .Y(_2031_));
 sky130_fd_sc_hd__o32a_1 _4159_ (.A1(_0719_),
    .A2(net75),
    .A3(_2029_),
    .B1(_2030_),
    .B2(_2031_),
    .X(_2032_));
 sky130_fd_sc_hd__o21ai_1 _4160_ (.A1(_2025_),
    .A2(_2032_),
    .B1(_1908_),
    .Y(_2033_));
 sky130_fd_sc_hd__o211a_1 _4161_ (.A1(\tms1x00.PC[0] ),
    .A2(_1908_),
    .B1(_2033_),
    .C1(_1966_),
    .X(_0571_));
 sky130_fd_sc_hd__o22a_1 _4162_ (.A1(_0743_),
    .A2(_1995_),
    .B1(_2027_),
    .B2(\tms1x00.SR[1] ),
    .X(_2034_));
 sky130_fd_sc_hd__o22a_1 _4163_ (.A1(\tms1x00.PC[1] ),
    .A2(_2030_),
    .B1(_2034_),
    .B2(_1971_),
    .X(_2035_));
 sky130_fd_sc_hd__xor2_1 _4164_ (.A(_2025_),
    .B(_2035_),
    .X(_2036_));
 sky130_fd_sc_hd__or2_1 _4165_ (.A(\tms1x00.PC[1] ),
    .B(_1908_),
    .X(_2037_));
 sky130_fd_sc_hd__o211a_1 _4166_ (.A1(_0760_),
    .A2(_2036_),
    .B1(_2037_),
    .C1(_1966_),
    .X(_0572_));
 sky130_fd_sc_hd__nand2_1 _4167_ (.A(\tms1x00.PC[1] ),
    .B(_2025_),
    .Y(_2038_));
 sky130_fd_sc_hd__o22a_1 _4168_ (.A1(\tms1x00.ins_in[4] ),
    .A2(_1995_),
    .B1(_2027_),
    .B2(\tms1x00.SR[2] ),
    .X(_2039_));
 sky130_fd_sc_hd__o22a_1 _4169_ (.A1(\tms1x00.PC[2] ),
    .A2(_2030_),
    .B1(_2039_),
    .B2(_1971_),
    .X(_2040_));
 sky130_fd_sc_hd__nor2_1 _4170_ (.A(_2038_),
    .B(_2040_),
    .Y(_2041_));
 sky130_fd_sc_hd__a221o_1 _4171_ (.A1(net148),
    .A2(_0721_),
    .B1(_2038_),
    .B2(_2040_),
    .C1(_2041_),
    .X(_2042_));
 sky130_fd_sc_hd__o211a_1 _4172_ (.A1(\tms1x00.PC[2] ),
    .A2(_1908_),
    .B1(_2042_),
    .C1(_1966_),
    .X(_0573_));
 sky130_fd_sc_hd__and3_1 _4173_ (.A(\tms1x00.PC[2] ),
    .B(\tms1x00.PC[1] ),
    .C(_2025_),
    .X(_2043_));
 sky130_fd_sc_hd__o22a_1 _4174_ (.A1(\tms1x00.ins_in[5] ),
    .A2(_1995_),
    .B1(_2027_),
    .B2(\tms1x00.SR[3] ),
    .X(_2044_));
 sky130_fd_sc_hd__o22a_1 _4175_ (.A1(\tms1x00.PC[3] ),
    .A2(_2030_),
    .B1(_2044_),
    .B2(_1971_),
    .X(_2045_));
 sky130_fd_sc_hd__xor2_1 _4176_ (.A(_2043_),
    .B(_2045_),
    .X(_2046_));
 sky130_fd_sc_hd__or2_1 _4177_ (.A(\tms1x00.PC[3] ),
    .B(_1908_),
    .X(_2047_));
 sky130_fd_sc_hd__o211a_1 _4178_ (.A1(_0760_),
    .A2(_2046_),
    .B1(_2047_),
    .C1(_1966_),
    .X(_0574_));
 sky130_fd_sc_hd__and2_1 _4179_ (.A(\tms1x00.PC[3] ),
    .B(_2043_),
    .X(_2048_));
 sky130_fd_sc_hd__o22a_1 _4180_ (.A1(_0748_),
    .A2(_1995_),
    .B1(_2027_),
    .B2(\tms1x00.SR[4] ),
    .X(_2049_));
 sky130_fd_sc_hd__o22a_1 _4181_ (.A1(\tms1x00.PC[4] ),
    .A2(_2030_),
    .B1(_2049_),
    .B2(_1971_),
    .X(_2050_));
 sky130_fd_sc_hd__xor2_1 _4182_ (.A(_2048_),
    .B(_2050_),
    .X(_2051_));
 sky130_fd_sc_hd__or2_1 _4183_ (.A(\tms1x00.PC[4] ),
    .B(_1908_),
    .X(_2052_));
 sky130_fd_sc_hd__o211a_1 _4184_ (.A1(_0760_),
    .A2(_2051_),
    .B1(_2052_),
    .C1(_1966_),
    .X(_0575_));
 sky130_fd_sc_hd__or3_1 _4185_ (.A(\tms1x00.SR[5] ),
    .B(_1971_),
    .C(_2027_),
    .X(_2053_));
 sky130_fd_sc_hd__o21ai_1 _4186_ (.A1(\tms1x00.PC[5] ),
    .A2(_2030_),
    .B1(_2053_),
    .Y(_2054_));
 sky130_fd_sc_hd__a21oi_1 _4187_ (.A1(\tms1x00.PC[4] ),
    .A2(_2048_),
    .B1(_2054_),
    .Y(_2055_));
 sky130_fd_sc_hd__a31o_1 _4188_ (.A1(\tms1x00.PC[4] ),
    .A2(_2048_),
    .A3(_2054_),
    .B1(_0760_),
    .X(_2056_));
 sky130_fd_sc_hd__o21a_1 _4189_ (.A1(\tms1x00.PC[5] ),
    .A2(_1908_),
    .B1(_0766_),
    .X(_2057_));
 sky130_fd_sc_hd__o21a_1 _4190_ (.A1(_2055_),
    .A2(_2056_),
    .B1(_2057_),
    .X(_0576_));
 sky130_fd_sc_hd__or3b_2 _4191_ (.A(_0748_),
    .B(\tms1x00.ins_in[5] ),
    .C_N(_0747_),
    .X(_2058_));
 sky130_fd_sc_hd__or3_1 _4192_ (.A(\tms1x00.ins_in[4] ),
    .B(\tms1x00.N[0] ),
    .C(_2058_),
    .X(_2059_));
 sky130_fd_sc_hd__o21ai_1 _4193_ (.A1(\tms1x00.ins_in[4] ),
    .A2(_2058_),
    .B1(\tms1x00.N[0] ),
    .Y(_2060_));
 sky130_fd_sc_hd__and2_1 _4194_ (.A(_2059_),
    .B(_2060_),
    .X(_2061_));
 sky130_fd_sc_hd__xor2_1 _4195_ (.A(\tms1x00.P[0] ),
    .B(_2061_),
    .X(_2062_));
 sky130_fd_sc_hd__nor4b_4 _4196_ (.A(\tms1x00.ins_in[4] ),
    .B(_0746_),
    .C(_1127_),
    .D_N(\tms1x00.ins_in[5] ),
    .Y(_2063_));
 sky130_fd_sc_hd__mux2_1 _4197_ (.A0(\tms1x00.Y[0] ),
    .A1(_2062_),
    .S(_2063_),
    .X(_2064_));
 sky130_fd_sc_hd__and2_1 _4198_ (.A(_0766_),
    .B(_2064_),
    .X(_2065_));
 sky130_fd_sc_hd__clkbuf_1 _4199_ (.A(_2065_),
    .X(_0577_));
 sky130_fd_sc_hd__nand2_1 _4200_ (.A(\tms1x00.P[1] ),
    .B(\tms1x00.N[1] ),
    .Y(_2066_));
 sky130_fd_sc_hd__or2_1 _4201_ (.A(\tms1x00.P[1] ),
    .B(\tms1x00.N[1] ),
    .X(_2067_));
 sky130_fd_sc_hd__nand2_1 _4202_ (.A(_2066_),
    .B(_2067_),
    .Y(_2068_));
 sky130_fd_sc_hd__a21bo_1 _4203_ (.A1(\tms1x00.P[0] ),
    .A2(_2059_),
    .B1_N(_2060_),
    .X(_2069_));
 sky130_fd_sc_hd__xnor2_1 _4204_ (.A(_2068_),
    .B(_2069_),
    .Y(_2070_));
 sky130_fd_sc_hd__mux2_1 _4205_ (.A0(\tms1x00.Y[1] ),
    .A1(_2070_),
    .S(_2063_),
    .X(_2071_));
 sky130_fd_sc_hd__and2_1 _4206_ (.A(_0766_),
    .B(_2071_),
    .X(_2072_));
 sky130_fd_sc_hd__clkbuf_1 _4207_ (.A(_2072_),
    .X(_0578_));
 sky130_fd_sc_hd__and2_1 _4208_ (.A(\tms1x00.P[2] ),
    .B(\tms1x00.N[2] ),
    .X(_2073_));
 sky130_fd_sc_hd__nor2_1 _4209_ (.A(\tms1x00.P[2] ),
    .B(\tms1x00.N[2] ),
    .Y(_2074_));
 sky130_fd_sc_hd__nor2_1 _4210_ (.A(_2073_),
    .B(_2074_),
    .Y(_2075_));
 sky130_fd_sc_hd__a21boi_1 _4211_ (.A1(_2067_),
    .A2(_2069_),
    .B1_N(_2066_),
    .Y(_2076_));
 sky130_fd_sc_hd__xnor2_1 _4212_ (.A(_2075_),
    .B(_2076_),
    .Y(_2077_));
 sky130_fd_sc_hd__mux2_1 _4213_ (.A0(\tms1x00.Y[2] ),
    .A1(_2077_),
    .S(_2063_),
    .X(_2078_));
 sky130_fd_sc_hd__and2_1 _4214_ (.A(_0766_),
    .B(_2078_),
    .X(_2079_));
 sky130_fd_sc_hd__clkbuf_1 _4215_ (.A(_2079_),
    .X(_0579_));
 sky130_fd_sc_hd__o21ba_1 _4216_ (.A1(_2074_),
    .A2(_2076_),
    .B1_N(_2073_),
    .X(_2080_));
 sky130_fd_sc_hd__xor2_1 _4217_ (.A(\tms1x00.P[3] ),
    .B(\tms1x00.N[3] ),
    .X(_2081_));
 sky130_fd_sc_hd__xnor2_1 _4218_ (.A(_2080_),
    .B(_2081_),
    .Y(_2082_));
 sky130_fd_sc_hd__mux2_1 _4219_ (.A0(_0732_),
    .A1(_2082_),
    .S(_2063_),
    .X(_2083_));
 sky130_fd_sc_hd__and2_1 _4220_ (.A(_0766_),
    .B(_2083_),
    .X(_2084_));
 sky130_fd_sc_hd__clkbuf_1 _4221_ (.A(_2084_),
    .X(_0580_));
 sky130_fd_sc_hd__or4_1 _4222_ (.A(_0743_),
    .B(\tms1x00.ins_in[2] ),
    .C(\tms1x00.ins_in[1] ),
    .D(_0742_),
    .X(_2085_));
 sky130_fd_sc_hd__o22a_1 _4223_ (.A1(_0744_),
    .A2(_0904_),
    .B1(_2085_),
    .B2(_0750_),
    .X(_2086_));
 sky130_fd_sc_hd__nor2_1 _4224_ (.A(_0746_),
    .B(_2086_),
    .Y(_2087_));
 sky130_fd_sc_hd__and2b_1 _4225_ (.A_N(\tms1x00.ins_in[5] ),
    .B(_2087_),
    .X(_2088_));
 sky130_fd_sc_hd__nand2_1 _4226_ (.A(\tms1x00.X[0] ),
    .B(_2087_),
    .Y(_2089_));
 sky130_fd_sc_hd__o211a_1 _4227_ (.A1(\tms1x00.X[0] ),
    .A2(_2088_),
    .B1(_2089_),
    .C1(_1966_),
    .X(_0581_));
 sky130_fd_sc_hd__nand2_1 _4228_ (.A(\tms1x00.X[1] ),
    .B(_2087_),
    .Y(_2090_));
 sky130_fd_sc_hd__o211a_1 _4229_ (.A1(\tms1x00.X[1] ),
    .A2(_2088_),
    .B1(_2090_),
    .C1(_0766_),
    .X(_0582_));
 sky130_fd_sc_hd__nand2_1 _4230_ (.A(\tms1x00.X[2] ),
    .B(_2087_),
    .Y(_2091_));
 sky130_fd_sc_hd__o211a_1 _4231_ (.A1(\tms1x00.X[2] ),
    .A2(_2088_),
    .B1(_2091_),
    .C1(_0766_),
    .X(_0583_));
 sky130_fd_sc_hd__or2_1 _4232_ (.A(\tms1x00.N[0] ),
    .B(_2007_),
    .X(_2092_));
 sky130_fd_sc_hd__clkbuf_1 _4233_ (.A(_2092_),
    .X(_0584_));
 sky130_fd_sc_hd__or2_1 _4234_ (.A(\tms1x00.N[1] ),
    .B(_2007_),
    .X(_2093_));
 sky130_fd_sc_hd__clkbuf_1 _4235_ (.A(_2093_),
    .X(_0585_));
 sky130_fd_sc_hd__or2_1 _4236_ (.A(\tms1x00.N[2] ),
    .B(_2007_),
    .X(_2094_));
 sky130_fd_sc_hd__clkbuf_1 _4237_ (.A(_2094_),
    .X(_0586_));
 sky130_fd_sc_hd__or2_1 _4238_ (.A(\tms1x00.N[3] ),
    .B(_2007_),
    .X(_2095_));
 sky130_fd_sc_hd__clkbuf_1 _4239_ (.A(_2095_),
    .X(_0587_));
 sky130_fd_sc_hd__nor4_4 _4240_ (.A(_0762_),
    .B(_0738_),
    .C(_0746_),
    .D(_2058_),
    .Y(_2096_));
 sky130_fd_sc_hd__mux2_1 _4241_ (.A0(\tms1x00.A[0] ),
    .A1(_2062_),
    .S(_2096_),
    .X(_2097_));
 sky130_fd_sc_hd__clkbuf_1 _4242_ (.A(_2097_),
    .X(_0588_));
 sky130_fd_sc_hd__mux2_1 _4243_ (.A0(\tms1x00.A[1] ),
    .A1(_2070_),
    .S(_2096_),
    .X(_2098_));
 sky130_fd_sc_hd__clkbuf_1 _4244_ (.A(_2098_),
    .X(_0589_));
 sky130_fd_sc_hd__mux2_1 _4245_ (.A0(\tms1x00.A[2] ),
    .A1(_2077_),
    .S(_2096_),
    .X(_2099_));
 sky130_fd_sc_hd__clkbuf_1 _4246_ (.A(_2099_),
    .X(_0590_));
 sky130_fd_sc_hd__mux2_1 _4247_ (.A0(\tms1x00.A[3] ),
    .A1(_2082_),
    .S(_2096_),
    .X(_2100_));
 sky130_fd_sc_hd__clkbuf_1 _4248_ (.A(_2100_),
    .X(_0591_));
 sky130_fd_sc_hd__nor2_2 _4249_ (.A(_1310_),
    .B(_1430_),
    .Y(_2101_));
 sky130_fd_sc_hd__mux2_1 _4250_ (.A0(\tms1x00.RAM[119][0] ),
    .A1(_1323_),
    .S(_2101_),
    .X(_2102_));
 sky130_fd_sc_hd__clkbuf_1 _4251_ (.A(_2102_),
    .X(_0592_));
 sky130_fd_sc_hd__mux2_1 _4252_ (.A0(\tms1x00.RAM[119][1] ),
    .A1(_1327_),
    .S(_2101_),
    .X(_2103_));
 sky130_fd_sc_hd__clkbuf_1 _4253_ (.A(_2103_),
    .X(_0593_));
 sky130_fd_sc_hd__mux2_1 _4254_ (.A0(\tms1x00.RAM[119][2] ),
    .A1(_1330_),
    .S(_2101_),
    .X(_2104_));
 sky130_fd_sc_hd__clkbuf_1 _4255_ (.A(_2104_),
    .X(_0594_));
 sky130_fd_sc_hd__mux2_1 _4256_ (.A0(\tms1x00.RAM[119][3] ),
    .A1(_1333_),
    .S(_2101_),
    .X(_2105_));
 sky130_fd_sc_hd__clkbuf_1 _4257_ (.A(_2105_),
    .X(_0595_));
 sky130_fd_sc_hd__nor2_2 _4258_ (.A(_1310_),
    .B(_1525_),
    .Y(_2106_));
 sky130_fd_sc_hd__mux2_1 _4259_ (.A0(\tms1x00.RAM[39][0] ),
    .A1(_1323_),
    .S(_2106_),
    .X(_2107_));
 sky130_fd_sc_hd__clkbuf_1 _4260_ (.A(_2107_),
    .X(_0596_));
 sky130_fd_sc_hd__mux2_1 _4261_ (.A0(\tms1x00.RAM[39][1] ),
    .A1(_1327_),
    .S(_2106_),
    .X(_2108_));
 sky130_fd_sc_hd__clkbuf_1 _4262_ (.A(_2108_),
    .X(_0597_));
 sky130_fd_sc_hd__mux2_1 _4263_ (.A0(\tms1x00.RAM[39][2] ),
    .A1(_1330_),
    .S(_2106_),
    .X(_2109_));
 sky130_fd_sc_hd__clkbuf_1 _4264_ (.A(_2109_),
    .X(_0598_));
 sky130_fd_sc_hd__mux2_1 _4265_ (.A0(\tms1x00.RAM[39][3] ),
    .A1(_1333_),
    .S(_2106_),
    .X(_2110_));
 sky130_fd_sc_hd__clkbuf_1 _4266_ (.A(_2110_),
    .X(_0599_));
 sky130_fd_sc_hd__nor2_2 _4267_ (.A(_1250_),
    .B(_1317_),
    .Y(_2111_));
 sky130_fd_sc_hd__mux2_1 _4268_ (.A0(\tms1x00.RAM[22][0] ),
    .A1(_1323_),
    .S(_2111_),
    .X(_2112_));
 sky130_fd_sc_hd__clkbuf_1 _4269_ (.A(_2112_),
    .X(_0600_));
 sky130_fd_sc_hd__mux2_1 _4270_ (.A0(\tms1x00.RAM[22][1] ),
    .A1(_1327_),
    .S(_2111_),
    .X(_2113_));
 sky130_fd_sc_hd__clkbuf_1 _4271_ (.A(_2113_),
    .X(_0601_));
 sky130_fd_sc_hd__mux2_1 _4272_ (.A0(\tms1x00.RAM[22][2] ),
    .A1(_1330_),
    .S(_2111_),
    .X(_2114_));
 sky130_fd_sc_hd__clkbuf_1 _4273_ (.A(_2114_),
    .X(_0602_));
 sky130_fd_sc_hd__mux2_1 _4274_ (.A0(\tms1x00.RAM[22][3] ),
    .A1(_1333_),
    .S(_2111_),
    .X(_2115_));
 sky130_fd_sc_hd__clkbuf_1 _4275_ (.A(_2115_),
    .X(_0603_));
 sky130_fd_sc_hd__or2_2 _4276_ (.A(_0917_),
    .B(_1249_),
    .X(_2116_));
 sky130_fd_sc_hd__mux2_1 _4277_ (.A0(_1816_),
    .A1(\tms1x00.RAM[29][0] ),
    .S(_2116_),
    .X(_2117_));
 sky130_fd_sc_hd__clkbuf_1 _4278_ (.A(_2117_),
    .X(_0604_));
 sky130_fd_sc_hd__mux2_1 _4279_ (.A0(_1819_),
    .A1(\tms1x00.RAM[29][1] ),
    .S(_2116_),
    .X(_2118_));
 sky130_fd_sc_hd__clkbuf_1 _4280_ (.A(_2118_),
    .X(_0605_));
 sky130_fd_sc_hd__mux2_1 _4281_ (.A0(_1821_),
    .A1(\tms1x00.RAM[29][2] ),
    .S(_2116_),
    .X(_2119_));
 sky130_fd_sc_hd__clkbuf_1 _4282_ (.A(_2119_),
    .X(_0606_));
 sky130_fd_sc_hd__mux2_1 _4283_ (.A0(_1823_),
    .A1(\tms1x00.RAM[29][3] ),
    .S(_2116_),
    .X(_2120_));
 sky130_fd_sc_hd__clkbuf_1 _4284_ (.A(_2120_),
    .X(_0607_));
 sky130_fd_sc_hd__nor2_2 _4285_ (.A(_1240_),
    .B(_1250_),
    .Y(_2121_));
 sky130_fd_sc_hd__mux2_1 _4286_ (.A0(\tms1x00.RAM[21][0] ),
    .A1(_1323_),
    .S(_2121_),
    .X(_2122_));
 sky130_fd_sc_hd__clkbuf_1 _4287_ (.A(_2122_),
    .X(_0608_));
 sky130_fd_sc_hd__mux2_1 _4288_ (.A0(\tms1x00.RAM[21][1] ),
    .A1(_1327_),
    .S(_2121_),
    .X(_2123_));
 sky130_fd_sc_hd__clkbuf_1 _4289_ (.A(_2123_),
    .X(_0609_));
 sky130_fd_sc_hd__mux2_1 _4290_ (.A0(\tms1x00.RAM[21][2] ),
    .A1(_1330_),
    .S(_2121_),
    .X(_2124_));
 sky130_fd_sc_hd__clkbuf_1 _4291_ (.A(_2124_),
    .X(_0610_));
 sky130_fd_sc_hd__mux2_1 _4292_ (.A0(\tms1x00.RAM[21][3] ),
    .A1(_1333_),
    .S(_2121_),
    .X(_2125_));
 sky130_fd_sc_hd__clkbuf_1 _4293_ (.A(_2125_),
    .X(_0611_));
 sky130_fd_sc_hd__or2_2 _4294_ (.A(_1249_),
    .B(_1345_),
    .X(_2126_));
 sky130_fd_sc_hd__mux2_1 _4295_ (.A0(_1816_),
    .A1(\tms1x00.RAM[16][0] ),
    .S(_2126_),
    .X(_2127_));
 sky130_fd_sc_hd__clkbuf_1 _4296_ (.A(_2127_),
    .X(_0612_));
 sky130_fd_sc_hd__mux2_1 _4297_ (.A0(_1819_),
    .A1(\tms1x00.RAM[16][1] ),
    .S(_2126_),
    .X(_2128_));
 sky130_fd_sc_hd__clkbuf_1 _4298_ (.A(_2128_),
    .X(_0613_));
 sky130_fd_sc_hd__mux2_1 _4299_ (.A0(_1821_),
    .A1(\tms1x00.RAM[16][2] ),
    .S(_2126_),
    .X(_2129_));
 sky130_fd_sc_hd__clkbuf_1 _4300_ (.A(_2129_),
    .X(_0614_));
 sky130_fd_sc_hd__mux2_1 _4301_ (.A0(_1823_),
    .A1(\tms1x00.RAM[16][3] ),
    .S(_2126_),
    .X(_2130_));
 sky130_fd_sc_hd__clkbuf_1 _4302_ (.A(_2130_),
    .X(_0615_));
 sky130_fd_sc_hd__nor2_2 _4303_ (.A(_1250_),
    .B(_1337_),
    .Y(_2131_));
 sky130_fd_sc_hd__mux2_1 _4304_ (.A0(\tms1x00.RAM[20][0] ),
    .A1(_1323_),
    .S(_2131_),
    .X(_2132_));
 sky130_fd_sc_hd__clkbuf_1 _4305_ (.A(_2132_),
    .X(_0616_));
 sky130_fd_sc_hd__mux2_1 _4306_ (.A0(\tms1x00.RAM[20][1] ),
    .A1(_1327_),
    .S(_2131_),
    .X(_2133_));
 sky130_fd_sc_hd__clkbuf_1 _4307_ (.A(_2133_),
    .X(_0617_));
 sky130_fd_sc_hd__mux2_1 _4308_ (.A0(\tms1x00.RAM[20][2] ),
    .A1(_1330_),
    .S(_2131_),
    .X(_2134_));
 sky130_fd_sc_hd__clkbuf_1 _4309_ (.A(_2134_),
    .X(_0618_));
 sky130_fd_sc_hd__mux2_1 _4310_ (.A0(\tms1x00.RAM[20][3] ),
    .A1(_1333_),
    .S(_2131_),
    .X(_2135_));
 sky130_fd_sc_hd__clkbuf_1 _4311_ (.A(_2135_),
    .X(_0619_));
 sky130_fd_sc_hd__or2_2 _4312_ (.A(_1344_),
    .B(_1409_),
    .X(_2136_));
 sky130_fd_sc_hd__mux2_1 _4313_ (.A0(_1816_),
    .A1(\tms1x00.RAM[12][0] ),
    .S(_2136_),
    .X(_2137_));
 sky130_fd_sc_hd__clkbuf_1 _4314_ (.A(_2137_),
    .X(_0620_));
 sky130_fd_sc_hd__mux2_1 _4315_ (.A0(_1819_),
    .A1(\tms1x00.RAM[12][1] ),
    .S(_2136_),
    .X(_2138_));
 sky130_fd_sc_hd__clkbuf_1 _4316_ (.A(_2138_),
    .X(_0621_));
 sky130_fd_sc_hd__mux2_1 _4317_ (.A0(_1821_),
    .A1(\tms1x00.RAM[12][2] ),
    .S(_2136_),
    .X(_2139_));
 sky130_fd_sc_hd__clkbuf_1 _4318_ (.A(_2139_),
    .X(_0622_));
 sky130_fd_sc_hd__mux2_1 _4319_ (.A0(_1823_),
    .A1(\tms1x00.RAM[12][3] ),
    .S(_2136_),
    .X(_2140_));
 sky130_fd_sc_hd__clkbuf_1 _4320_ (.A(_2140_),
    .X(_0623_));
 sky130_fd_sc_hd__or2_2 _4321_ (.A(_1267_),
    .B(_1375_),
    .X(_2141_));
 sky130_fd_sc_hd__mux2_1 _4322_ (.A0(_1816_),
    .A1(\tms1x00.RAM[127][0] ),
    .S(_2141_),
    .X(_2142_));
 sky130_fd_sc_hd__clkbuf_1 _4323_ (.A(_2142_),
    .X(_0624_));
 sky130_fd_sc_hd__mux2_1 _4324_ (.A0(_1819_),
    .A1(\tms1x00.RAM[127][1] ),
    .S(_2141_),
    .X(_2143_));
 sky130_fd_sc_hd__clkbuf_1 _4325_ (.A(_2143_),
    .X(_0625_));
 sky130_fd_sc_hd__mux2_1 _4326_ (.A0(_1821_),
    .A1(\tms1x00.RAM[127][2] ),
    .S(_2141_),
    .X(_2144_));
 sky130_fd_sc_hd__clkbuf_1 _4327_ (.A(_2144_),
    .X(_0626_));
 sky130_fd_sc_hd__mux2_1 _4328_ (.A0(_1823_),
    .A1(\tms1x00.RAM[127][3] ),
    .S(_2141_),
    .X(_2145_));
 sky130_fd_sc_hd__clkbuf_1 _4329_ (.A(_2145_),
    .X(_0627_));
 sky130_fd_sc_hd__or2_2 _4330_ (.A(_1267_),
    .B(_1343_),
    .X(_2146_));
 sky130_fd_sc_hd__mux2_1 _4331_ (.A0(_1235_),
    .A1(\tms1x00.RAM[15][0] ),
    .S(_2146_),
    .X(_2147_));
 sky130_fd_sc_hd__clkbuf_1 _4332_ (.A(_2147_),
    .X(_0628_));
 sky130_fd_sc_hd__mux2_1 _4333_ (.A0(_1243_),
    .A1(\tms1x00.RAM[15][1] ),
    .S(_2146_),
    .X(_2148_));
 sky130_fd_sc_hd__clkbuf_1 _4334_ (.A(_2148_),
    .X(_0629_));
 sky130_fd_sc_hd__mux2_1 _4335_ (.A0(_1245_),
    .A1(\tms1x00.RAM[15][2] ),
    .S(_2146_),
    .X(_2149_));
 sky130_fd_sc_hd__clkbuf_1 _4336_ (.A(_2149_),
    .X(_0630_));
 sky130_fd_sc_hd__mux2_1 _4337_ (.A0(_1247_),
    .A1(\tms1x00.RAM[15][3] ),
    .S(_2146_),
    .X(_2150_));
 sky130_fd_sc_hd__clkbuf_1 _4338_ (.A(_2150_),
    .X(_0631_));
 sky130_fd_sc_hd__or2_2 _4339_ (.A(_1251_),
    .B(_1343_),
    .X(_2151_));
 sky130_fd_sc_hd__mux2_1 _4340_ (.A0(_1235_),
    .A1(\tms1x00.RAM[1][0] ),
    .S(_2151_),
    .X(_2152_));
 sky130_fd_sc_hd__clkbuf_1 _4341_ (.A(_2152_),
    .X(_0632_));
 sky130_fd_sc_hd__mux2_1 _4342_ (.A0(_1243_),
    .A1(\tms1x00.RAM[1][1] ),
    .S(_2151_),
    .X(_2153_));
 sky130_fd_sc_hd__clkbuf_1 _4343_ (.A(_2153_),
    .X(_0633_));
 sky130_fd_sc_hd__mux2_1 _4344_ (.A0(_1245_),
    .A1(\tms1x00.RAM[1][2] ),
    .S(_2151_),
    .X(_2154_));
 sky130_fd_sc_hd__clkbuf_1 _4345_ (.A(_2154_),
    .X(_0634_));
 sky130_fd_sc_hd__mux2_1 _4346_ (.A0(_1247_),
    .A1(\tms1x00.RAM[1][3] ),
    .S(_2151_),
    .X(_2155_));
 sky130_fd_sc_hd__clkbuf_1 _4347_ (.A(_2155_),
    .X(_0635_));
 sky130_fd_sc_hd__or2_2 _4348_ (.A(_0917_),
    .B(_1343_),
    .X(_2156_));
 sky130_fd_sc_hd__mux2_1 _4349_ (.A0(_1235_),
    .A1(\tms1x00.RAM[13][0] ),
    .S(_2156_),
    .X(_2157_));
 sky130_fd_sc_hd__clkbuf_1 _4350_ (.A(_2157_),
    .X(_0636_));
 sky130_fd_sc_hd__mux2_1 _4351_ (.A0(_1243_),
    .A1(\tms1x00.RAM[13][1] ),
    .S(_2156_),
    .X(_2158_));
 sky130_fd_sc_hd__clkbuf_1 _4352_ (.A(_2158_),
    .X(_0637_));
 sky130_fd_sc_hd__mux2_1 _4353_ (.A0(_1245_),
    .A1(\tms1x00.RAM[13][2] ),
    .S(_2156_),
    .X(_2159_));
 sky130_fd_sc_hd__clkbuf_1 _4354_ (.A(_2159_),
    .X(_0638_));
 sky130_fd_sc_hd__mux2_1 _4355_ (.A0(_1247_),
    .A1(\tms1x00.RAM[13][3] ),
    .S(_2156_),
    .X(_2160_));
 sky130_fd_sc_hd__clkbuf_1 _4356_ (.A(_2160_),
    .X(_0639_));
 sky130_fd_sc_hd__or2_2 _4357_ (.A(_1343_),
    .B(_1396_),
    .X(_2161_));
 sky130_fd_sc_hd__mux2_1 _4358_ (.A0(_1235_),
    .A1(\tms1x00.RAM[14][0] ),
    .S(_2161_),
    .X(_2162_));
 sky130_fd_sc_hd__clkbuf_1 _4359_ (.A(_2162_),
    .X(_0640_));
 sky130_fd_sc_hd__mux2_1 _4360_ (.A0(_1243_),
    .A1(\tms1x00.RAM[14][1] ),
    .S(_2161_),
    .X(_2163_));
 sky130_fd_sc_hd__clkbuf_1 _4361_ (.A(_2163_),
    .X(_0641_));
 sky130_fd_sc_hd__mux2_1 _4362_ (.A0(_1245_),
    .A1(\tms1x00.RAM[14][2] ),
    .S(_2161_),
    .X(_2164_));
 sky130_fd_sc_hd__clkbuf_1 _4363_ (.A(_2164_),
    .X(_0642_));
 sky130_fd_sc_hd__mux2_1 _4364_ (.A0(_1247_),
    .A1(\tms1x00.RAM[14][3] ),
    .S(_2161_),
    .X(_2165_));
 sky130_fd_sc_hd__clkbuf_1 _4365_ (.A(_2165_),
    .X(_0643_));
 sky130_fd_sc_hd__nor2_2 _4366_ (.A(_1261_),
    .B(_1344_),
    .Y(_2166_));
 sky130_fd_sc_hd__mux2_1 _4367_ (.A0(\tms1x00.RAM[9][0] ),
    .A1(_1323_),
    .S(_2166_),
    .X(_2167_));
 sky130_fd_sc_hd__clkbuf_1 _4368_ (.A(_2167_),
    .X(_0644_));
 sky130_fd_sc_hd__mux2_1 _4369_ (.A0(\tms1x00.RAM[9][1] ),
    .A1(_1327_),
    .S(_2166_),
    .X(_2168_));
 sky130_fd_sc_hd__clkbuf_1 _4370_ (.A(_2168_),
    .X(_0645_));
 sky130_fd_sc_hd__mux2_1 _4371_ (.A0(\tms1x00.RAM[9][2] ),
    .A1(_1330_),
    .S(_2166_),
    .X(_2169_));
 sky130_fd_sc_hd__clkbuf_1 _4372_ (.A(_2169_),
    .X(_0646_));
 sky130_fd_sc_hd__mux2_1 _4373_ (.A0(\tms1x00.RAM[9][3] ),
    .A1(_1333_),
    .S(_2166_),
    .X(_2170_));
 sky130_fd_sc_hd__clkbuf_1 _4374_ (.A(_2170_),
    .X(_0647_));
 sky130_fd_sc_hd__mux2_1 _4375_ (.A0(\tms1x00.PC[2] ),
    .A1(net95),
    .S(_2006_),
    .X(_2171_));
 sky130_fd_sc_hd__clkbuf_1 _4376_ (.A(_2171_),
    .X(_0648_));
 sky130_fd_sc_hd__mux2_1 _4377_ (.A0(\tms1x00.PC[3] ),
    .A1(net96),
    .S(_2006_),
    .X(_2172_));
 sky130_fd_sc_hd__clkbuf_1 _4378_ (.A(_2172_),
    .X(_0649_));
 sky130_fd_sc_hd__mux2_1 _4379_ (.A0(\tms1x00.PC[4] ),
    .A1(net97),
    .S(_2006_),
    .X(_2173_));
 sky130_fd_sc_hd__clkbuf_1 _4380_ (.A(_2173_),
    .X(_0650_));
 sky130_fd_sc_hd__mux2_1 _4381_ (.A0(\tms1x00.PC[5] ),
    .A1(net98),
    .S(_2006_),
    .X(_2174_));
 sky130_fd_sc_hd__clkbuf_1 _4382_ (.A(_2174_),
    .X(_0651_));
 sky130_fd_sc_hd__mux2_1 _4383_ (.A0(\tms1x00.PA[0] ),
    .A1(net99),
    .S(_2006_),
    .X(_2175_));
 sky130_fd_sc_hd__clkbuf_1 _4384_ (.A(_2175_),
    .X(_0652_));
 sky130_fd_sc_hd__mux2_1 _4385_ (.A0(\tms1x00.PA[1] ),
    .A1(net100),
    .S(_2006_),
    .X(_2176_));
 sky130_fd_sc_hd__clkbuf_1 _4386_ (.A(_2176_),
    .X(_0653_));
 sky130_fd_sc_hd__mux2_1 _4387_ (.A0(\tms1x00.PA[2] ),
    .A1(net101),
    .S(_2006_),
    .X(_2177_));
 sky130_fd_sc_hd__clkbuf_1 _4388_ (.A(_2177_),
    .X(_0654_));
 sky130_fd_sc_hd__mux2_1 _4389_ (.A0(\tms1x00.PA[3] ),
    .A1(net102),
    .S(_2006_),
    .X(_2178_));
 sky130_fd_sc_hd__clkbuf_1 _4390_ (.A(_2178_),
    .X(_0655_));
 sky130_fd_sc_hd__dfxtp_2 _4391_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0049_),
    .Q(net77));
 sky130_fd_sc_hd__dfxtp_4 _4392_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0000_),
    .Q(net94));
 sky130_fd_sc_hd__dfxtp_2 _4393_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0002_),
    .Q(\tms1x00.wb_step ));
 sky130_fd_sc_hd__dfxtp_1 _4394_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0001_),
    .Q(wb_rst_override));
 sky130_fd_sc_hd__dfxtp_1 _4395_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0050_),
    .Q(chip_sel_override));
 sky130_fd_sc_hd__dfxtp_1 _4396_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0003_),
    .Q(\wbs_o_buff[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4397_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0014_),
    .Q(\wbs_o_buff[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4398_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0025_),
    .Q(\wbs_o_buff[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4399_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0028_),
    .Q(\wbs_o_buff[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4400_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0029_),
    .Q(\wbs_o_buff[4] ));
 sky130_fd_sc_hd__dfxtp_1 _4401_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0030_),
    .Q(\wbs_o_buff[5] ));
 sky130_fd_sc_hd__dfxtp_1 _4402_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0031_),
    .Q(\wbs_o_buff[6] ));
 sky130_fd_sc_hd__dfxtp_1 _4403_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0032_),
    .Q(\wbs_o_buff[7] ));
 sky130_fd_sc_hd__dfxtp_1 _4404_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0033_),
    .Q(\wbs_o_buff[8] ));
 sky130_fd_sc_hd__dfxtp_1 _4405_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0034_),
    .Q(\wbs_o_buff[9] ));
 sky130_fd_sc_hd__dfxtp_1 _4406_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0004_),
    .Q(\wbs_o_buff[10] ));
 sky130_fd_sc_hd__dfxtp_1 _4407_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0005_),
    .Q(\wbs_o_buff[11] ));
 sky130_fd_sc_hd__dfxtp_1 _4408_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0006_),
    .Q(\wbs_o_buff[12] ));
 sky130_fd_sc_hd__dfxtp_1 _4409_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0007_),
    .Q(\wbs_o_buff[13] ));
 sky130_fd_sc_hd__dfxtp_1 _4410_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0008_),
    .Q(\wbs_o_buff[14] ));
 sky130_fd_sc_hd__dfxtp_1 _4411_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0009_),
    .Q(\wbs_o_buff[15] ));
 sky130_fd_sc_hd__dfxtp_1 _4412_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0010_),
    .Q(\wbs_o_buff[16] ));
 sky130_fd_sc_hd__dfxtp_1 _4413_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0011_),
    .Q(\wbs_o_buff[17] ));
 sky130_fd_sc_hd__dfxtp_1 _4414_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0012_),
    .Q(\wbs_o_buff[18] ));
 sky130_fd_sc_hd__dfxtp_1 _4415_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0013_),
    .Q(\wbs_o_buff[19] ));
 sky130_fd_sc_hd__dfxtp_1 _4416_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0015_),
    .Q(\wbs_o_buff[20] ));
 sky130_fd_sc_hd__dfxtp_1 _4417_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0016_),
    .Q(\wbs_o_buff[21] ));
 sky130_fd_sc_hd__dfxtp_1 _4418_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0017_),
    .Q(\wbs_o_buff[22] ));
 sky130_fd_sc_hd__dfxtp_1 _4419_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0018_),
    .Q(\wbs_o_buff[23] ));
 sky130_fd_sc_hd__dfxtp_1 _4420_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0019_),
    .Q(\wbs_o_buff[24] ));
 sky130_fd_sc_hd__dfxtp_1 _4421_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0020_),
    .Q(\wbs_o_buff[25] ));
 sky130_fd_sc_hd__dfxtp_1 _4422_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0021_),
    .Q(\wbs_o_buff[26] ));
 sky130_fd_sc_hd__dfxtp_1 _4423_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0022_),
    .Q(\wbs_o_buff[27] ));
 sky130_fd_sc_hd__dfxtp_1 _4424_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0023_),
    .Q(\wbs_o_buff[28] ));
 sky130_fd_sc_hd__dfxtp_1 _4425_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0024_),
    .Q(\wbs_o_buff[29] ));
 sky130_fd_sc_hd__dfxtp_1 _4426_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0026_),
    .Q(\wbs_o_buff[30] ));
 sky130_fd_sc_hd__dfxtp_1 _4427_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0027_),
    .Q(\wbs_o_buff[31] ));
 sky130_fd_sc_hd__dfxtp_1 _4428_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(net200),
    .Q(net115));
 sky130_fd_sc_hd__dfxtp_1 _4429_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(valid),
    .Q(feedback_delay));
 sky130_fd_sc_hd__dfxtp_1 _4430_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0051_),
    .Q(\tms1x00.RAM[109][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4431_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0052_),
    .Q(\tms1x00.RAM[109][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4432_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0053_),
    .Q(\tms1x00.RAM[109][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4433_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0054_),
    .Q(\tms1x00.RAM[109][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4434_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0055_),
    .Q(\tms1x00.RAM[99][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4435_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0056_),
    .Q(\tms1x00.RAM[99][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4436_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0057_),
    .Q(\tms1x00.RAM[99][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4437_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0058_),
    .Q(\tms1x00.RAM[99][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4438_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0059_),
    .Q(\tms1x00.RAM[69][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4439_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0060_),
    .Q(\tms1x00.RAM[69][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4440_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0061_),
    .Q(\tms1x00.RAM[69][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4441_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0062_),
    .Q(\tms1x00.RAM[69][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4442_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0063_),
    .Q(\tms1x00.RAM[17][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4443_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0064_),
    .Q(\tms1x00.RAM[17][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4444_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0065_),
    .Q(\tms1x00.RAM[17][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4445_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0066_),
    .Q(\tms1x00.RAM[17][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4446_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0067_),
    .Q(\tms1x00.RAM[89][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4447_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0068_),
    .Q(\tms1x00.RAM[89][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4448_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0069_),
    .Q(\tms1x00.RAM[89][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4449_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0070_),
    .Q(\tms1x00.RAM[89][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4450_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0071_),
    .Q(\tms1x00.RAM[79][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4451_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0072_),
    .Q(\tms1x00.RAM[79][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4452_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0073_),
    .Q(\tms1x00.RAM[79][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4453_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0074_),
    .Q(\tms1x00.RAM[79][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4454_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0075_),
    .Q(\tms1x00.RAM[18][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4455_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0076_),
    .Q(\tms1x00.RAM[18][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4456_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0077_),
    .Q(\tms1x00.RAM[18][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4457_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0078_),
    .Q(\tms1x00.RAM[18][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4458_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0079_),
    .Q(\K_override[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4459_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0080_),
    .Q(\K_override[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4460_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0081_),
    .Q(\K_override[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4461_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0082_),
    .Q(\K_override[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4462_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0083_),
    .Q(\tms1x00.RAM[59][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4463_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0084_),
    .Q(\tms1x00.RAM[59][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4464_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0085_),
    .Q(\tms1x00.RAM[59][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4465_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0086_),
    .Q(\tms1x00.RAM[59][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4466_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0087_),
    .Q(\tms1x00.RAM[49][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4467_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0088_),
    .Q(\tms1x00.RAM[49][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4468_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0089_),
    .Q(\tms1x00.RAM[49][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4469_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0090_),
    .Q(\tms1x00.RAM[49][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4470_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0091_),
    .Q(\tms1x00.RAM[19][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4471_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0092_),
    .Q(\tms1x00.RAM[19][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4472_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0093_),
    .Q(\tms1x00.RAM[19][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4473_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0094_),
    .Q(\tms1x00.RAM[19][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4474_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0095_),
    .Q(\tms1x00.RAM[104][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4475_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0096_),
    .Q(\tms1x00.RAM[104][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4476_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0097_),
    .Q(\tms1x00.RAM[104][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4477_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0098_),
    .Q(\tms1x00.RAM[104][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4478_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0099_),
    .Q(\tms1x00.RAM[103][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4479_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0100_),
    .Q(\tms1x00.RAM[103][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4480_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0101_),
    .Q(\tms1x00.RAM[103][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4481_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0102_),
    .Q(\tms1x00.RAM[103][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4482_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0103_),
    .Q(\tms1x00.RAM[102][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4483_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0104_),
    .Q(\tms1x00.RAM[102][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4484_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0105_),
    .Q(\tms1x00.RAM[102][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4485_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0106_),
    .Q(\tms1x00.RAM[102][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4486_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0107_),
    .Q(\tms1x00.RAM[101][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4487_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0108_),
    .Q(\tms1x00.RAM[101][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4488_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0109_),
    .Q(\tms1x00.RAM[101][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4489_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0110_),
    .Q(\tms1x00.RAM[101][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4490_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0111_),
    .Q(\tms1x00.RAM[100][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4491_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0112_),
    .Q(\tms1x00.RAM[100][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4492_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0113_),
    .Q(\tms1x00.RAM[100][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4493_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0114_),
    .Q(\tms1x00.RAM[100][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4494_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0115_),
    .Q(\tms1x00.RAM[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4495_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0116_),
    .Q(\tms1x00.RAM[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4496_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0117_),
    .Q(\tms1x00.RAM[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4497_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0118_),
    .Q(\tms1x00.RAM[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4498_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0119_),
    .Q(\tms1x00.RAM[98][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4499_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0120_),
    .Q(\tms1x00.RAM[98][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4500_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0121_),
    .Q(\tms1x00.RAM[98][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4501_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0122_),
    .Q(\tms1x00.RAM[98][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4502_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0123_),
    .Q(\tms1x00.RAM[97][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4503_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0124_),
    .Q(\tms1x00.RAM[97][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4504_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0125_),
    .Q(\tms1x00.RAM[97][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4505_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0126_),
    .Q(\tms1x00.RAM[97][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4506_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0127_),
    .Q(\tms1x00.RAM[96][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4507_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0128_),
    .Q(\tms1x00.RAM[96][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4508_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0129_),
    .Q(\tms1x00.RAM[96][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4509_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0130_),
    .Q(\tms1x00.RAM[96][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4510_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0131_),
    .Q(\tms1x00.RAM[95][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4511_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0132_),
    .Q(\tms1x00.RAM[95][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4512_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0133_),
    .Q(\tms1x00.RAM[95][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4513_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0134_),
    .Q(\tms1x00.RAM[95][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4514_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0135_),
    .Q(\tms1x00.RAM[114][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4515_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0136_),
    .Q(\tms1x00.RAM[114][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4516_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0137_),
    .Q(\tms1x00.RAM[114][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4517_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0138_),
    .Q(\tms1x00.RAM[114][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4518_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0139_),
    .Q(\tms1x00.RAM[113][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4519_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0140_),
    .Q(\tms1x00.RAM[113][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4520_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0141_),
    .Q(\tms1x00.RAM[113][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4521_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0142_),
    .Q(\tms1x00.RAM[113][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4522_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0143_),
    .Q(\tms1x00.RAM[112][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4523_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0144_),
    .Q(\tms1x00.RAM[112][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4524_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0145_),
    .Q(\tms1x00.RAM[112][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4525_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0146_),
    .Q(\tms1x00.RAM[112][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4526_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0147_),
    .Q(\tms1x00.RAM[111][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4527_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0148_),
    .Q(\tms1x00.RAM[111][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4528_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0149_),
    .Q(\tms1x00.RAM[111][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4529_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0150_),
    .Q(\tms1x00.RAM[111][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4530_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0151_),
    .Q(\tms1x00.RAM[110][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4531_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0152_),
    .Q(\tms1x00.RAM[110][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4532_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0153_),
    .Q(\tms1x00.RAM[110][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4533_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0154_),
    .Q(\tms1x00.RAM[110][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4534_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0155_),
    .Q(\tms1x00.RAM[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4535_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0156_),
    .Q(\tms1x00.RAM[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4536_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0157_),
    .Q(\tms1x00.RAM[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4537_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0158_),
    .Q(\tms1x00.RAM[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4538_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0159_),
    .Q(\tms1x00.RAM[108][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4539_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0160_),
    .Q(\tms1x00.RAM[108][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4540_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0161_),
    .Q(\tms1x00.RAM[108][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4541_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0162_),
    .Q(\tms1x00.RAM[108][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4542_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0163_),
    .Q(\tms1x00.RAM[107][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4543_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0164_),
    .Q(\tms1x00.RAM[107][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4544_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0165_),
    .Q(\tms1x00.RAM[107][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4545_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0166_),
    .Q(\tms1x00.RAM[107][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4546_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0167_),
    .Q(\tms1x00.RAM[106][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4547_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0168_),
    .Q(\tms1x00.RAM[106][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4548_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0169_),
    .Q(\tms1x00.RAM[106][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4549_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0170_),
    .Q(\tms1x00.RAM[106][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4550_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0171_),
    .Q(\tms1x00.RAM[105][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4551_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0172_),
    .Q(\tms1x00.RAM[105][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4552_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0173_),
    .Q(\tms1x00.RAM[105][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4553_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0174_),
    .Q(\tms1x00.RAM[105][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4554_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0175_),
    .Q(\tms1x00.RAM[124][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4555_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0176_),
    .Q(\tms1x00.RAM[124][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4556_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0177_),
    .Q(\tms1x00.RAM[124][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4557_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0178_),
    .Q(\tms1x00.RAM[124][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4558_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0179_),
    .Q(\tms1x00.RAM[123][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4559_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0180_),
    .Q(\tms1x00.RAM[123][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4560_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0181_),
    .Q(\tms1x00.RAM[123][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4561_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0182_),
    .Q(\tms1x00.RAM[123][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4562_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0183_),
    .Q(\tms1x00.RAM[122][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4563_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0184_),
    .Q(\tms1x00.RAM[122][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4564_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0185_),
    .Q(\tms1x00.RAM[122][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4565_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0186_),
    .Q(\tms1x00.RAM[122][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4566_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0187_),
    .Q(\tms1x00.RAM[121][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4567_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0188_),
    .Q(\tms1x00.RAM[121][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4568_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0189_),
    .Q(\tms1x00.RAM[121][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4569_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0190_),
    .Q(\tms1x00.RAM[121][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4570_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0191_),
    .Q(\tms1x00.RAM[120][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4571_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0192_),
    .Q(\tms1x00.RAM[120][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4572_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0193_),
    .Q(\tms1x00.RAM[120][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4573_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0194_),
    .Q(\tms1x00.RAM[120][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4574_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0195_),
    .Q(\tms1x00.RAM[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4575_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0196_),
    .Q(\tms1x00.RAM[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4576_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0197_),
    .Q(\tms1x00.RAM[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4577_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0198_),
    .Q(\tms1x00.RAM[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4578_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0199_),
    .Q(\tms1x00.RAM[118][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4579_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0200_),
    .Q(\tms1x00.RAM[118][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4580_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0201_),
    .Q(\tms1x00.RAM[118][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4581_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0202_),
    .Q(\tms1x00.RAM[118][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4582_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0203_),
    .Q(\tms1x00.RAM[117][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4583_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0204_),
    .Q(\tms1x00.RAM[117][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4584_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0205_),
    .Q(\tms1x00.RAM[117][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4585_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0206_),
    .Q(\tms1x00.RAM[117][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4586_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0207_),
    .Q(\tms1x00.RAM[116][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4587_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0208_),
    .Q(\tms1x00.RAM[116][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4588_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0209_),
    .Q(\tms1x00.RAM[116][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4589_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0210_),
    .Q(\tms1x00.RAM[116][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4590_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0211_),
    .Q(\tms1x00.RAM[115][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4591_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0212_),
    .Q(\tms1x00.RAM[115][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4592_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0213_),
    .Q(\tms1x00.RAM[115][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4593_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0214_),
    .Q(\tms1x00.RAM[115][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4594_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0215_),
    .Q(\tms1x00.RAM[126][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4595_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0216_),
    .Q(\tms1x00.RAM[126][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4596_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0217_),
    .Q(\tms1x00.RAM[126][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4597_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0218_),
    .Q(\tms1x00.RAM[126][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4598_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0219_),
    .Q(\tms1x00.RAM[125][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4599_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0220_),
    .Q(\tms1x00.RAM[125][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4600_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0221_),
    .Q(\tms1x00.RAM[125][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4601_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0222_),
    .Q(\tms1x00.RAM[125][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4602_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0223_),
    .Q(\tms1x00.RAM[25][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4603_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0224_),
    .Q(\tms1x00.RAM[25][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4604_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0225_),
    .Q(\tms1x00.RAM[25][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4605_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0226_),
    .Q(\tms1x00.RAM[25][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4606_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0227_),
    .Q(\tms1x00.RAM[24][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4607_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0228_),
    .Q(\tms1x00.RAM[24][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4608_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0229_),
    .Q(\tms1x00.RAM[24][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4609_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0230_),
    .Q(\tms1x00.RAM[24][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4610_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0231_),
    .Q(\tms1x00.RAM[28][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4611_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0232_),
    .Q(\tms1x00.RAM[28][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4612_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0233_),
    .Q(\tms1x00.RAM[28][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4613_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0234_),
    .Q(\tms1x00.RAM[28][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4614_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0235_),
    .Q(\tms1x00.RAM[27][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4615_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0236_),
    .Q(\tms1x00.RAM[27][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4616_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0237_),
    .Q(\tms1x00.RAM[27][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4617_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0238_),
    .Q(\tms1x00.RAM[27][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4618_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0239_),
    .Q(\tms1x00.RAM[26][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4619_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0240_),
    .Q(\tms1x00.RAM[26][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4620_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0241_),
    .Q(\tms1x00.RAM[26][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4621_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0242_),
    .Q(\tms1x00.RAM[26][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4622_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0243_),
    .Q(\tms1x00.RAM[32][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4623_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0244_),
    .Q(\tms1x00.RAM[32][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4624_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0245_),
    .Q(\tms1x00.RAM[32][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4625_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0246_),
    .Q(\tms1x00.RAM[32][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4626_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0247_),
    .Q(\tms1x00.RAM[31][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4627_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0248_),
    .Q(\tms1x00.RAM[31][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4628_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0249_),
    .Q(\tms1x00.RAM[31][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4629_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0250_),
    .Q(\tms1x00.RAM[31][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4630_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0251_),
    .Q(\tms1x00.RAM[30][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4631_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0252_),
    .Q(\tms1x00.RAM[30][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4632_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0253_),
    .Q(\tms1x00.RAM[30][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4633_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0254_),
    .Q(\tms1x00.RAM[30][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4634_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0255_),
    .Q(\tms1x00.RAM[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4635_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0256_),
    .Q(\tms1x00.RAM[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4636_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0257_),
    .Q(\tms1x00.RAM[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4637_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0258_),
    .Q(\tms1x00.RAM[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4638_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0259_),
    .Q(\tms1x00.RAM[37][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4639_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0260_),
    .Q(\tms1x00.RAM[37][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4640_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0261_),
    .Q(\tms1x00.RAM[37][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4641_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0262_),
    .Q(\tms1x00.RAM[37][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4642_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0263_),
    .Q(\tms1x00.RAM[36][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4643_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0264_),
    .Q(\tms1x00.RAM[36][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4644_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0265_),
    .Q(\tms1x00.RAM[36][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4645_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0266_),
    .Q(\tms1x00.RAM[36][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4646_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0267_),
    .Q(\tms1x00.RAM[35][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4647_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0268_),
    .Q(\tms1x00.RAM[35][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4648_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0269_),
    .Q(\tms1x00.RAM[35][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4649_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0270_),
    .Q(\tms1x00.RAM[35][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4650_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0271_),
    .Q(\tms1x00.RAM[34][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4651_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0272_),
    .Q(\tms1x00.RAM[34][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4652_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0273_),
    .Q(\tms1x00.RAM[34][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4653_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0274_),
    .Q(\tms1x00.RAM[34][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4654_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0275_),
    .Q(\tms1x00.RAM[33][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4655_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0276_),
    .Q(\tms1x00.RAM[33][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4656_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0277_),
    .Q(\tms1x00.RAM[33][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4657_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0278_),
    .Q(\tms1x00.RAM[33][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4658_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0279_),
    .Q(\tms1x00.RAM[41][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4659_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0280_),
    .Q(\tms1x00.RAM[41][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4660_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0281_),
    .Q(\tms1x00.RAM[41][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4661_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0282_),
    .Q(\tms1x00.RAM[41][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4662_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0283_),
    .Q(\tms1x00.RAM[40][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4663_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0284_),
    .Q(\tms1x00.RAM[40][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4664_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0285_),
    .Q(\tms1x00.RAM[40][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4665_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0286_),
    .Q(\tms1x00.RAM[40][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4666_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0287_),
    .Q(\tms1x00.RAM[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4667_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0288_),
    .Q(\tms1x00.RAM[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4668_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0289_),
    .Q(\tms1x00.RAM[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4669_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0290_),
    .Q(\tms1x00.RAM[3][3] ));
 sky130_fd_sc_hd__dfxtp_2 _4670_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0042_),
    .Q(_0035_));
 sky130_fd_sc_hd__dfxtp_1 _4671_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0043_),
    .Q(_0036_));
 sky130_fd_sc_hd__dfxtp_1 _4672_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0044_),
    .Q(_0037_));
 sky130_fd_sc_hd__dfxtp_2 _4673_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0045_),
    .Q(_0038_));
 sky130_fd_sc_hd__dfxtp_1 _4674_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0046_),
    .Q(_0039_));
 sky130_fd_sc_hd__dfxtp_4 _4675_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0047_),
    .Q(_0040_));
 sky130_fd_sc_hd__dfxtp_1 _4676_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0048_),
    .Q(_0041_));
 sky130_fd_sc_hd__dfxtp_1 _4677_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0291_),
    .Q(\tms1x00.RAM[38][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4678_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0292_),
    .Q(\tms1x00.RAM[38][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4679_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0293_),
    .Q(\tms1x00.RAM[38][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4680_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0294_),
    .Q(\tms1x00.RAM[38][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4681_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0295_),
    .Q(\tms1x00.RAM[45][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4682_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0296_),
    .Q(\tms1x00.RAM[45][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4683_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0297_),
    .Q(\tms1x00.RAM[45][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4684_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0298_),
    .Q(\tms1x00.RAM[45][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4685_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0299_),
    .Q(\tms1x00.RAM[44][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4686_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0300_),
    .Q(\tms1x00.RAM[44][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4687_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0301_),
    .Q(\tms1x00.RAM[44][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4688_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0302_),
    .Q(\tms1x00.RAM[44][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4689_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0303_),
    .Q(\tms1x00.RAM[43][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4690_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0304_),
    .Q(\tms1x00.RAM[43][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4691_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0305_),
    .Q(\tms1x00.RAM[43][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4692_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0306_),
    .Q(\tms1x00.RAM[43][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4693_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0307_),
    .Q(\tms1x00.RAM[42][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4694_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0308_),
    .Q(\tms1x00.RAM[42][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4695_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0309_),
    .Q(\tms1x00.RAM[42][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4696_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0310_),
    .Q(\tms1x00.RAM[42][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4697_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0311_),
    .Q(\tms1x00.RAM[50][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4698_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0312_),
    .Q(\tms1x00.RAM[50][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4699_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0313_),
    .Q(\tms1x00.RAM[50][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4700_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0314_),
    .Q(\tms1x00.RAM[50][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4701_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0315_),
    .Q(\tms1x00.RAM[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4702_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0316_),
    .Q(\tms1x00.RAM[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4703_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0317_),
    .Q(\tms1x00.RAM[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4704_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0318_),
    .Q(\tms1x00.RAM[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4705_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0319_),
    .Q(\tms1x00.RAM[48][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4706_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0320_),
    .Q(\tms1x00.RAM[48][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4707_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0321_),
    .Q(\tms1x00.RAM[48][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4708_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0322_),
    .Q(\tms1x00.RAM[48][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4709_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0323_),
    .Q(\tms1x00.RAM[47][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4710_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0324_),
    .Q(\tms1x00.RAM[47][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4711_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0325_),
    .Q(\tms1x00.RAM[47][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4712_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0326_),
    .Q(\tms1x00.RAM[47][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4713_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0327_),
    .Q(\tms1x00.RAM[46][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4714_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0328_),
    .Q(\tms1x00.RAM[46][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4715_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0329_),
    .Q(\tms1x00.RAM[46][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4716_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0330_),
    .Q(\tms1x00.RAM[46][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4717_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0331_),
    .Q(\tms1x00.RAM[54][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4718_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0332_),
    .Q(\tms1x00.RAM[54][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4719_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0333_),
    .Q(\tms1x00.RAM[54][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4720_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0334_),
    .Q(\tms1x00.RAM[54][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4721_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0335_),
    .Q(\tms1x00.RAM[53][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4722_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0336_),
    .Q(\tms1x00.RAM[53][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4723_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0337_),
    .Q(\tms1x00.RAM[53][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4724_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0338_),
    .Q(\tms1x00.RAM[53][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4725_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0339_),
    .Q(\tms1x00.RAM[52][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4726_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0340_),
    .Q(\tms1x00.RAM[52][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4727_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0341_),
    .Q(\tms1x00.RAM[52][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4728_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0342_),
    .Q(\tms1x00.RAM[52][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4729_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0343_),
    .Q(\tms1x00.RAM[51][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4730_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0344_),
    .Q(\tms1x00.RAM[51][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4731_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0345_),
    .Q(\tms1x00.RAM[51][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4732_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0346_),
    .Q(\tms1x00.RAM[51][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4733_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0347_),
    .Q(\tms1x00.RAM[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4734_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0348_),
    .Q(\tms1x00.RAM[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4735_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0349_),
    .Q(\tms1x00.RAM[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4736_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0350_),
    .Q(\tms1x00.RAM[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4737_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0351_),
    .Q(\tms1x00.RAM[58][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4738_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0352_),
    .Q(\tms1x00.RAM[58][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4739_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0353_),
    .Q(\tms1x00.RAM[58][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4740_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0354_),
    .Q(\tms1x00.RAM[58][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4741_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0355_),
    .Q(\tms1x00.RAM[57][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4742_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0356_),
    .Q(\tms1x00.RAM[57][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4743_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0357_),
    .Q(\tms1x00.RAM[57][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4744_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0358_),
    .Q(\tms1x00.RAM[57][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4745_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0359_),
    .Q(\tms1x00.RAM[56][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4746_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0360_),
    .Q(\tms1x00.RAM[56][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4747_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0361_),
    .Q(\tms1x00.RAM[56][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4748_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0362_),
    .Q(\tms1x00.RAM[56][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4749_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0363_),
    .Q(\tms1x00.RAM[55][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4750_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0364_),
    .Q(\tms1x00.RAM[55][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4751_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0365_),
    .Q(\tms1x00.RAM[55][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4752_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0366_),
    .Q(\tms1x00.RAM[55][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4753_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0367_),
    .Q(\tms1x00.RAM[63][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4754_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0368_),
    .Q(\tms1x00.RAM[63][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4755_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0369_),
    .Q(\tms1x00.RAM[63][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4756_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0370_),
    .Q(\tms1x00.RAM[63][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4757_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0371_),
    .Q(\tms1x00.RAM[62][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4758_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0372_),
    .Q(\tms1x00.RAM[62][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4759_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0373_),
    .Q(\tms1x00.RAM[62][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4760_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0374_),
    .Q(\tms1x00.RAM[62][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4761_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0375_),
    .Q(\tms1x00.RAM[61][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4762_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0376_),
    .Q(\tms1x00.RAM[61][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4763_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0377_),
    .Q(\tms1x00.RAM[61][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4764_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0378_),
    .Q(\tms1x00.RAM[61][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4765_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0379_),
    .Q(\tms1x00.RAM[60][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4766_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0380_),
    .Q(\tms1x00.RAM[60][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4767_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0381_),
    .Q(\tms1x00.RAM[60][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4768_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0382_),
    .Q(\tms1x00.RAM[60][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4769_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0383_),
    .Q(\tms1x00.RAM[67][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4770_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0384_),
    .Q(\tms1x00.RAM[67][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4771_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0385_),
    .Q(\tms1x00.RAM[67][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4772_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0386_),
    .Q(\tms1x00.RAM[67][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4773_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0387_),
    .Q(\tms1x00.RAM[66][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4774_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0388_),
    .Q(\tms1x00.RAM[66][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4775_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0389_),
    .Q(\tms1x00.RAM[66][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4776_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0390_),
    .Q(\tms1x00.RAM[66][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4777_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0391_),
    .Q(\tms1x00.RAM[65][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4778_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0392_),
    .Q(\tms1x00.RAM[65][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4779_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0393_),
    .Q(\tms1x00.RAM[65][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4780_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0394_),
    .Q(\tms1x00.RAM[65][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4781_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0395_),
    .Q(\tms1x00.RAM[64][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4782_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0396_),
    .Q(\tms1x00.RAM[64][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4783_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0397_),
    .Q(\tms1x00.RAM[64][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4784_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0398_),
    .Q(\tms1x00.RAM[64][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4785_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0399_),
    .Q(\tms1x00.RAM[72][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4786_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0400_),
    .Q(\tms1x00.RAM[72][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4787_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0401_),
    .Q(\tms1x00.RAM[72][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4788_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0402_),
    .Q(\tms1x00.RAM[72][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4789_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0403_),
    .Q(\tms1x00.RAM[71][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4790_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0404_),
    .Q(\tms1x00.RAM[71][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4791_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0405_),
    .Q(\tms1x00.RAM[71][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4792_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0406_),
    .Q(\tms1x00.RAM[71][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4793_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0407_),
    .Q(\tms1x00.RAM[70][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4794_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0408_),
    .Q(\tms1x00.RAM[70][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4795_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0409_),
    .Q(\tms1x00.RAM[70][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4796_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0410_),
    .Q(\tms1x00.RAM[70][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4797_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0411_),
    .Q(\tms1x00.RAM[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4798_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0412_),
    .Q(\tms1x00.RAM[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4799_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0413_),
    .Q(\tms1x00.RAM[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4800_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0414_),
    .Q(\tms1x00.RAM[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4801_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0415_),
    .Q(\tms1x00.RAM[68][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4802_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0416_),
    .Q(\tms1x00.RAM[68][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4803_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0417_),
    .Q(\tms1x00.RAM[68][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4804_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0418_),
    .Q(\tms1x00.RAM[68][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4805_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0419_),
    .Q(\tms1x00.RAM[76][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4806_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0420_),
    .Q(\tms1x00.RAM[76][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4807_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0421_),
    .Q(\tms1x00.RAM[76][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4808_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0422_),
    .Q(\tms1x00.RAM[76][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4809_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0423_),
    .Q(\tms1x00.RAM[75][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4810_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0424_),
    .Q(\tms1x00.RAM[75][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4811_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0425_),
    .Q(\tms1x00.RAM[75][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4812_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0426_),
    .Q(\tms1x00.RAM[75][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4813_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0427_),
    .Q(\tms1x00.RAM[74][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4814_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0428_),
    .Q(\tms1x00.RAM[74][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4815_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0429_),
    .Q(\tms1x00.RAM[74][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4816_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0430_),
    .Q(\tms1x00.RAM[74][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4817_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0431_),
    .Q(\tms1x00.RAM[73][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4818_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0432_),
    .Q(\tms1x00.RAM[73][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4819_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0433_),
    .Q(\tms1x00.RAM[73][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4820_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0434_),
    .Q(\tms1x00.RAM[73][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4821_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0435_),
    .Q(\tms1x00.RAM[80][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4822_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0436_),
    .Q(\tms1x00.RAM[80][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4823_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0437_),
    .Q(\tms1x00.RAM[80][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4824_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0438_),
    .Q(\tms1x00.RAM[80][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4825_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0439_),
    .Q(\tms1x00.RAM[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4826_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0440_),
    .Q(\tms1x00.RAM[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4827_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0441_),
    .Q(\tms1x00.RAM[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4828_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0442_),
    .Q(\tms1x00.RAM[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4829_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0443_),
    .Q(\tms1x00.RAM[78][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4830_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0444_),
    .Q(\tms1x00.RAM[78][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4831_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0445_),
    .Q(\tms1x00.RAM[78][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4832_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0446_),
    .Q(\tms1x00.RAM[78][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4833_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0447_),
    .Q(\tms1x00.RAM[77][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4834_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0448_),
    .Q(\tms1x00.RAM[77][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4835_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0449_),
    .Q(\tms1x00.RAM[77][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4836_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0450_),
    .Q(\tms1x00.RAM[77][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4837_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0451_),
    .Q(\tms1x00.RAM[85][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4838_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0452_),
    .Q(\tms1x00.RAM[85][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4839_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0453_),
    .Q(\tms1x00.RAM[85][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4840_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0454_),
    .Q(\tms1x00.RAM[85][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4841_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0455_),
    .Q(\tms1x00.RAM[84][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4842_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0456_),
    .Q(\tms1x00.RAM[84][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4843_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0457_),
    .Q(\tms1x00.RAM[84][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4844_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0458_),
    .Q(\tms1x00.RAM[84][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4845_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0459_),
    .Q(\tms1x00.RAM[83][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4846_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0460_),
    .Q(\tms1x00.RAM[83][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4847_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0461_),
    .Q(\tms1x00.RAM[83][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4848_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0462_),
    .Q(\tms1x00.RAM[83][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4849_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0463_),
    .Q(\tms1x00.RAM[82][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4850_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0464_),
    .Q(\tms1x00.RAM[82][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4851_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0465_),
    .Q(\tms1x00.RAM[82][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4852_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0466_),
    .Q(\tms1x00.RAM[82][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4853_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0467_),
    .Q(\tms1x00.RAM[81][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4854_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0468_),
    .Q(\tms1x00.RAM[81][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4855_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0469_),
    .Q(\tms1x00.RAM[81][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4856_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0470_),
    .Q(\tms1x00.RAM[81][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4857_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0471_),
    .Q(\tms1x00.RAM[86][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4858_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0472_),
    .Q(\tms1x00.RAM[86][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4859_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0473_),
    .Q(\tms1x00.RAM[86][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4860_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0474_),
    .Q(\tms1x00.RAM[86][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4861_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0475_),
    .Q(\tms1x00.RAM[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4862_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0476_),
    .Q(\tms1x00.RAM[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4863_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0477_),
    .Q(\tms1x00.RAM[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4864_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0478_),
    .Q(\tms1x00.RAM[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4865_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0479_),
    .Q(\tms1x00.RAM[88][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4866_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0480_),
    .Q(\tms1x00.RAM[88][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4867_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0481_),
    .Q(\tms1x00.RAM[88][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4868_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0482_),
    .Q(\tms1x00.RAM[88][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4869_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0483_),
    .Q(\tms1x00.RAM[87][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4870_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0484_),
    .Q(\tms1x00.RAM[87][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4871_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0485_),
    .Q(\tms1x00.RAM[87][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4872_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0486_),
    .Q(\tms1x00.RAM[87][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4873_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0487_),
    .Q(\tms1x00.RAM[94][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4874_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0488_),
    .Q(\tms1x00.RAM[94][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4875_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0489_),
    .Q(\tms1x00.RAM[94][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4876_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0490_),
    .Q(\tms1x00.RAM[94][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4877_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0491_),
    .Q(\tms1x00.RAM[93][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4878_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0492_),
    .Q(\tms1x00.RAM[93][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4879_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0493_),
    .Q(\tms1x00.RAM[93][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4880_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0494_),
    .Q(\tms1x00.RAM[93][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4881_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0495_),
    .Q(\tms1x00.RAM[92][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4882_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0496_),
    .Q(\tms1x00.RAM[92][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4883_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0497_),
    .Q(\tms1x00.RAM[92][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4884_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0498_),
    .Q(\tms1x00.RAM[92][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4885_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0499_),
    .Q(\tms1x00.RAM[91][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4886_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0500_),
    .Q(\tms1x00.RAM[91][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4887_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0501_),
    .Q(\tms1x00.RAM[91][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4888_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0502_),
    .Q(\tms1x00.RAM[91][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4889_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0503_),
    .Q(\tms1x00.RAM[90][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4890_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0504_),
    .Q(\tms1x00.RAM[90][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4891_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0505_),
    .Q(\tms1x00.RAM[90][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4892_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0506_),
    .Q(\tms1x00.RAM[90][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4893_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0507_),
    .Q(\tms1x00.RAM[23][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4894_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0508_),
    .Q(\tms1x00.RAM[23][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4895_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0509_),
    .Q(\tms1x00.RAM[23][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4896_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0510_),
    .Q(\tms1x00.RAM[23][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4897_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0511_),
    .Q(\tms1x00.ram_addr_buff[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4898_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0512_),
    .Q(\tms1x00.ram_addr_buff[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4899_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0513_),
    .Q(\tms1x00.ram_addr_buff[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4900_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0514_),
    .Q(\tms1x00.ram_addr_buff[3] ));
 sky130_fd_sc_hd__dfxtp_4 _4901_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0515_),
    .Q(\tms1x00.ram_addr_buff[4] ));
 sky130_fd_sc_hd__dfxtp_4 _4902_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0516_),
    .Q(\tms1x00.ram_addr_buff[5] ));
 sky130_fd_sc_hd__dfxtp_4 _4903_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0517_),
    .Q(\tms1x00.ram_addr_buff[6] ));
 sky130_fd_sc_hd__dfxtp_1 _4904_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0518_),
    .Q(\tms1x00.wb_step_state ));
 sky130_fd_sc_hd__dfxtp_2 _4905_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0519_),
    .Q(net93));
 sky130_fd_sc_hd__dfxtp_1 _4906_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0520_),
    .Q(\tms1x00.ins_in[0] ));
 sky130_fd_sc_hd__dfxtp_2 _4907_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0521_),
    .Q(\tms1x00.ins_in[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4908_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0522_),
    .Q(\tms1x00.ins_in[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4909_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0523_),
    .Q(\tms1x00.ins_in[3] ));
 sky130_fd_sc_hd__dfxtp_4 _4910_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0524_),
    .Q(\tms1x00.ins_in[4] ));
 sky130_fd_sc_hd__dfxtp_2 _4911_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0525_),
    .Q(\tms1x00.ins_in[5] ));
 sky130_fd_sc_hd__dfxtp_1 _4912_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0526_),
    .Q(\tms1x00.ins_in[6] ));
 sky130_fd_sc_hd__dfxtp_1 _4913_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0527_),
    .Q(\tms1x00.ins_in[7] ));
 sky130_fd_sc_hd__dfxtp_2 _4914_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0528_),
    .Q(net74));
 sky130_fd_sc_hd__dfxtp_4 _4915_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0529_),
    .Q(net75));
 sky130_fd_sc_hd__dfxtp_4 _4916_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0530_),
    .Q(net76));
 sky130_fd_sc_hd__dfxtp_1 _4917_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(\tms1x00.K_in[0] ),
    .Q(\tms1x00.K_latch[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4918_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(\tms1x00.K_in[1] ),
    .Q(\tms1x00.K_latch[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4919_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(\tms1x00.K_in[2] ),
    .Q(\tms1x00.K_latch[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4920_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(\tms1x00.K_in[3] ),
    .Q(\tms1x00.K_latch[3] ));
 sky130_fd_sc_hd__dfxtp_2 _4921_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0531_),
    .Q(net78));
 sky130_fd_sc_hd__dfxtp_2 _4922_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0532_),
    .Q(net79));
 sky130_fd_sc_hd__dfxtp_2 _4923_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0533_),
    .Q(net80));
 sky130_fd_sc_hd__dfxtp_2 _4924_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0534_),
    .Q(net81));
 sky130_fd_sc_hd__dfxtp_2 _4925_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0535_),
    .Q(net82));
 sky130_fd_sc_hd__dfxtp_2 _4926_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0536_),
    .Q(net83));
 sky130_fd_sc_hd__dfxtp_2 _4927_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0537_),
    .Q(net84));
 sky130_fd_sc_hd__dfxtp_2 _4928_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0538_),
    .Q(net85));
 sky130_fd_sc_hd__dfxtp_2 _4929_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0539_),
    .Q(net86));
 sky130_fd_sc_hd__dfxtp_2 _4930_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0540_),
    .Q(net87));
 sky130_fd_sc_hd__dfxtp_2 _4931_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0541_),
    .Q(net88));
 sky130_fd_sc_hd__dfxtp_2 _4932_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0542_),
    .Q(net89));
 sky130_fd_sc_hd__dfxtp_2 _4933_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0543_),
    .Q(net90));
 sky130_fd_sc_hd__dfxtp_2 _4934_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0544_),
    .Q(net91));
 sky130_fd_sc_hd__dfxtp_4 _4935_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0545_),
    .Q(net92));
 sky130_fd_sc_hd__dfxtp_2 _4936_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0546_),
    .Q(net69));
 sky130_fd_sc_hd__dfxtp_2 _4937_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0547_),
    .Q(net70));
 sky130_fd_sc_hd__dfxtp_2 _4938_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0548_),
    .Q(net71));
 sky130_fd_sc_hd__dfxtp_2 _4939_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0549_),
    .Q(net72));
 sky130_fd_sc_hd__dfxtp_2 _4940_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0550_),
    .Q(net73));
 sky130_fd_sc_hd__dfxtp_1 _4941_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0551_),
    .Q(\tms1x00.CL ));
 sky130_fd_sc_hd__dfxtp_1 _4942_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0552_),
    .Q(\tms1x00.status ));
 sky130_fd_sc_hd__dfxtp_1 _4943_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0553_),
    .Q(\tms1x00.SR[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4944_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0554_),
    .Q(\tms1x00.SR[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4945_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0555_),
    .Q(\tms1x00.SR[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4946_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0556_),
    .Q(\tms1x00.SR[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4947_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0557_),
    .Q(\tms1x00.SR[4] ));
 sky130_fd_sc_hd__dfxtp_1 _4948_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0558_),
    .Q(\tms1x00.SR[5] ));
 sky130_fd_sc_hd__dfxtp_1 _4949_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0559_),
    .Q(\tms1x00.PB[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4950_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0560_),
    .Q(\tms1x00.PB[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4951_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0561_),
    .Q(\tms1x00.PB[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4952_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0562_),
    .Q(\tms1x00.PB[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4953_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0563_),
    .Q(\tms1x00.PA[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4954_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0564_),
    .Q(\tms1x00.PA[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4955_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0565_),
    .Q(\tms1x00.PA[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4956_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0566_),
    .Q(\tms1x00.PA[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4957_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0567_),
    .Q(\tms1x00.P[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4958_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0568_),
    .Q(\tms1x00.P[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4959_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0569_),
    .Q(\tms1x00.P[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4960_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0570_),
    .Q(\tms1x00.P[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4961_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0571_),
    .Q(\tms1x00.PC[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4962_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0572_),
    .Q(\tms1x00.PC[1] ));
 sky130_fd_sc_hd__dfxtp_2 _4963_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0573_),
    .Q(\tms1x00.PC[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4964_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0574_),
    .Q(\tms1x00.PC[3] ));
 sky130_fd_sc_hd__dfxtp_2 _4965_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0575_),
    .Q(\tms1x00.PC[4] ));
 sky130_fd_sc_hd__dfxtp_1 _4966_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0576_),
    .Q(\tms1x00.PC[5] ));
 sky130_fd_sc_hd__dfxtp_2 _4967_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0577_),
    .Q(\tms1x00.Y[0] ));
 sky130_fd_sc_hd__dfxtp_2 _4968_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0578_),
    .Q(\tms1x00.Y[1] ));
 sky130_fd_sc_hd__dfxtp_2 _4969_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0579_),
    .Q(\tms1x00.Y[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4970_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0580_),
    .Q(\tms1x00.Y[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4971_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0581_),
    .Q(\tms1x00.X[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4972_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0582_),
    .Q(\tms1x00.X[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4973_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0583_),
    .Q(\tms1x00.X[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4974_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0584_),
    .Q(\tms1x00.N[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4975_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0585_),
    .Q(\tms1x00.N[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4976_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0586_),
    .Q(\tms1x00.N[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4977_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0587_),
    .Q(\tms1x00.N[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4978_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0588_),
    .Q(\tms1x00.A[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4979_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0589_),
    .Q(\tms1x00.A[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4980_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0590_),
    .Q(\tms1x00.A[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4981_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0591_),
    .Q(\tms1x00.A[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4982_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0592_),
    .Q(\tms1x00.RAM[119][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4983_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0593_),
    .Q(\tms1x00.RAM[119][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4984_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0594_),
    .Q(\tms1x00.RAM[119][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4985_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0595_),
    .Q(\tms1x00.RAM[119][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4986_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0596_),
    .Q(\tms1x00.RAM[39][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4987_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0597_),
    .Q(\tms1x00.RAM[39][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4988_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0598_),
    .Q(\tms1x00.RAM[39][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4989_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0599_),
    .Q(\tms1x00.RAM[39][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4990_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0600_),
    .Q(\tms1x00.RAM[22][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4991_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0601_),
    .Q(\tms1x00.RAM[22][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4992_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0602_),
    .Q(\tms1x00.RAM[22][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4993_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0603_),
    .Q(\tms1x00.RAM[22][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4994_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0604_),
    .Q(\tms1x00.RAM[29][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4995_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0605_),
    .Q(\tms1x00.RAM[29][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4996_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0606_),
    .Q(\tms1x00.RAM[29][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4997_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0607_),
    .Q(\tms1x00.RAM[29][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4998_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0608_),
    .Q(\tms1x00.RAM[21][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4999_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0609_),
    .Q(\tms1x00.RAM[21][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5000_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0610_),
    .Q(\tms1x00.RAM[21][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5001_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0611_),
    .Q(\tms1x00.RAM[21][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5002_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0612_),
    .Q(\tms1x00.RAM[16][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5003_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0613_),
    .Q(\tms1x00.RAM[16][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5004_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0614_),
    .Q(\tms1x00.RAM[16][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5005_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0615_),
    .Q(\tms1x00.RAM[16][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5006_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0616_),
    .Q(\tms1x00.RAM[20][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5007_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0617_),
    .Q(\tms1x00.RAM[20][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5008_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0618_),
    .Q(\tms1x00.RAM[20][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5009_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0619_),
    .Q(\tms1x00.RAM[20][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5010_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0620_),
    .Q(\tms1x00.RAM[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5011_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0621_),
    .Q(\tms1x00.RAM[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5012_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0622_),
    .Q(\tms1x00.RAM[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5013_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0623_),
    .Q(\tms1x00.RAM[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5014_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0624_),
    .Q(\tms1x00.RAM[127][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5015_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0625_),
    .Q(\tms1x00.RAM[127][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5016_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0626_),
    .Q(\tms1x00.RAM[127][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5017_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0627_),
    .Q(\tms1x00.RAM[127][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5018_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0628_),
    .Q(\tms1x00.RAM[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5019_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0629_),
    .Q(\tms1x00.RAM[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5020_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0630_),
    .Q(\tms1x00.RAM[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5021_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0631_),
    .Q(\tms1x00.RAM[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5022_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0632_),
    .Q(\tms1x00.RAM[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5023_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0633_),
    .Q(\tms1x00.RAM[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5024_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0634_),
    .Q(\tms1x00.RAM[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5025_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0635_),
    .Q(\tms1x00.RAM[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5026_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0636_),
    .Q(\tms1x00.RAM[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5027_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0637_),
    .Q(\tms1x00.RAM[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5028_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0638_),
    .Q(\tms1x00.RAM[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5029_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0639_),
    .Q(\tms1x00.RAM[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5030_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0640_),
    .Q(\tms1x00.RAM[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5031_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0641_),
    .Q(\tms1x00.RAM[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5032_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0642_),
    .Q(\tms1x00.RAM[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5033_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0643_),
    .Q(\tms1x00.RAM[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5034_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0644_),
    .Q(\tms1x00.RAM[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5035_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0645_),
    .Q(\tms1x00.RAM[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5036_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0646_),
    .Q(\tms1x00.RAM[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5037_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0647_),
    .Q(\tms1x00.RAM[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5038_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0648_),
    .Q(net95));
 sky130_fd_sc_hd__dfxtp_1 _5039_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0649_),
    .Q(net96));
 sky130_fd_sc_hd__dfxtp_1 _5040_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0650_),
    .Q(net97));
 sky130_fd_sc_hd__dfxtp_1 _5041_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0651_),
    .Q(net98));
 sky130_fd_sc_hd__dfxtp_1 _5042_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0652_),
    .Q(net99));
 sky130_fd_sc_hd__dfxtp_1 _5043_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0653_),
    .Q(net100));
 sky130_fd_sc_hd__dfxtp_1 _5044_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0654_),
    .Q(net101));
 sky130_fd_sc_hd__dfxtp_1 _5045_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0655_),
    .Q(net102));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_191 (.HI(net191));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_192 (.HI(net192));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_193 (.HI(net193));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_194 (.HI(net194));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_195 (.HI(net195));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_196 (.HI(net196));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_197 (.HI(net197));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_198 (.HI(net198));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_199 (.HI(net199));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_150 (.LO(net150));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_151 (.LO(net151));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_152 (.LO(net152));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_153 (.LO(net153));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_154 (.LO(net154));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_155 (.LO(net155));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_156 (.LO(net156));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_157 (.LO(net157));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_158 (.LO(net158));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_159 (.LO(net159));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_160 (.LO(net160));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_161 (.LO(net161));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_162 (.LO(net162));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_163 (.LO(net163));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_164 (.LO(net164));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_165 (.LO(net165));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_166 (.LO(net166));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_167 (.LO(net167));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_168 (.LO(net168));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_169 (.LO(net169));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_170 (.LO(net170));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_171 (.LO(net171));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_172 (.LO(net172));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_173 (.LO(net173));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_174 (.LO(net174));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_175 (.LO(net175));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_176 (.LO(net176));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_177 (.LO(net177));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_178 (.LO(net178));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_179 (.LO(net179));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_180 (.LO(net180));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_181 (.LO(net181));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_182 (.LO(net182));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_183 (.LO(net183));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_184 (.LO(net184));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_185 (.LO(net185));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_186 (.LO(net186));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_187 (.LO(net187));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_188 (.LO(net188));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_189 (.LO(net189));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_190 (.HI(net190));
 sky130_fd_sc_hd__clkbuf_2 _5097_ (.A(net50),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_2 _5098_ (.A(net51),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_2 _5099_ (.A(net52),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_2 _5100_ (.A(net53),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_2 _5101_ (.A(net54),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_2 _5102_ (.A(net55),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_2 _5103_ (.A(net56),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_2 _5104_ (.A(net57),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_2 _5105_ (.A(net47),
    .X(net112));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(io_in[5]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(io_in[6]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(io_in[7]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(io_in[8]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(io_in[9]),
    .X(net5));
 sky130_fd_sc_hd__dlymetal6s2s_1 input6 (.A(oram_value[0]),
    .X(net6));
 sky130_fd_sc_hd__dlymetal6s2s_1 input7 (.A(oram_value[1]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(oram_value[2]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(oram_value[3]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(oram_value[4]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(oram_value[5]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(oram_value[6]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(oram_value[7]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(ram_val[0]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(ram_val[10]),
    .X(net15));
 sky130_fd_sc_hd__dlymetal6s2s_1 input16 (.A(ram_val[11]),
    .X(net16));
 sky130_fd_sc_hd__dlymetal6s2s_1 input17 (.A(ram_val[12]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(ram_val[13]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(ram_val[14]),
    .X(net19));
 sky130_fd_sc_hd__dlymetal6s2s_1 input20 (.A(ram_val[15]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(ram_val[16]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(ram_val[17]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(ram_val[18]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(ram_val[19]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(ram_val[1]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(ram_val[20]),
    .X(net26));
 sky130_fd_sc_hd__dlymetal6s2s_1 input27 (.A(ram_val[21]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(ram_val[22]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(ram_val[23]),
    .X(net29));
 sky130_fd_sc_hd__dlymetal6s2s_1 input30 (.A(ram_val[24]),
    .X(net30));
 sky130_fd_sc_hd__dlymetal6s2s_1 input31 (.A(ram_val[25]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(ram_val[26]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(ram_val[27]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(ram_val[28]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(ram_val[29]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 input36 (.A(ram_val[2]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(ram_val[30]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(ram_val[31]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_2 input39 (.A(ram_val[3]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_2 input40 (.A(ram_val[4]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_2 input41 (.A(ram_val[5]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_2 input42 (.A(ram_val[6]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_2 input43 (.A(ram_val[7]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_2 input44 (.A(ram_val[8]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_2 input45 (.A(ram_val[9]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_4 input46 (.A(wb_rst_i),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(wbs_adr_i[10]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(wbs_adr_i[16]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_4 input49 (.A(wbs_adr_i[23]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(wbs_adr_i[2]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(wbs_adr_i[3]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(wbs_adr_i[4]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(wbs_adr_i[5]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(wbs_adr_i[6]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(wbs_adr_i[7]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(wbs_adr_i[8]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 input57 (.A(wbs_adr_i[9]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(wbs_cyc_i),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(wbs_dat_i[0]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(wbs_dat_i[10]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(wbs_dat_i[11]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(wbs_dat_i[1]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 input63 (.A(wbs_dat_i[2]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 input64 (.A(wbs_dat_i[3]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 input65 (.A(wbs_dat_i[8]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 input66 (.A(wbs_dat_i[9]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 input67 (.A(wbs_stb_i),
    .X(net67));
 sky130_fd_sc_hd__dlymetal6s2s_1 input68 (.A(wbs_we_i),
    .X(net68));
 sky130_fd_sc_hd__buf_2 output69 (.A(net69),
    .X(io_out[10]));
 sky130_fd_sc_hd__buf_2 output70 (.A(net70),
    .X(io_out[11]));
 sky130_fd_sc_hd__buf_2 output71 (.A(net71),
    .X(io_out[12]));
 sky130_fd_sc_hd__buf_2 output72 (.A(net72),
    .X(io_out[13]));
 sky130_fd_sc_hd__buf_2 output73 (.A(net73),
    .X(io_out[14]));
 sky130_fd_sc_hd__buf_2 output74 (.A(net74),
    .X(io_out[15]));
 sky130_fd_sc_hd__buf_2 output75 (.A(net75),
    .X(io_out[16]));
 sky130_fd_sc_hd__buf_2 output76 (.A(net76),
    .X(io_out[17]));
 sky130_fd_sc_hd__buf_2 output77 (.A(net77),
    .X(io_out[18]));
 sky130_fd_sc_hd__buf_2 output78 (.A(net78),
    .X(io_out[19]));
 sky130_fd_sc_hd__buf_2 output79 (.A(net79),
    .X(io_out[20]));
 sky130_fd_sc_hd__buf_2 output80 (.A(net80),
    .X(io_out[21]));
 sky130_fd_sc_hd__buf_2 output81 (.A(net81),
    .X(io_out[22]));
 sky130_fd_sc_hd__buf_2 output82 (.A(net82),
    .X(io_out[23]));
 sky130_fd_sc_hd__buf_2 output83 (.A(net83),
    .X(io_out[24]));
 sky130_fd_sc_hd__buf_2 output84 (.A(net84),
    .X(io_out[25]));
 sky130_fd_sc_hd__buf_2 output85 (.A(net85),
    .X(io_out[26]));
 sky130_fd_sc_hd__buf_2 output86 (.A(net86),
    .X(io_out[27]));
 sky130_fd_sc_hd__buf_2 output87 (.A(net87),
    .X(io_out[28]));
 sky130_fd_sc_hd__buf_2 output88 (.A(net88),
    .X(io_out[29]));
 sky130_fd_sc_hd__buf_2 output89 (.A(net89),
    .X(io_out[30]));
 sky130_fd_sc_hd__buf_2 output90 (.A(net90),
    .X(io_out[31]));
 sky130_fd_sc_hd__buf_2 output91 (.A(net91),
    .X(io_out[32]));
 sky130_fd_sc_hd__buf_2 output92 (.A(net92),
    .X(io_out[33]));
 sky130_fd_sc_hd__buf_2 output93 (.A(net93),
    .X(io_out[36]));
 sky130_fd_sc_hd__buf_2 output94 (.A(net94),
    .X(io_out[37]));
 sky130_fd_sc_hd__buf_2 output95 (.A(net95),
    .X(oram_addr[0]));
 sky130_fd_sc_hd__buf_2 output96 (.A(net96),
    .X(oram_addr[1]));
 sky130_fd_sc_hd__buf_2 output97 (.A(net97),
    .X(oram_addr[2]));
 sky130_fd_sc_hd__buf_2 output98 (.A(net98),
    .X(oram_addr[3]));
 sky130_fd_sc_hd__buf_2 output99 (.A(net99),
    .X(oram_addr[4]));
 sky130_fd_sc_hd__buf_2 output100 (.A(net100),
    .X(oram_addr[5]));
 sky130_fd_sc_hd__buf_2 output101 (.A(net101),
    .X(oram_addr[6]));
 sky130_fd_sc_hd__buf_2 output102 (.A(net102),
    .X(oram_addr[7]));
 sky130_fd_sc_hd__buf_2 output103 (.A(net103),
    .X(oram_csb));
 sky130_fd_sc_hd__buf_2 output104 (.A(net104),
    .X(ram_adrb[0]));
 sky130_fd_sc_hd__buf_2 output105 (.A(net105),
    .X(ram_adrb[1]));
 sky130_fd_sc_hd__buf_2 output106 (.A(net106),
    .X(ram_adrb[2]));
 sky130_fd_sc_hd__buf_2 output107 (.A(net107),
    .X(ram_adrb[3]));
 sky130_fd_sc_hd__buf_2 output108 (.A(net108),
    .X(ram_adrb[4]));
 sky130_fd_sc_hd__buf_2 output109 (.A(net109),
    .X(ram_adrb[5]));
 sky130_fd_sc_hd__buf_2 output110 (.A(net110),
    .X(ram_adrb[6]));
 sky130_fd_sc_hd__buf_2 output111 (.A(net111),
    .X(ram_adrb[7]));
 sky130_fd_sc_hd__buf_2 output112 (.A(net112),
    .X(ram_adrb[8]));
 sky130_fd_sc_hd__buf_2 output113 (.A(net113),
    .X(ram_csb));
 sky130_fd_sc_hd__buf_2 output114 (.A(net114),
    .X(ram_web));
 sky130_fd_sc_hd__buf_2 output115 (.A(net115),
    .X(wbs_ack_o));
 sky130_fd_sc_hd__buf_2 output116 (.A(net116),
    .X(wbs_dat_o[0]));
 sky130_fd_sc_hd__buf_2 output117 (.A(net117),
    .X(wbs_dat_o[10]));
 sky130_fd_sc_hd__buf_2 output118 (.A(net118),
    .X(wbs_dat_o[11]));
 sky130_fd_sc_hd__buf_2 output119 (.A(net119),
    .X(wbs_dat_o[12]));
 sky130_fd_sc_hd__buf_2 output120 (.A(net120),
    .X(wbs_dat_o[13]));
 sky130_fd_sc_hd__buf_2 output121 (.A(net121),
    .X(wbs_dat_o[14]));
 sky130_fd_sc_hd__buf_2 output122 (.A(net122),
    .X(wbs_dat_o[15]));
 sky130_fd_sc_hd__buf_2 output123 (.A(net123),
    .X(wbs_dat_o[16]));
 sky130_fd_sc_hd__buf_2 output124 (.A(net124),
    .X(wbs_dat_o[17]));
 sky130_fd_sc_hd__buf_2 output125 (.A(net125),
    .X(wbs_dat_o[18]));
 sky130_fd_sc_hd__buf_2 output126 (.A(net126),
    .X(wbs_dat_o[19]));
 sky130_fd_sc_hd__buf_2 output127 (.A(net127),
    .X(wbs_dat_o[1]));
 sky130_fd_sc_hd__buf_2 output128 (.A(net128),
    .X(wbs_dat_o[20]));
 sky130_fd_sc_hd__buf_2 output129 (.A(net129),
    .X(wbs_dat_o[21]));
 sky130_fd_sc_hd__buf_2 output130 (.A(net130),
    .X(wbs_dat_o[22]));
 sky130_fd_sc_hd__buf_2 output131 (.A(net131),
    .X(wbs_dat_o[23]));
 sky130_fd_sc_hd__buf_2 output132 (.A(net132),
    .X(wbs_dat_o[24]));
 sky130_fd_sc_hd__buf_2 output133 (.A(net133),
    .X(wbs_dat_o[25]));
 sky130_fd_sc_hd__buf_2 output134 (.A(net134),
    .X(wbs_dat_o[26]));
 sky130_fd_sc_hd__buf_2 output135 (.A(net135),
    .X(wbs_dat_o[27]));
 sky130_fd_sc_hd__buf_2 output136 (.A(net136),
    .X(wbs_dat_o[28]));
 sky130_fd_sc_hd__buf_2 output137 (.A(net137),
    .X(wbs_dat_o[29]));
 sky130_fd_sc_hd__buf_2 output138 (.A(net138),
    .X(wbs_dat_o[2]));
 sky130_fd_sc_hd__buf_2 output139 (.A(net139),
    .X(wbs_dat_o[30]));
 sky130_fd_sc_hd__buf_2 output140 (.A(net140),
    .X(wbs_dat_o[31]));
 sky130_fd_sc_hd__buf_2 output141 (.A(net141),
    .X(wbs_dat_o[3]));
 sky130_fd_sc_hd__buf_2 output142 (.A(net142),
    .X(wbs_dat_o[4]));
 sky130_fd_sc_hd__buf_2 output143 (.A(net143),
    .X(wbs_dat_o[5]));
 sky130_fd_sc_hd__buf_2 output144 (.A(net144),
    .X(wbs_dat_o[6]));
 sky130_fd_sc_hd__buf_2 output145 (.A(net145),
    .X(wbs_dat_o[7]));
 sky130_fd_sc_hd__buf_2 output146 (.A(net146),
    .X(wbs_dat_o[8]));
 sky130_fd_sc_hd__buf_2 output147 (.A(net147),
    .X(wbs_dat_o[9]));
 sky130_fd_sc_hd__buf_4 fanout148 (.A(net94),
    .X(net148));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_149 (.LO(net149));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_21_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_23_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_25_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_26_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_28_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_29_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_32_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_33_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_34_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(feedback_delay),
    .X(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__2914__A0 (.DIODE(\K_override[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2248__A1 (.DIODE(\K_override[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2916__A0 (.DIODE(\K_override[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2250__A1 (.DIODE(\K_override[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2918__A0 (.DIODE(\K_override[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2252__A1 (.DIODE(\K_override[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2920__A0 (.DIODE(\K_override[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2254__A1 (.DIODE(\K_override[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2628__B1 (.DIODE(_0038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2501__B1 (.DIODE(_0038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2455__B1 (.DIODE(_0038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2413__A (.DIODE(_0038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2409__A (.DIODE(_0038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2381__A (.DIODE(_0038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2688__A (.DIODE(_0039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2509__A1 (.DIODE(_0039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2489__B1 (.DIODE(_0039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2428__A (.DIODE(_0039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2411__A (.DIODE(_0039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2830__A1 (.DIODE(_0040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2785__B1 (.DIODE(_0040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2734__A1 (.DIODE(_0040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2665__B1 (.DIODE(_0040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2637__A1 (.DIODE(_0040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2590__B1 (.DIODE(_0040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2568__B1 (.DIODE(_0040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2509__C1 (.DIODE(_0040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2464__C1 (.DIODE(_0040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2380__A (.DIODE(_0040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4963__D (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2221__S (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2219__S (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2217__S (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2215__S (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2213__S (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2211__S (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2209__S (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2207__S (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2205__S (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2203__S (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2204__A (.DIODE(_0669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2206__A (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2210__A (.DIODE(_0672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2216__A (.DIODE(_0675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2222__A (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2289__A2 (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2288__A2 (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2287__A2 (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2286__A2 (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2273__A (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2260__B (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2259__A (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2304__B (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2302__B (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2285__A (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2274__A (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2261__A (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4156__C1 (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4151__A_N (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4134__A (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4130__A (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3998__A1 (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3994__A (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3993__A (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3977__A (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2319__A_N (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2268__A1 (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2284__B1 (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2283__B1 (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2282__B1 (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2281__B1 (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2280__B1 (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2279__B1 (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2278__B1 (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2277__B1 (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2276__B1 (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2275__B1 (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2300__B (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2298__B (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2296__B (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2294__B (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2292__B (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2290__B (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2289__B1 (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2288__B1 (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2287__B1 (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2286__B1 (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2920__S (.DIODE(_0715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2918__S (.DIODE(_0715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2916__S (.DIODE(_0715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2914__S (.DIODE(_0715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2309__B (.DIODE(_0715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4087__A (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4070__A (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4043__A (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4031__A (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4022__A (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3995__A (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3979__A (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2371__A (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2341__A (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2321__A (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3991__A2 (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3989__A2 (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3985__S (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3984__A2 (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3982__A2 (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3980__A2 (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3974__S (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3971__S (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2321__B (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3956__S (.DIODE(_0726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3954__S (.DIODE(_0726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3952__S (.DIODE(_0726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2339__S (.DIODE(_0726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2337__S (.DIODE(_0726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2335__S (.DIODE(_0726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2333__S (.DIODE(_0726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2329__S (.DIODE(_0726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2326__S (.DIODE(_0726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2323__S (.DIODE(_0726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4145__A1 (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4052__B (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4049__B (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4038__B (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4035__B (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4017__A2 (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4008__B (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4004__B (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3956__A0 (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2329__A0 (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4219__A0 (.DIODE(_0732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4148__B2 (.DIODE(_0732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4041__A1 (.DIODE(_0732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4026__A (.DIODE(_0732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4021__A (.DIODE(_0732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4016__A (.DIODE(_0732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4014__A (.DIODE(_0732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4008__A (.DIODE(_0732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4004__A (.DIODE(_0732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2332__A (.DIODE(_0732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4240__B (.DIODE(_0738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4128__A (.DIODE(_0738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4126__A (.DIODE(_0738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4123__A (.DIODE(_0738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4103__B (.DIODE(_0738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4085__B (.DIODE(_0738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3969__S (.DIODE(_0738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2512__B (.DIODE(_0738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2378__A (.DIODE(_0738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2342__A (.DIODE(_0738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4222__D (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4075__A_N (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4072__A_N (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4068__A_N (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4065__A_N (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4061__A_N (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3971__A0 (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2515__B (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2362__C_N (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2357__B (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4191__C_N (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4114__B (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4080__B (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3991__A1 (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2832__A (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2736__B_N (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2639__A_N (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2511__A (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2379__A (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2354__A (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4191__A (.DIODE(_0748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4180__A1 (.DIODE(_0748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4080__C (.DIODE(_0748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3989__A1 (.DIODE(_0748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2832__B (.DIODE(_0748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2736__A (.DIODE(_0748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2639__B (.DIODE(_0748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2511__C (.DIODE(_0748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2379__B (.DIODE(_0748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2354__B (.DIODE(_0748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4053__B (.DIODE(_0752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4050__B (.DIODE(_0752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4042__B (.DIODE(_0752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4030__B (.DIODE(_0752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4008__C (.DIODE(_0752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4004__C (.DIODE(_0752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2358__A (.DIODE(_0752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4188__B1 (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4184__A1 (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4178__A1 (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4166__A1 (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4128__B (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4081__A (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4079__A (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3977__B (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2378__B (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2366__A (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4052__C (.DIODE(_0763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4049__C (.DIODE(_0763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4041__A2 (.DIODE(_0763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4029__A2 (.DIODE(_0763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4012__B (.DIODE(_0763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4007__C (.DIODE(_0763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2369__A (.DIODE(_0763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4231__C1 (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4229__C1 (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4220__A (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4214__A (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4206__A (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4198__A (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4189__B1 (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4034__C1 (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3966__B (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2372__C1 (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4156__A1 (.DIODE(_0768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4132__B (.DIODE(_0768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4059__B (.DIODE(_0768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2377__B (.DIODE(_0768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2809__C1 (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2765__C1 (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2713__C1 (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2689__C1 (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2636__A (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2510__A1 (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2465__A1 (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2801__C1 (.DIODE(_0775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2757__C1 (.DIODE(_0775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2705__C1 (.DIODE(_0775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2623__B1 (.DIODE(_0775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2552__A (.DIODE(_0775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2497__C1 (.DIODE(_0775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2488__C1 (.DIODE(_0775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2451__C1 (.DIODE(_0775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2440__C1 (.DIODE(_0775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2383__A (.DIODE(_0775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2745__C1 (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2733__A1 (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2669__C1 (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2664__A1 (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2653__C1 (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2608__B1 (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2589__C1 (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2542__B1 (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2475__A1 (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2412__A1 (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2500__S0 (.DIODE(_0777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2498__S0 (.DIODE(_0777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2495__S0 (.DIODE(_0777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2491__S0 (.DIODE(_0777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2444__S0 (.DIODE(_0777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2437__A (.DIODE(_0777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2415__A (.DIODE(_0777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2406__A (.DIODE(_0777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2395__A (.DIODE(_0777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2385__A (.DIODE(_0777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2805__S (.DIODE(_0778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2798__S (.DIODE(_0778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2760__A1 (.DIODE(_0778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2759__B_N (.DIODE(_0778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2631__S (.DIODE(_0778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2583__A (.DIODE(_0778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2503__A1 (.DIODE(_0778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2502__B_N (.DIODE(_0778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2389__S0 (.DIODE(_0778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2388__S0 (.DIODE(_0778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2500__S1 (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2498__S1 (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2495__S1 (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2491__S1 (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2457__A (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2449__S1 (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2444__S1 (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2438__A (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2407__A (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2387__A (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2815__S1 (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2804__B1 (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2633__S1 (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2630__B1 (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2618__S1 (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2476__S1 (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2416__S1 (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2398__A (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2389__S1 (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2388__S1 (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2827__A (.DIODE(_0783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2816__A (.DIODE(_0783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2782__A (.DIODE(_0783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2731__A (.DIODE(_0783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2722__A (.DIODE(_0783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2634__A1 (.DIODE(_0783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2626__A (.DIODE(_0783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2556__A (.DIODE(_0783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2468__S (.DIODE(_0783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2391__S (.DIODE(_0783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2806__B2 (.DIODE(_0786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2762__B2 (.DIODE(_0786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2755__A1 (.DIODE(_0786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2710__B2 (.DIODE(_0786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2703__A1 (.DIODE(_0786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2486__A1 (.DIODE(_0786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2472__A1 (.DIODE(_0786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2460__B2 (.DIODE(_0786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2436__A1 (.DIODE(_0786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2394__A (.DIODE(_0786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2822__B2 (.DIODE(_0787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2793__A1 (.DIODE(_0787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2777__B2 (.DIODE(_0787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2749__A1 (.DIODE(_0787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2697__A1 (.DIODE(_0787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2611__A1 (.DIODE(_0787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2606__A1 (.DIODE(_0787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2549__B2 (.DIODE(_0787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2534__A (.DIODE(_0787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2403__A1 (.DIODE(_0787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2796__S (.DIODE(_0788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2709__S (.DIODE(_0788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2702__S (.DIODE(_0788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2700__S (.DIODE(_0788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2684__A1 (.DIODE(_0788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2683__B_N (.DIODE(_0788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2633__S0 (.DIODE(_0788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2459__S (.DIODE(_0788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2399__S (.DIODE(_0788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2396__A (.DIODE(_0788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2776__S (.DIODE(_0789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2748__S (.DIODE(_0789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2716__S (.DIODE(_0789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2694__S (.DIODE(_0789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2672__S (.DIODE(_0789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2479__A1 (.DIODE(_0789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2478__B_N (.DIODE(_0789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2421__A1 (.DIODE(_0789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2418__B_N (.DIODE(_0789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2397__S (.DIODE(_0789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2820__B1 (.DIODE(_0791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2814__S1 (.DIODE(_0791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2599__S1 (.DIODE(_0791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2593__S1 (.DIODE(_0791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2592__S1 (.DIODE(_0791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2571__S1 (.DIODE(_0791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2569__S1 (.DIODE(_0791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2555__S1 (.DIODE(_0791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2554__S1 (.DIODE(_0791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2402__A1 (.DIODE(_0791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2806__C1 (.DIODE(_0794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2799__B1 (.DIODE(_0794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2710__C1 (.DIODE(_0794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2703__B1 (.DIODE(_0794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2632__C1 (.DIODE(_0794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2628__A1 (.DIODE(_0794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2604__A (.DIODE(_0794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2561__A (.DIODE(_0794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2455__A1 (.DIODE(_0794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2402__B1 (.DIODE(_0794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2768__A (.DIODE(_0798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2763__A1 (.DIODE(_0798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2705__B2 (.DIODE(_0798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2659__A (.DIODE(_0798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2621__A (.DIODE(_0798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2575__A (.DIODE(_0798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2497__A1 (.DIODE(_0798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2474__B2 (.DIODE(_0798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2451__A1 (.DIODE(_0798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2410__A1 (.DIODE(_0798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2758__S0 (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2667__S0 (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2658__S0 (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2651__S0 (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2616__S0 (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2574__S0 (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2563__A (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2494__S0 (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2443__S0 (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2408__S0 (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2682__S1 (.DIODE(_0800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2667__S1 (.DIODE(_0800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2658__S1 (.DIODE(_0800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2651__S1 (.DIODE(_0800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2616__S1 (.DIODE(_0800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2564__A (.DIODE(_0800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2494__S1 (.DIODE(_0800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2473__S1 (.DIODE(_0800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2443__S1 (.DIODE(_0800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2408__S1 (.DIODE(_0800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2763__C1 (.DIODE(_0802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2711__C1 (.DIODE(_0802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2687__C1 (.DIODE(_0802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2663__C1 (.DIODE(_0802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2619__B1 (.DIODE(_0802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2550__A (.DIODE(_0802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2493__C1 (.DIODE(_0802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2474__C1 (.DIODE(_0802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2446__C1 (.DIODE(_0802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2410__B1 (.DIODE(_0802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2784__B1 (.DIODE(_0804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2724__B1 (.DIODE(_0804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2664__B1 (.DIODE(_0804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2635__C1 (.DIODE(_0804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2624__C1 (.DIODE(_0804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2528__A (.DIODE(_0804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2508__C1 (.DIODE(_0804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2475__C1 (.DIODE(_0804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2463__C1 (.DIODE(_0804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2412__C1 (.DIODE(_0804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2828__C1 (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2817__C1 (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2807__C1 (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2783__C1 (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2732__C1 (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2723__C1 (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2600__C1 (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2581__C1 (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2489__A1 (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2441__A1 (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2757__B2 (.DIODE(_0807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2687__A1 (.DIODE(_0807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2681__B2 (.DIODE(_0807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2648__A (.DIODE(_0807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2619__A1 (.DIODE(_0807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2580__A (.DIODE(_0807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2488__B2 (.DIODE(_0807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2477__A (.DIODE(_0807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2440__B2 (.DIODE(_0807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2417__A (.DIODE(_0807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2680__S0 (.DIODE(_0808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2622__S0 (.DIODE(_0808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2618__S0 (.DIODE(_0808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2579__S0 (.DIODE(_0808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2553__A (.DIODE(_0808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2490__S0 (.DIODE(_0808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2476__S0 (.DIODE(_0808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2458__A1 (.DIODE(_0808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2456__B_N (.DIODE(_0808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2416__S0 (.DIODE(_0808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2760__B1 (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2684__B1 (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2661__S1 (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2506__S1 (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2503__B1 (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2461__S1 (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2454__S1 (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2452__S1 (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2429__A (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2420__A (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2767__S1 (.DIODE(_0813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2758__S1 (.DIODE(_0813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2743__S1 (.DIODE(_0813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2704__S1 (.DIODE(_0813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2677__A (.DIODE(_0813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2620__S1 (.DIODE(_0813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2574__S1 (.DIODE(_0813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2479__B1 (.DIODE(_0813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2448__S1 (.DIODE(_0813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2421__B1 (.DIODE(_0813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2676__S (.DIODE(_0815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2661__S0 (.DIODE(_0815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2506__S0 (.DIODE(_0815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2480__A (.DIODE(_0815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2461__S0 (.DIODE(_0815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2454__S0 (.DIODE(_0815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2452__S0 (.DIODE(_0815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2449__S0 (.DIODE(_0815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2447__A (.DIODE(_0815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2423__A (.DIODE(_0815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2823__S0 (.DIODE(_0816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2812__S0 (.DIODE(_0816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2810__S0 (.DIODE(_0816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2802__S0 (.DIODE(_0816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2800__S0 (.DIODE(_0816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2729__S0 (.DIODE(_0816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2720__S0 (.DIODE(_0816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2597__S (.DIODE(_0816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2558__S (.DIODE(_0816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2424__S (.DIODE(_0816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2799__A1 (.DIODE(_0818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2717__B2 (.DIODE(_0818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2673__A1 (.DIODE(_0818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2657__B2 (.DIODE(_0818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2632__B2 (.DIODE(_0818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2596__A (.DIODE(_0818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2588__B2 (.DIODE(_0818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2559__A (.DIODE(_0818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2482__B2 (.DIODE(_0818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2427__B2 (.DIODE(_0818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2668__A (.DIODE(_0819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2652__A (.DIODE(_0819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2623__A1 (.DIODE(_0819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2598__B1 (.DIODE(_0819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2588__C1 (.DIODE(_0819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2548__A (.DIODE(_0819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2493__A1 (.DIODE(_0819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2482__C1 (.DIODE(_0819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2446__A1 (.DIODE(_0819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2427__C1 (.DIODE(_0819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2818__B1 (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2808__A (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2785__A1 (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2764__A (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2733__B1 (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2712__A (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2665__A1 (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2577__B1 (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2464__A1 (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2441__B1 (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2753__A (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2727__S1 (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2725__S1 (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2718__S1 (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2706__S1 (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2660__S1 (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2540__A (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2484__A (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2470__A (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2432__A (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2781__S0 (.DIODE(_0823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2752__S (.DIODE(_0823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2730__S0 (.DIODE(_0823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2721__S0 (.DIODE(_0823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2685__S (.DIODE(_0823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2678__S (.DIODE(_0823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2625__S0 (.DIODE(_0823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2483__S (.DIODE(_0823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2469__S (.DIODE(_0823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2431__S (.DIODE(_0823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2826__S0 (.DIODE(_0826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2815__S0 (.DIODE(_0826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2761__S (.DIODE(_0826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2754__S (.DIODE(_0826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2627__S0 (.DIODE(_0826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2531__A (.DIODE(_0826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2504__S (.DIODE(_0826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2485__S (.DIODE(_0826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2471__S (.DIODE(_0826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2434__S (.DIODE(_0826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2762__C1 (.DIODE(_0828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2755__B1 (.DIODE(_0828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2505__C1 (.DIODE(_0828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2501__A1 (.DIODE(_0828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2496__A (.DIODE(_0828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2486__B1 (.DIODE(_0828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2472__B1 (.DIODE(_0828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2460__C1 (.DIODE(_0828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2450__A (.DIODE(_0828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2436__B1 (.DIODE(_0828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2756__S0 (.DIODE(_0830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2708__A1 (.DIODE(_0830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2707__B_N (.DIODE(_0830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2682__S0 (.DIODE(_0830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2647__S0 (.DIODE(_0830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2487__S0 (.DIODE(_0830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2473__S0 (.DIODE(_0830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2467__S0 (.DIODE(_0830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2466__S0 (.DIODE(_0830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2439__S0 (.DIODE(_0830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2756__S1 (.DIODE(_0831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2680__S1 (.DIODE(_0831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2647__S1 (.DIODE(_0831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2622__S1 (.DIODE(_0831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2579__S1 (.DIODE(_0831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2490__S1 (.DIODE(_0831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2487__S1 (.DIODE(_0831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2467__S1 (.DIODE(_0831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2466__S1 (.DIODE(_0831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2439__S1 (.DIODE(_0831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2804__A1 (.DIODE(_0840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2803__B_N (.DIODE(_0840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2767__S0 (.DIODE(_0840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2743__S0 (.DIODE(_0840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2704__S0 (.DIODE(_0840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2660__S0 (.DIODE(_0840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2630__A1 (.DIODE(_0840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2620__S0 (.DIODE(_0840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2539__A (.DIODE(_0840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2448__S0 (.DIODE(_0840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2451__A2 (.DIODE(_0841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2453__B (.DIODE(_0845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2826__S1 (.DIODE(_0850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2781__S1 (.DIODE(_0850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2730__S1 (.DIODE(_0850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2721__S1 (.DIODE(_0850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2708__B1 (.DIODE(_0850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2627__S1 (.DIODE(_0850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2625__S1 (.DIODE(_0850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2585__A (.DIODE(_0850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2535__A (.DIODE(_0850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2458__B1 (.DIODE(_0850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2462__A2 (.DIODE(_0854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4131__A (.DIODE(_0858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2514__A2 (.DIODE(_0858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2468__A0 (.DIODE(_0859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2468__A1 (.DIODE(_0860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2474__B1 (.DIODE(_0866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2778__S0 (.DIODE(_0873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2771__S0 (.DIODE(_0873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2727__S0 (.DIODE(_0873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2725__S0 (.DIODE(_0873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2718__S0 (.DIODE(_0873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2706__S0 (.DIODE(_0873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2691__S0 (.DIODE(_0873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2629__B_N (.DIODE(_0873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2595__S (.DIODE(_0873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2481__S (.DIODE(_0873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2493__A2 (.DIODE(_0883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2497__A2 (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4131__B (.DIODE(_0903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2514__A3 (.DIODE(_0903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3831__A (.DIODE(_0911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3755__A (.DIODE(_0911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3634__A (.DIODE(_0911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3576__A (.DIODE(_0911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3428__A (.DIODE(_0911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3406__A (.DIODE(_0911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3256__A (.DIODE(_0911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3044__A (.DIODE(_0911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2850__A (.DIODE(_0911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2519__A (.DIODE(_0911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3036__A0 (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3027__A0 (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3018__A0 (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2945__A0 (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2936__A0 (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2906__A0 (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2896__A0 (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2872__A0 (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2842__A0 (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2526__A0 (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3125__A (.DIODE(_0913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3104__A (.DIODE(_0913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3094__A (.DIODE(_0913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3045__A (.DIODE(_0913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3035__A (.DIODE(_0913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3026__A (.DIODE(_0913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2521__A (.DIODE(_0913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3152__A (.DIODE(_0914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3143__A (.DIODE(_0914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3134__A (.DIODE(_0914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3005__A (.DIODE(_0914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2988__A (.DIODE(_0914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2977__A (.DIODE(_0914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2966__A (.DIODE(_0914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2955__A (.DIODE(_0914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2841__A (.DIODE(_0914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2525__A (.DIODE(_0914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4348__A (.DIODE(_0917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4276__A (.DIODE(_0917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3907__A (.DIODE(_0917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3804__A (.DIODE(_0917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3635__A (.DIODE(_0917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3450__A (.DIODE(_0917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3269__A (.DIODE(_0917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2525__B (.DIODE(_0917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2829__B1 (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2809__A1 (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2765__A1 (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2713__A1 (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2689__A1 (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2615__C1 (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2601__C1 (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2590__A1 (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2568__A1 (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2567__C1 (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2824__A (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2813__A (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2807__A1 (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2801__B2 (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2779__A (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2728__A (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2719__A (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2711__A1 (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2594__S (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2530__A (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2795__B2 (.DIODE(_0922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2789__A1 (.DIODE(_0922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2773__A1 (.DIODE(_0922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2751__B2 (.DIODE(_0922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2745__A1 (.DIODE(_0922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2699__B2 (.DIODE(_0922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2693__A1 (.DIODE(_0922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2551__A1 (.DIODE(_0922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2543__A1 (.DIODE(_0922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2542__A1 (.DIODE(_0922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2825__S0 (.DIODE(_0923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2814__S0 (.DIODE(_0923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2787__S0 (.DIODE(_0923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2780__S0 (.DIODE(_0923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2746__S (.DIODE(_0923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2670__S (.DIODE(_0923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2656__S (.DIODE(_0923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2587__S (.DIODE(_0923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2560__S (.DIODE(_0923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2532__A (.DIODE(_0923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2794__S0 (.DIODE(_0924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2786__S0 (.DIODE(_0924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2609__S (.DIODE(_0924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2602__S (.DIODE(_0924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2547__S (.DIODE(_0924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2546__A1 (.DIODE(_0924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2545__B_N (.DIODE(_0924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2544__S0 (.DIODE(_0924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2537__S (.DIODE(_0924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2533__S (.DIODE(_0924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2825__S1 (.DIODE(_0927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2812__S1 (.DIODE(_0927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2810__S1 (.DIODE(_0927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2802__S1 (.DIODE(_0927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2797__A (.DIODE(_0927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2787__S1 (.DIODE(_0927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2780__S1 (.DIODE(_0927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2775__B1 (.DIODE(_0927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2715__B1 (.DIODE(_0927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2536__A (.DIODE(_0927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2794__S1 (.DIODE(_0928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2791__A (.DIODE(_0928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2786__S1 (.DIODE(_0928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2747__A (.DIODE(_0928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2695__A (.DIODE(_0928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2612__A1 (.DIODE(_0928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2605__A1 (.DIODE(_0928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2562__A1 (.DIODE(_0928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2544__S1 (.DIODE(_0928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2538__A (.DIODE(_0928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2820__A1 (.DIODE(_0931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2819__B_N (.DIODE(_0931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2770__S0 (.DIODE(_0931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2766__S0 (.DIODE(_0931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2750__S0 (.DIODE(_0931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2742__S0 (.DIODE(_0931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2698__S0 (.DIODE(_0931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2690__S0 (.DIODE(_0931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2613__S0 (.DIODE(_0931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2541__S0 (.DIODE(_0931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2770__S1 (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2766__S1 (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2750__S1 (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2742__S1 (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2698__S1 (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2690__S1 (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2671__A (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2598__A1 (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2546__B1 (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2541__S1 (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2828__A1 (.DIODE(_0940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2817__A1 (.DIODE(_0940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2793__B1 (.DIODE(_0940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2783__A1 (.DIODE(_0940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2769__A1 (.DIODE(_0940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2649__A1 (.DIODE(_0940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2581__A1 (.DIODE(_0940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2576__A1 (.DIODE(_0940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2570__A (.DIODE(_0940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2549__C1 (.DIODE(_0940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2795__C1 (.DIODE(_0942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2769__C1 (.DIODE(_0942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2751__C1 (.DIODE(_0942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2699__C1 (.DIODE(_0942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2675__C1 (.DIODE(_0942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2649__C1 (.DIODE(_0942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2614__B1 (.DIODE(_0942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2576__C1 (.DIODE(_0942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2566__C1 (.DIODE(_0942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2551__C1 (.DIODE(_0942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2829__A1 (.DIODE(_0944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2818__A1 (.DIODE(_0944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2789__C1 (.DIODE(_0944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2784__A1 (.DIODE(_0944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2773__C1 (.DIODE(_0944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2724__A1 (.DIODE(_0944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2693__C1 (.DIODE(_0944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2601__A1 (.DIODE(_0944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2577__A1 (.DIODE(_0944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2567__A1 (.DIODE(_0944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2792__S (.DIODE(_0945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2790__S (.DIODE(_0945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2715__A1 (.DIODE(_0945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2714__B_N (.DIODE(_0945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2599__S0 (.DIODE(_0945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2578__S0 (.DIODE(_0945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2571__S0 (.DIODE(_0945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2569__S0 (.DIODE(_0945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2555__S0 (.DIODE(_0945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2554__S0 (.DIODE(_0945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2675__B2 (.DIODE(_0948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2669__A1 (.DIODE(_0948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2653__A1 (.DIODE(_0948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2614__A1 (.DIODE(_0948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2608__A1 (.DIODE(_0948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2600__B2 (.DIODE(_0948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2589__A1 (.DIODE(_0948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2572__A (.DIODE(_0948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2566__B2 (.DIODE(_0948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2557__S (.DIODE(_0948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2749__B1 (.DIODE(_0953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2744__A (.DIODE(_0953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2726__A (.DIODE(_0953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2717__C1 (.DIODE(_0953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2692__A (.DIODE(_0953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2673__B1 (.DIODE(_0953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2663__A1 (.DIODE(_0953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2657__C1 (.DIODE(_0953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2617__A (.DIODE(_0953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2562__B1 (.DIODE(_0953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2775__A1 (.DIODE(_0955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2774__B_N (.DIODE(_0955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2674__S0 (.DIODE(_0955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2666__S0 (.DIODE(_0955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2650__S0 (.DIODE(_0955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2646__S0 (.DIODE(_0955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2607__S0 (.DIODE(_0955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2582__S0 (.DIODE(_0955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2573__S0 (.DIODE(_0955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2565__S0 (.DIODE(_0955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2674__S1 (.DIODE(_0956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2666__S1 (.DIODE(_0956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2650__S1 (.DIODE(_0956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2646__S1 (.DIODE(_0956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2613__S1 (.DIODE(_0956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2607__S1 (.DIODE(_0956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2582__S1 (.DIODE(_0956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2578__S1 (.DIODE(_0956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2573__S1 (.DIODE(_0956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2565__S1 (.DIODE(_0956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2638__A1 (.DIODE(_0960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2572__B (.DIODE(_0963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2580__B (.DIODE(_0971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2589__A2 (.DIODE(_0974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2821__S (.DIODE(_0975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2696__S (.DIODE(_0975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2655__A1 (.DIODE(_0975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2654__B_N (.DIODE(_0975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2610__S (.DIODE(_0975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2603__S (.DIODE(_0975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2593__S0 (.DIODE(_0975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2592__S0 (.DIODE(_0975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2586__A1 (.DIODE(_0975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2584__B_N (.DIODE(_0975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2823__S1 (.DIODE(_0977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2800__S1 (.DIODE(_0977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2778__S1 (.DIODE(_0977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2771__S1 (.DIODE(_0977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2729__S1 (.DIODE(_0977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2720__S1 (.DIODE(_0977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2701__A (.DIODE(_0977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2691__S1 (.DIODE(_0977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2655__B1 (.DIODE(_0977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2586__B1 (.DIODE(_0977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2594__A1 (.DIODE(_0985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2598__A2 (.DIODE(_0989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2600__B1 (.DIODE(_0991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2822__C1 (.DIODE(_0996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2811__A (.DIODE(_0996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2788__A (.DIODE(_0996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2777__C1 (.DIODE(_0996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2772__A (.DIODE(_0996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2732__A1 (.DIODE(_0996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2723__A1 (.DIODE(_0996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2697__B1 (.DIODE(_0996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2611__B1 (.DIODE(_0996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2605__B1 (.DIODE(_0996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2617__B (.DIODE(_1008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2621__B (.DIODE(_1012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2623__A2 (.DIODE(_1014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2634__A2 (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4139__B (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2641__A2 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3835__A (.DIODE(_1034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3759__A (.DIODE(_1034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3638__A (.DIODE(_1034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3580__A (.DIODE(_1034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3432__A (.DIODE(_1034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3410__A (.DIODE(_1034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3260__A (.DIODE(_1034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3048__A (.DIODE(_1034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2859__A (.DIODE(_1034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2643__A (.DIODE(_1034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3038__A0 (.DIODE(_1035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3029__A0 (.DIODE(_1035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3020__A0 (.DIODE(_1035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2947__A0 (.DIODE(_1035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2938__A0 (.DIODE(_1035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2908__A0 (.DIODE(_1035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2898__A0 (.DIODE(_1035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2874__A0 (.DIODE(_1035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2844__A0 (.DIODE(_1035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2644__A0 (.DIODE(_1035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2649__A2 (.DIODE(_1037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2653__A2 (.DIODE(_1041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2652__B (.DIODE(_1042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2659__B (.DIODE(_1049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2669__A2 (.DIODE(_1057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2668__B (.DIODE(_1058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2675__B1 (.DIODE(_1065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2693__A2 (.DIODE(_1081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2735__B1 (.DIODE(_1104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2724__A2 (.DIODE(_1108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2724__A3 (.DIODE(_1110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2722__B (.DIODE(_1112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2728__B (.DIODE(_1118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2731__B (.DIODE(_1121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4143__B (.DIODE(_1126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2737__A2 (.DIODE(_1126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3838__A (.DIODE(_1129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3762__A (.DIODE(_1129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3641__A (.DIODE(_1129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3583__A (.DIODE(_1129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3435__A (.DIODE(_1129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3413__A (.DIODE(_1129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3263__A (.DIODE(_1129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3051__A (.DIODE(_1129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2862__A (.DIODE(_1129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2739__A (.DIODE(_1129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3040__A0 (.DIODE(_1130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3031__A0 (.DIODE(_1130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3022__A0 (.DIODE(_1130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2949__A0 (.DIODE(_1130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2940__A0 (.DIODE(_1130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2910__A0 (.DIODE(_1130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2900__A0 (.DIODE(_1130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2876__A0 (.DIODE(_1130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2846__A0 (.DIODE(_1130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2740__A0 (.DIODE(_1130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2745__A2 (.DIODE(_1132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2831__A2 (.DIODE(_1155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2768__B (.DIODE(_1157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2773__A2 (.DIODE(_1160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2784__A2 (.DIODE(_1167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2782__B (.DIODE(_1171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2788__B (.DIODE(_1177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2795__B1 (.DIODE(_1184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2801__B1 (.DIODE(_1190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2813__B (.DIODE(_1202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2817__A2 (.DIODE(_1204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2824__B (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4147__B (.DIODE(_1221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2833__B1 (.DIODE(_1221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3841__A (.DIODE(_1224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3765__A (.DIODE(_1224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3644__A (.DIODE(_1224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3586__A (.DIODE(_1224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3438__A (.DIODE(_1224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3416__A (.DIODE(_1224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3266__A (.DIODE(_1224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3054__A (.DIODE(_1224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2865__A (.DIODE(_1224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2835__A (.DIODE(_1224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3042__A0 (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3033__A0 (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3024__A0 (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2951__A0 (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2942__A0 (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2912__A0 (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2902__A0 (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2878__A0 (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2848__A0 (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2836__A0 (.DIODE(_1225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3832__A (.DIODE(_1229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3656__A (.DIODE(_1229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3558__A (.DIODE(_1229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3429__A (.DIODE(_1229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3379__A (.DIODE(_1229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3247__A (.DIODE(_1229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2944__A (.DIODE(_1229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2841__B (.DIODE(_1229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4358__A0 (.DIODE(_1235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4349__A0 (.DIODE(_1235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4340__A0 (.DIODE(_1235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4331__A0 (.DIODE(_1235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2978__A1 (.DIODE(_1235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2967__A1 (.DIODE(_1235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2956__A1 (.DIODE(_1235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2927__A1 (.DIODE(_1235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2886__A1 (.DIODE(_1235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2857__A1 (.DIODE(_1235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3804__B (.DIODE(_1236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3795__A (.DIODE(_1236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3737__A (.DIODE(_1236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3683__A (.DIODE(_1236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3674__A (.DIODE(_1236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3656__B (.DIODE(_1236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2852__A (.DIODE(_1236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3768__A (.DIODE(_1237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3756__A (.DIODE(_1237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3746__A (.DIODE(_1237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3728__A (.DIODE(_1237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3710__A (.DIODE(_1237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3701__A (.DIODE(_1237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3692__A (.DIODE(_1237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3665__A (.DIODE(_1237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2895__A (.DIODE(_1237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2856__A (.DIODE(_1237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4285__A (.DIODE(_1240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3813__A (.DIODE(_1240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3567__A (.DIODE(_1240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3540__A (.DIODE(_1240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3361__A (.DIODE(_1240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3229__A (.DIODE(_1240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2988__B (.DIODE(_1240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2856__B (.DIODE(_1240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4360__A0 (.DIODE(_1243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4351__A0 (.DIODE(_1243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4342__A0 (.DIODE(_1243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4333__A0 (.DIODE(_1243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2980__A1 (.DIODE(_1243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2969__A1 (.DIODE(_1243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2958__A1 (.DIODE(_1243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2929__A1 (.DIODE(_1243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2888__A1 (.DIODE(_1243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2860__A1 (.DIODE(_1243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4362__A0 (.DIODE(_1245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4353__A0 (.DIODE(_1245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4344__A0 (.DIODE(_1245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4335__A0 (.DIODE(_1245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2982__A1 (.DIODE(_1245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2971__A1 (.DIODE(_1245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2960__A1 (.DIODE(_1245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2931__A1 (.DIODE(_1245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2890__A1 (.DIODE(_1245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2863__A1 (.DIODE(_1245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4364__A0 (.DIODE(_1247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4355__A0 (.DIODE(_1247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4346__A0 (.DIODE(_1247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4337__A0 (.DIODE(_1247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2984__A1 (.DIODE(_1247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2973__A1 (.DIODE(_1247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2962__A1 (.DIODE(_1247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2933__A1 (.DIODE(_1247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2892__A1 (.DIODE(_1247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2866__A1 (.DIODE(_1247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4294__A (.DIODE(_1249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4276__B (.DIODE(_1249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3343__A (.DIODE(_1249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3334__A (.DIODE(_1249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3296__A (.DIODE(_1249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2944__B (.DIODE(_1249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2869__A (.DIODE(_1249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4303__A (.DIODE(_1250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4285__B (.DIODE(_1250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4267__A (.DIODE(_1250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3943__A (.DIODE(_1250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3314__A (.DIODE(_1250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3305__A (.DIODE(_1250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3287__A (.DIODE(_1250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3278__A (.DIODE(_1250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2905__A (.DIODE(_1250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2871__A (.DIODE(_1250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4339__A (.DIODE(_1251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3853__A (.DIODE(_1251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3674__B (.DIODE(_1251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3397__A (.DIODE(_1251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3076__A (.DIODE(_1251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3035__B (.DIODE(_1251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2935__A (.DIODE(_1251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2871__B (.DIODE(_1251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3916__A (.DIODE(_1257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3907__B (.DIODE(_1257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3898__A (.DIODE(_1257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3853__B (.DIODE(_1257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3844__A (.DIODE(_1257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3832__B (.DIODE(_1257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2881__A (.DIODE(_1257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3934__A (.DIODE(_1258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3925__A (.DIODE(_1258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3889__A (.DIODE(_1258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3880__A (.DIODE(_1258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3862__A (.DIODE(_1258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3822__A (.DIODE(_1258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3813__B (.DIODE(_1258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3777__A (.DIODE(_1258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3057__A (.DIODE(_1258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2885__A (.DIODE(_1258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4366__A (.DIODE(_1261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3768__B (.DIODE(_1261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3589__A (.DIODE(_1261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3407__A (.DIODE(_1261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3278__B (.DIODE(_1261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3189__A (.DIODE(_1261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3152__B (.DIODE(_1261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2885__B (.DIODE(_1261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4330__A (.DIODE(_1267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4321__A (.DIODE(_1267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3616__A (.DIODE(_1267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3513__A (.DIODE(_1267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3334__B (.DIODE(_1267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3094__B (.DIODE(_1267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3057__B (.DIODE(_1267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2895__B (.DIODE(_1267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3844__B (.DIODE(_1273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3665__B (.DIODE(_1273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3486__A (.DIODE(_1273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3388__A (.DIODE(_1273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3352__A (.DIODE(_1273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3067__A (.DIODE(_1273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3026__B (.DIODE(_1273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2905__B (.DIODE(_1273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3647__A (.DIODE(_1283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3635__B (.DIODE(_1283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3616__B (.DIODE(_1283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3558__B (.DIODE(_1283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3486__B (.DIODE(_1283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2935__B (.DIODE(_1283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2923__A (.DIODE(_1283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3625__A (.DIODE(_1284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3607__A (.DIODE(_1284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3598__A (.DIODE(_1284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3589__B (.DIODE(_1284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3577__A (.DIODE(_1284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3549__A (.DIODE(_1284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3540__B (.DIODE(_1284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3531__A (.DIODE(_1284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3504__A (.DIODE(_1284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2926__A (.DIODE(_1284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3925__B (.DIODE(_1286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3746__B (.DIODE(_1286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3468__A (.DIODE(_1286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3305__B (.DIODE(_1286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3208__A (.DIODE(_1286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3171__A (.DIODE(_1286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3134__B (.DIODE(_1286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2926__B (.DIODE(_1286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3880__B (.DIODE(_1303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3871__A (.DIODE(_1303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3692__B (.DIODE(_1303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3598__B (.DIODE(_1303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3419__A (.DIODE(_1303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3287__B (.DIODE(_1303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3198__A (.DIODE(_1303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2955__B (.DIODE(_1303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4258__A (.DIODE(_1310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4249__A (.DIODE(_1310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3943__B (.DIODE(_1310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3889__B (.DIODE(_1310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3786__A (.DIODE(_1310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3701__B (.DIODE(_1310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3607__B (.DIODE(_1310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2966__B (.DIODE(_1310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4267__B (.DIODE(_1317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3862__B (.DIODE(_1317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3719__A (.DIODE(_1317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3710__B (.DIODE(_1317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3531__B (.DIODE(_1317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3441__A (.DIODE(_1317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3220__A (.DIODE(_1317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2977__B (.DIODE(_1317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4367__A1 (.DIODE(_1323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4304__A1 (.DIODE(_1323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4286__A1 (.DIODE(_1323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4268__A1 (.DIODE(_1323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4259__A1 (.DIODE(_1323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4250__A1 (.DIODE(_1323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3944__A1 (.DIODE(_1323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3935__A1 (.DIODE(_1323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3207__A (.DIODE(_1323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2987__A (.DIODE(_1323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3199__A1 (.DIODE(_1324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3190__A1 (.DIODE(_1324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3181__A1 (.DIODE(_1324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3172__A1 (.DIODE(_1324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3153__A1 (.DIODE(_1324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3144__A1 (.DIODE(_1324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3135__A1 (.DIODE(_1324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3116__A1 (.DIODE(_1324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3006__A1 (.DIODE(_1324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2989__A1 (.DIODE(_1324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4369__A1 (.DIODE(_1327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4306__A1 (.DIODE(_1327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4288__A1 (.DIODE(_1327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4270__A1 (.DIODE(_1327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4261__A1 (.DIODE(_1327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4252__A1 (.DIODE(_1327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3946__A1 (.DIODE(_1327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3937__A1 (.DIODE(_1327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3211__A (.DIODE(_1327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2992__A (.DIODE(_1327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3201__A1 (.DIODE(_1328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3192__A1 (.DIODE(_1328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3183__A1 (.DIODE(_1328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3174__A1 (.DIODE(_1328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3155__A1 (.DIODE(_1328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3146__A1 (.DIODE(_1328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3137__A1 (.DIODE(_1328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3118__A1 (.DIODE(_1328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3008__A1 (.DIODE(_1328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2993__A1 (.DIODE(_1328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4371__A1 (.DIODE(_1330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4308__A1 (.DIODE(_1330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4290__A1 (.DIODE(_1330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4272__A1 (.DIODE(_1330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4263__A1 (.DIODE(_1330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4254__A1 (.DIODE(_1330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3948__A1 (.DIODE(_1330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3939__A1 (.DIODE(_1330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3214__A (.DIODE(_1330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2996__A (.DIODE(_1330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3203__A1 (.DIODE(_1331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3194__A1 (.DIODE(_1331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3185__A1 (.DIODE(_1331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3176__A1 (.DIODE(_1331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3157__A1 (.DIODE(_1331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3148__A1 (.DIODE(_1331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3139__A1 (.DIODE(_1331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3120__A1 (.DIODE(_1331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3010__A1 (.DIODE(_1331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2997__A1 (.DIODE(_1331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4373__A1 (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4310__A1 (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4292__A1 (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4274__A1 (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4265__A1 (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4256__A1 (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3950__A1 (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3941__A1 (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3217__A (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3000__A (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3205__A1 (.DIODE(_1334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3196__A1 (.DIODE(_1334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3187__A1 (.DIODE(_1334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3178__A1 (.DIODE(_1334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3159__A1 (.DIODE(_1334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3150__A1 (.DIODE(_1334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3141__A1 (.DIODE(_1334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3122__A1 (.DIODE(_1334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3012__A1 (.DIODE(_1334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3001__A1 (.DIODE(_1334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4303__B (.DIODE(_1337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3822__B (.DIODE(_1337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3728__B (.DIODE(_1337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3549__B (.DIODE(_1337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3495__A (.DIODE(_1337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3370__A (.DIODE(_1337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3238__A (.DIODE(_1337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3005__B (.DIODE(_1337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4357__A (.DIODE(_1343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4348__B (.DIODE(_1343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4339__B (.DIODE(_1343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4330__B (.DIODE(_1343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3429__B (.DIODE(_1343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3352__B (.DIODE(_1343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3015__A (.DIODE(_1343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4366__B (.DIODE(_1344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4312__A (.DIODE(_1344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3871__B (.DIODE(_1344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3786__B (.DIODE(_1344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3719__B (.DIODE(_1344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3567__B (.DIODE(_1344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3495__B (.DIODE(_1344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3208__B (.DIODE(_1344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3115__A (.DIODE(_1344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3017__A (.DIODE(_1344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4294__B (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3777__B (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3683__B (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3504__B (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3325__A (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3085__A (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3045__B (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3017__B (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3248__A0 (.DIODE(_1361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3163__A0 (.DIODE(_1361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3126__A0 (.DIODE(_1361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3105__A0 (.DIODE(_1361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3095__A0 (.DIODE(_1361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3086__A0 (.DIODE(_1361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3077__A0 (.DIODE(_1361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3068__A0 (.DIODE(_1361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3058__A0 (.DIODE(_1361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3046__A0 (.DIODE(_1361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3250__A0 (.DIODE(_1364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3165__A0 (.DIODE(_1364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3128__A0 (.DIODE(_1364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3107__A0 (.DIODE(_1364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3097__A0 (.DIODE(_1364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3088__A0 (.DIODE(_1364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3079__A0 (.DIODE(_1364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3070__A0 (.DIODE(_1364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3060__A0 (.DIODE(_1364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3049__A0 (.DIODE(_1364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3252__A0 (.DIODE(_1366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3167__A0 (.DIODE(_1366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3130__A0 (.DIODE(_1366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3109__A0 (.DIODE(_1366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3099__A0 (.DIODE(_1366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3090__A0 (.DIODE(_1366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3081__A0 (.DIODE(_1366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3072__A0 (.DIODE(_1366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3062__A0 (.DIODE(_1366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3052__A0 (.DIODE(_1366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3254__A0 (.DIODE(_1368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3169__A0 (.DIODE(_1368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3132__A0 (.DIODE(_1368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3111__A0 (.DIODE(_1368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3101__A0 (.DIODE(_1368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3092__A0 (.DIODE(_1368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3083__A0 (.DIODE(_1368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3074__A0 (.DIODE(_1368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3064__A0 (.DIODE(_1368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3055__A0 (.DIODE(_1368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4321__B (.DIODE(_1375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3269__B (.DIODE(_1375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3247__B (.DIODE(_1375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3161__A (.DIODE(_1375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3085__B (.DIODE(_1375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3076__B (.DIODE(_1375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3067__B (.DIODE(_1375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4357__B (.DIODE(_1396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3898__B (.DIODE(_1396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3795__B (.DIODE(_1396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3625__B (.DIODE(_1396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3522__A (.DIODE(_1396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3343__B (.DIODE(_1396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3257__B (.DIODE(_1396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3104__B (.DIODE(_1396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3934__B (.DIODE(_1403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3756__B (.DIODE(_1403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3577__B (.DIODE(_1403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3477__A (.DIODE(_1403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3314__B (.DIODE(_1403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3180__B (.DIODE(_1403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3143__B (.DIODE(_1403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3115__B (.DIODE(_1403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4312__B (.DIODE(_1409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3916__B (.DIODE(_1409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3737__B (.DIODE(_1409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3647__B (.DIODE(_1409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3459__A (.DIODE(_1409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3296__B (.DIODE(_1409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3162__B (.DIODE(_1409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3125__B (.DIODE(_1409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4249__B (.DIODE(_1430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3257__A (.DIODE(_1430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3238__B (.DIODE(_1430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3229__B (.DIODE(_1430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3220__B (.DIODE(_1430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3198__B (.DIODE(_1430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3189__B (.DIODE(_1430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3180__A (.DIODE(_1430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3171__B (.DIODE(_1430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3162__A (.DIODE(_1430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3371__A1 (.DIODE(_1456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3362__A1 (.DIODE(_1456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3315__A1 (.DIODE(_1456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3306__A1 (.DIODE(_1456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3288__A1 (.DIODE(_1456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3279__A1 (.DIODE(_1456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3239__A1 (.DIODE(_1456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3230__A1 (.DIODE(_1456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3221__A1 (.DIODE(_1456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3209__A1 (.DIODE(_1456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3373__A1 (.DIODE(_1459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3364__A1 (.DIODE(_1459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3317__A1 (.DIODE(_1459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3308__A1 (.DIODE(_1459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3290__A1 (.DIODE(_1459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3281__A1 (.DIODE(_1459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3241__A1 (.DIODE(_1459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3232__A1 (.DIODE(_1459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3223__A1 (.DIODE(_1459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3212__A1 (.DIODE(_1459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3375__A1 (.DIODE(_1461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3366__A1 (.DIODE(_1461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3319__A1 (.DIODE(_1461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3310__A1 (.DIODE(_1461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3292__A1 (.DIODE(_1461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3283__A1 (.DIODE(_1461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3243__A1 (.DIODE(_1461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3234__A1 (.DIODE(_1461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3225__A1 (.DIODE(_1461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3215__A1 (.DIODE(_1461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3377__A1 (.DIODE(_1463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3368__A1 (.DIODE(_1463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3321__A1 (.DIODE(_1463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3312__A1 (.DIODE(_1463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3294__A1 (.DIODE(_1463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3285__A1 (.DIODE(_1463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3245__A1 (.DIODE(_1463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3236__A1 (.DIODE(_1463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3227__A1 (.DIODE(_1463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3218__A1 (.DIODE(_1463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3398__A0 (.DIODE(_1485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3389__A0 (.DIODE(_1485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3380__A0 (.DIODE(_1485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3353__A0 (.DIODE(_1485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3344__A0 (.DIODE(_1485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3335__A0 (.DIODE(_1485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3326__A0 (.DIODE(_1485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3297__A0 (.DIODE(_1485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3270__A0 (.DIODE(_1485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3258__A0 (.DIODE(_1485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3400__A0 (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3391__A0 (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3382__A0 (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3355__A0 (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3346__A0 (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3337__A0 (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3328__A0 (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3299__A0 (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3272__A0 (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3261__A0 (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3402__A0 (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3393__A0 (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3384__A0 (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3357__A0 (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3348__A0 (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3339__A0 (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3330__A0 (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3301__A0 (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3274__A0 (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3264__A0 (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3404__A0 (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3395__A0 (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3386__A0 (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3359__A0 (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3350__A0 (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3341__A0 (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3332__A0 (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3303__A0 (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3276__A0 (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3267__A0 (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3312__S (.DIODE(_1514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3310__S (.DIODE(_1514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3308__S (.DIODE(_1514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3306__S (.DIODE(_1514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3321__S (.DIODE(_1519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3319__S (.DIODE(_1519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3317__S (.DIODE(_1519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3315__S (.DIODE(_1519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4258__B (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3477__B (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3468__B (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3441__B (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3419__B (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3407__B (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3379__B (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3370__B (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3361__B (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3325__B (.DIODE(_1525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3568__A1 (.DIODE(_1571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3550__A1 (.DIODE(_1571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3541__A1 (.DIODE(_1571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3532__A1 (.DIODE(_1571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3496__A1 (.DIODE(_1571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3478__A1 (.DIODE(_1571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3469__A1 (.DIODE(_1571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3442__A1 (.DIODE(_1571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3420__A1 (.DIODE(_1571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3408__A1 (.DIODE(_1571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3570__A1 (.DIODE(_1574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3552__A1 (.DIODE(_1574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3543__A1 (.DIODE(_1574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3534__A1 (.DIODE(_1574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3498__A1 (.DIODE(_1574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3480__A1 (.DIODE(_1574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3471__A1 (.DIODE(_1574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3444__A1 (.DIODE(_1574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3422__A1 (.DIODE(_1574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3411__A1 (.DIODE(_1574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3572__A1 (.DIODE(_1576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3554__A1 (.DIODE(_1576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3545__A1 (.DIODE(_1576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3536__A1 (.DIODE(_1576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3500__A1 (.DIODE(_1576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3482__A1 (.DIODE(_1576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3473__A1 (.DIODE(_1576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3446__A1 (.DIODE(_1576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3424__A1 (.DIODE(_1576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3414__A1 (.DIODE(_1576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3574__A1 (.DIODE(_1578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3556__A1 (.DIODE(_1578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3547__A1 (.DIODE(_1578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3538__A1 (.DIODE(_1578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3502__A1 (.DIODE(_1578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3484__A1 (.DIODE(_1578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3475__A1 (.DIODE(_1578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3448__A1 (.DIODE(_1578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3426__A1 (.DIODE(_1578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3417__A1 (.DIODE(_1578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3626__A0 (.DIODE(_1585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3617__A0 (.DIODE(_1585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3559__A0 (.DIODE(_1585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3523__A0 (.DIODE(_1585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3514__A0 (.DIODE(_1585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3505__A0 (.DIODE(_1585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3487__A0 (.DIODE(_1585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3460__A0 (.DIODE(_1585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3451__A0 (.DIODE(_1585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3430__A0 (.DIODE(_1585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3628__A0 (.DIODE(_1588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3619__A0 (.DIODE(_1588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3561__A0 (.DIODE(_1588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3525__A0 (.DIODE(_1588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3516__A0 (.DIODE(_1588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3507__A0 (.DIODE(_1588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3489__A0 (.DIODE(_1588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3462__A0 (.DIODE(_1588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3453__A0 (.DIODE(_1588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3433__A0 (.DIODE(_1588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3630__A0 (.DIODE(_1590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3621__A0 (.DIODE(_1590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3563__A0 (.DIODE(_1590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3527__A0 (.DIODE(_1590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3518__A0 (.DIODE(_1590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3509__A0 (.DIODE(_1590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3491__A0 (.DIODE(_1590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3464__A0 (.DIODE(_1590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3455__A0 (.DIODE(_1590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3436__A0 (.DIODE(_1590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3632__A0 (.DIODE(_1592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3623__A0 (.DIODE(_1592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3565__A0 (.DIODE(_1592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3529__A0 (.DIODE(_1592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3520__A0 (.DIODE(_1592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3511__A0 (.DIODE(_1592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3493__A0 (.DIODE(_1592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3466__A0 (.DIODE(_1592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3457__A0 (.DIODE(_1592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3439__A0 (.DIODE(_1592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3457__S (.DIODE(_1599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3455__S (.DIODE(_1599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3453__S (.DIODE(_1599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3451__S (.DIODE(_1599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3520__S (.DIODE(_1634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3518__S (.DIODE(_1634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3516__S (.DIODE(_1634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3514__S (.DIODE(_1634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3529__S (.DIODE(_1639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3527__S (.DIODE(_1639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3525__S (.DIODE(_1639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3523__S (.DIODE(_1639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3747__A1 (.DIODE(_1669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3729__A1 (.DIODE(_1669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3720__A1 (.DIODE(_1669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3711__A1 (.DIODE(_1669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3702__A1 (.DIODE(_1669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3693__A1 (.DIODE(_1669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3608__A1 (.DIODE(_1669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3599__A1 (.DIODE(_1669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3590__A1 (.DIODE(_1669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3578__A1 (.DIODE(_1669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3749__A1 (.DIODE(_1672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3731__A1 (.DIODE(_1672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3722__A1 (.DIODE(_1672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3713__A1 (.DIODE(_1672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3704__A1 (.DIODE(_1672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3695__A1 (.DIODE(_1672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3610__A1 (.DIODE(_1672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3601__A1 (.DIODE(_1672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3592__A1 (.DIODE(_1672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3581__A1 (.DIODE(_1672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3751__A1 (.DIODE(_1674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3733__A1 (.DIODE(_1674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3724__A1 (.DIODE(_1674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3715__A1 (.DIODE(_1674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3706__A1 (.DIODE(_1674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3697__A1 (.DIODE(_1674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3612__A1 (.DIODE(_1674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3603__A1 (.DIODE(_1674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3594__A1 (.DIODE(_1674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3584__A1 (.DIODE(_1674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3753__A1 (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3735__A1 (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3726__A1 (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3717__A1 (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3708__A1 (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3699__A1 (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3614__A1 (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3605__A1 (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3596__A1 (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3587__A1 (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3805__A0 (.DIODE(_1703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3796__A0 (.DIODE(_1703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3778__A0 (.DIODE(_1703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3738__A0 (.DIODE(_1703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3684__A0 (.DIODE(_1703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3675__A0 (.DIODE(_1703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3666__A0 (.DIODE(_1703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3657__A0 (.DIODE(_1703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3648__A0 (.DIODE(_1703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3636__A0 (.DIODE(_1703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3807__A0 (.DIODE(_1706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3798__A0 (.DIODE(_1706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3780__A0 (.DIODE(_1706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3740__A0 (.DIODE(_1706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3686__A0 (.DIODE(_1706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3677__A0 (.DIODE(_1706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3668__A0 (.DIODE(_1706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3659__A0 (.DIODE(_1706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3650__A0 (.DIODE(_1706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3639__A0 (.DIODE(_1706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3809__A0 (.DIODE(_1708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3800__A0 (.DIODE(_1708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3782__A0 (.DIODE(_1708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3742__A0 (.DIODE(_1708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3688__A0 (.DIODE(_1708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3679__A0 (.DIODE(_1708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3670__A0 (.DIODE(_1708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3661__A0 (.DIODE(_1708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3652__A0 (.DIODE(_1708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3642__A0 (.DIODE(_1708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3811__A0 (.DIODE(_1710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3802__A0 (.DIODE(_1710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3784__A0 (.DIODE(_1710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3744__A0 (.DIODE(_1710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3690__A0 (.DIODE(_1710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3681__A0 (.DIODE(_1710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3672__A0 (.DIODE(_1710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3663__A0 (.DIODE(_1710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3654__A0 (.DIODE(_1710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3645__A0 (.DIODE(_1710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3926__A1 (.DIODE(_1772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3890__A1 (.DIODE(_1772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3881__A1 (.DIODE(_1772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3872__A1 (.DIODE(_1772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3863__A1 (.DIODE(_1772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3823__A1 (.DIODE(_1772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3814__A1 (.DIODE(_1772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3787__A1 (.DIODE(_1772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3769__A1 (.DIODE(_1772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3757__A1 (.DIODE(_1772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3766__S (.DIODE(_1773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3763__S (.DIODE(_1773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3760__S (.DIODE(_1773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3757__S (.DIODE(_1773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3928__A1 (.DIODE(_1775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3892__A1 (.DIODE(_1775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3883__A1 (.DIODE(_1775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3874__A1 (.DIODE(_1775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3865__A1 (.DIODE(_1775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3825__A1 (.DIODE(_1775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3816__A1 (.DIODE(_1775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3789__A1 (.DIODE(_1775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3771__A1 (.DIODE(_1775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3760__A1 (.DIODE(_1775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3930__A1 (.DIODE(_1777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3894__A1 (.DIODE(_1777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3885__A1 (.DIODE(_1777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3876__A1 (.DIODE(_1777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3867__A1 (.DIODE(_1777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3827__A1 (.DIODE(_1777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3818__A1 (.DIODE(_1777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3791__A1 (.DIODE(_1777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3773__A1 (.DIODE(_1777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3763__A1 (.DIODE(_1777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3932__A1 (.DIODE(_1779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3896__A1 (.DIODE(_1779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3887__A1 (.DIODE(_1779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3878__A1 (.DIODE(_1779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3869__A1 (.DIODE(_1779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3829__A1 (.DIODE(_1779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3820__A1 (.DIODE(_1779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3793__A1 (.DIODE(_1779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3775__A1 (.DIODE(_1779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3766__A1 (.DIODE(_1779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3820__S (.DIODE(_1806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3818__S (.DIODE(_1806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3816__S (.DIODE(_1806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3814__S (.DIODE(_1806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3829__S (.DIODE(_1811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3827__S (.DIODE(_1811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3825__S (.DIODE(_1811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3823__S (.DIODE(_1811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4322__A0 (.DIODE(_1816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4313__A0 (.DIODE(_1816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4295__A0 (.DIODE(_1816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4277__A0 (.DIODE(_1816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3917__A0 (.DIODE(_1816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3908__A0 (.DIODE(_1816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3899__A0 (.DIODE(_1816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3854__A0 (.DIODE(_1816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3845__A0 (.DIODE(_1816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3833__A0 (.DIODE(_1816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4324__A0 (.DIODE(_1819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4315__A0 (.DIODE(_1819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4297__A0 (.DIODE(_1819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4279__A0 (.DIODE(_1819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3919__A0 (.DIODE(_1819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3910__A0 (.DIODE(_1819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3901__A0 (.DIODE(_1819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3856__A0 (.DIODE(_1819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3847__A0 (.DIODE(_1819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3836__A0 (.DIODE(_1819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4326__A0 (.DIODE(_1821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4317__A0 (.DIODE(_1821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4299__A0 (.DIODE(_1821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4281__A0 (.DIODE(_1821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3921__A0 (.DIODE(_1821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3912__A0 (.DIODE(_1821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3903__A0 (.DIODE(_1821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3858__A0 (.DIODE(_1821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3849__A0 (.DIODE(_1821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3839__A0 (.DIODE(_1821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4328__A0 (.DIODE(_1823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4319__A0 (.DIODE(_1823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4301__A0 (.DIODE(_1823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4283__A0 (.DIODE(_1823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3923__A0 (.DIODE(_1823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3914__A0 (.DIODE(_1823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3905__A0 (.DIODE(_1823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3860__A0 (.DIODE(_1823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3851__A0 (.DIODE(_1823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3842__A0 (.DIODE(_1823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3950__S (.DIODE(_1880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3948__S (.DIODE(_1880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3946__S (.DIODE(_1880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3944__S (.DIODE(_1880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3980__B1 (.DIODE(_1900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4018__C1 (.DIODE(_1901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4015__C1 (.DIODE(_1901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4009__C1 (.DIODE(_1901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4005__C1 (.DIODE(_1901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3999__C1 (.DIODE(_1901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3991__C1 (.DIODE(_1901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3989__C1 (.DIODE(_1901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3984__C1 (.DIODE(_1901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3982__C1 (.DIODE(_1901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3980__C1 (.DIODE(_1901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3982__B1 (.DIODE(_1902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3984__B1 (.DIODE(_1903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4067__C1 (.DIODE(_1931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4064__C1 (.DIODE(_1931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4057__C1 (.DIODE(_1931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4054__C1 (.DIODE(_1931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4051__C1 (.DIODE(_1931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4048__C1 (.DIODE(_1931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4040__C1 (.DIODE(_1931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4037__C1 (.DIODE(_1931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4027__C1 (.DIODE(_1931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4023__C1 (.DIODE(_1931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4227__C1 (.DIODE(_1966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4184__C1 (.DIODE(_1966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4178__C1 (.DIODE(_1966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4172__C1 (.DIODE(_1966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4166__C1 (.DIODE(_1966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4161__C1 (.DIODE(_1966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4084__C1 (.DIODE(_1966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4077__C1 (.DIODE(_1966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4074__C1 (.DIODE(_1966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4071__C1 (.DIODE(_1966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4389__S (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4387__S (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4385__S (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4383__S (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4381__S (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4379__S (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4377__S (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4375__S (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4134__B (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4130__B (.DIODE(_2006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4238__B (.DIODE(_2007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4236__B (.DIODE(_2007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4234__B (.DIODE(_2007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4232__B (.DIODE(_2007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4150__A2 (.DIODE(_2007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4146__A2 (.DIODE(_2007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4142__A2 (.DIODE(_2007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4138__A2 (.DIODE(_2007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4265__S (.DIODE(_2106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4263__S (.DIODE(_2106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4261__S (.DIODE(_2106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4259__S (.DIODE(_2106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4274__S (.DIODE(_2111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4272__S (.DIODE(_2111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4270__S (.DIODE(_2111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4268__S (.DIODE(_2111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3968__A1 (.DIODE(chip_sel_override));
 sky130_fd_sc_hd__diode_2 ANTENNA__2373__A1 (.DIODE(chip_sel_override));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(io_in[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(io_in[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(io_in[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(io_in[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(io_in[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA__4587__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4896__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5009__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4583__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4993__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5008__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5001__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4619__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5000__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4618__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4895__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4614__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4992__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4990__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4893__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4640__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4998__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4639__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4988__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(oram_value[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(oram_value[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(oram_value[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(oram_value[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(oram_value[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(oram_value[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(oram_value[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(oram_value[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(ram_val[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(ram_val[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(ram_val[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(ram_val[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(ram_val[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(ram_val[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(ram_val[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(ram_val[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(ram_val[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(ram_val[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(ram_val[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(ram_val[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(ram_val[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(ram_val[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(ram_val[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(ram_val[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(ram_val[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(ram_val[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(ram_val[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(ram_val[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(ram_val[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(ram_val[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(ram_val[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(ram_val[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(ram_val[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(ram_val[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(ram_val[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(ram_val[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(ram_val[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(ram_val[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(ram_val[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(ram_val[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA__4383__A0 (.DIODE(\tms1x00.PA[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4116__A1 (.DIODE(\tms1x00.PA[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4104__A1 (.DIODE(\tms1x00.PA[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4375__A0 (.DIODE(\tms1x00.PC[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4173__A (.DIODE(\tms1x00.PC[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4172__A1 (.DIODE(\tms1x00.PC[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4169__A1 (.DIODE(\tms1x00.PC[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4093__A1 (.DIODE(\tms1x00.PC[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4377__A0 (.DIODE(\tms1x00.PC[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4179__A (.DIODE(\tms1x00.PC[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4177__A (.DIODE(\tms1x00.PC[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4175__A1 (.DIODE(\tms1x00.PC[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4095__A1 (.DIODE(\tms1x00.PC[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4379__A0 (.DIODE(\tms1x00.PC[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4188__A1 (.DIODE(\tms1x00.PC[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4187__A1 (.DIODE(\tms1x00.PC[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4183__A (.DIODE(\tms1x00.PC[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4181__A1 (.DIODE(\tms1x00.PC[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4097__A1 (.DIODE(\tms1x00.PC[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4381__A0 (.DIODE(\tms1x00.PC[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4189__A1 (.DIODE(\tms1x00.PC[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4186__A1 (.DIODE(\tms1x00.PC[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4099__A1 (.DIODE(\tms1x00.PC[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3446__A0 (.DIODE(\tms1x00.RAM[38][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2651__A2 (.DIODE(\tms1x00.RAM[38][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2938__A1 (.DIODE(\tms1x00.RAM[49][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2633__A1 (.DIODE(\tms1x00.RAM[49][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3628__A1 (.DIODE(\tms1x00.RAM[62][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2627__A2 (.DIODE(\tms1x00.RAM[62][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3630__A1 (.DIODE(\tms1x00.RAM[62][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2660__A2 (.DIODE(\tms1x00.RAM[62][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3632__A1 (.DIODE(\tms1x00.RAM[62][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2825__A2 (.DIODE(\tms1x00.RAM[62][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3617__A1 (.DIODE(\tms1x00.RAM[63][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2500__A3 (.DIODE(\tms1x00.RAM[63][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3619__A1 (.DIODE(\tms1x00.RAM[63][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2627__A3 (.DIODE(\tms1x00.RAM[63][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3621__A1 (.DIODE(\tms1x00.RAM[63][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2660__A3 (.DIODE(\tms1x00.RAM[63][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3935__A0 (.DIODE(\tms1x00.RAM[90][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2408__A2 (.DIODE(\tms1x00.RAM[90][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3937__A0 (.DIODE(\tms1x00.RAM[90][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2565__A2 (.DIODE(\tms1x00.RAM[90][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3939__A0 (.DIODE(\tms1x00.RAM[90][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2698__A2 (.DIODE(\tms1x00.RAM[90][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3941__A0 (.DIODE(\tms1x00.RAM[90][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2750__A2 (.DIODE(\tms1x00.RAM[90][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4197__A0 (.DIODE(\tms1x00.Y[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4136__B2 (.DIODE(\tms1x00.Y[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4010__B (.DIODE(\tms1x00.Y[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4006__A_N (.DIODE(\tms1x00.Y[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4002__B (.DIODE(\tms1x00.Y[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3952__A0 (.DIODE(\tms1x00.Y[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2345__B (.DIODE(\tms1x00.Y[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2323__A0 (.DIODE(\tms1x00.Y[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4205__A0 (.DIODE(\tms1x00.Y[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4140__B2 (.DIODE(\tms1x00.Y[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4010__A (.DIODE(\tms1x00.Y[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4006__B (.DIODE(\tms1x00.Y[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4002__A_N (.DIODE(\tms1x00.Y[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3954__A0 (.DIODE(\tms1x00.Y[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2345__A (.DIODE(\tms1x00.Y[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2326__A0 (.DIODE(\tms1x00.Y[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4213__A0 (.DIODE(\tms1x00.Y[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4045__B (.DIODE(\tms1x00.Y[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4024__A (.DIODE(\tms1x00.Y[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4019__A (.DIODE(\tms1x00.Y[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4011__A (.DIODE(\tms1x00.Y[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2344__A (.DIODE(\tms1x00.Y[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2328__A (.DIODE(\tms1x00.Y[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4222__C (.DIODE(\tms1x00.ins_in[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4082__A (.DIODE(\tms1x00.ins_in[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4059__C (.DIODE(\tms1x00.ins_in[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3974__A0 (.DIODE(\tms1x00.ins_in[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2515__A (.DIODE(\tms1x00.ins_in[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2374__C (.DIODE(\tms1x00.ins_in[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2362__B (.DIODE(\tms1x00.ins_in[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2357__A (.DIODE(\tms1x00.ins_in[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4196__A (.DIODE(\tms1x00.ins_in[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4193__A1 (.DIODE(\tms1x00.ins_in[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4192__A (.DIODE(\tms1x00.ins_in[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4168__A1 (.DIODE(\tms1x00.ins_in[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4137__A1 (.DIODE(\tms1x00.ins_in[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4058__A (.DIODE(\tms1x00.ins_in[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3984__A1 (.DIODE(\tms1x00.ins_in[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2376__B (.DIODE(\tms1x00.ins_in[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2367__A (.DIODE(\tms1x00.ins_in[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2355__A (.DIODE(\tms1x00.ins_in[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4225__A_N (.DIODE(\tms1x00.ins_in[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4196__D_N (.DIODE(\tms1x00.ins_in[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4191__B (.DIODE(\tms1x00.ins_in[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4174__A1 (.DIODE(\tms1x00.ins_in[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4141__A1 (.DIODE(\tms1x00.ins_in[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3985__A0 (.DIODE(\tms1x00.ins_in[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2511__D_N (.DIODE(\tms1x00.ins_in[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2376__A_N (.DIODE(\tms1x00.ins_in[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2354__C (.DIODE(\tms1x00.ins_in[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3956__A1 (.DIODE(\tms1x00.ram_addr_buff[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2882__A (.DIODE(\tms1x00.ram_addr_buff[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2853__C_N (.DIODE(\tms1x00.ram_addr_buff[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2839__A (.DIODE(\tms1x00.ram_addr_buff[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2523__C (.DIODE(\tms1x00.ram_addr_buff[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2329__A1 (.DIODE(\tms1x00.ram_addr_buff[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3958__A1 (.DIODE(\tms1x00.ram_addr_buff[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2882__C_N (.DIODE(\tms1x00.ram_addr_buff[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2853__A (.DIODE(\tms1x00.ram_addr_buff[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2839__B (.DIODE(\tms1x00.ram_addr_buff[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2523__B (.DIODE(\tms1x00.ram_addr_buff[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2333__A1 (.DIODE(\tms1x00.ram_addr_buff[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3966__A (.DIODE(\tms1x00.wb_step ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2317__A (.DIODE(\tms1x00.wb_step ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2311__A1 (.DIODE(\tms1x00.wb_step ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4429__D (.DIODE(valid));
 sky130_fd_sc_hd__diode_2 ANTENNA__2343__B (.DIODE(valid));
 sky130_fd_sc_hd__diode_2 ANTENNA__2308__C (.DIODE(valid));
 sky130_fd_sc_hd__diode_2 ANTENNA__2307__C (.DIODE(valid));
 sky130_fd_sc_hd__diode_2 ANTENNA__2257__C (.DIODE(valid));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_wb_clk_i_A (.DIODE(wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(wb_rst_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(wbs_adr_i[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(wbs_adr_i[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(wbs_adr_i[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(wbs_adr_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(wbs_adr_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(wbs_adr_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(wbs_adr_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(wbs_adr_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(wbs_adr_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(wbs_adr_i[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(wbs_adr_i[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(wbs_cyc_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(wbs_dat_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(wbs_dat_i[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(wbs_dat_i[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(wbs_dat_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input63_A (.DIODE(wbs_dat_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input64_A (.DIODE(wbs_dat_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input65_A (.DIODE(wbs_dat_i[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input66_A (.DIODE(wbs_dat_i[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA__2270__B2 (.DIODE(\wbs_o_buff[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2196__A1 (.DIODE(\wbs_o_buff[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2271__B2 (.DIODE(\wbs_o_buff[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2198__A1 (.DIODE(\wbs_o_buff[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2272__B2 (.DIODE(\wbs_o_buff[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2200__A1 (.DIODE(\wbs_o_buff[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_input67_A (.DIODE(wbs_stb_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_input68_A (.DIODE(wbs_we_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__3971__A1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__3974__A1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__3978__A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__3981__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__2182__A0 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__2203__A0 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__2205__A0 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__2207__A0 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__2211__A0 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__2213__A0 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__2184__A0 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__2224__A0 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__2226__A0 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__2228__A0 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__2230__A0 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__2232__A0 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__2234__A0 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__2236__A0 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__2238__A0 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__2240__A0 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__2186__A0 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__2244__A0 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__2246__A0 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__2188__A0 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__2190__A0 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__2192__A0 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__2194__A0 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__2196__A0 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__2198__A0 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__2200__A0 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__5105__A (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__2308__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__2307__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__2257__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__2246__S (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__2244__S (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__2223__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__2202__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__2181__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__5097__A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__5098__A (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__5099__A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__5100__A (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__5101__A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__5102__A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_output69_A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__4063__A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__2262__A1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_output70_A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__4066__A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__2263__A1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_output71_A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__4069__A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__2264__A1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_output72_A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__4073__A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__2265__A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_output73_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__4076__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__2266__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_output74_A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__4078__A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__2374__B (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__2350__C (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__2267__A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_output75_A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__4159__A2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__3998__B1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__3997__B (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__2374__D_N (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__2350__B (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__2316__B (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__2269__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_output76_A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__4000__A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__3997__A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__2374__A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__2350__A_N (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__2315__A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__2270__A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_output77_A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__2370__B1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__2271__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_output78_A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__4005__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__2272__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_output79_A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__4009__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__2275__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_output80_A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__4015__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__2276__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_output81_A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__4017__B1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__2277__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_output82_A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__4023__A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__2278__A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_output83_A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__4027__A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__2279__A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_output84_A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__4029__B1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__2280__A1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_output85_A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4033__B1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__2281__A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_output86_A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__4036__B1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__2282__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_output87_A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__4039__B1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__2283__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_output88_A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__4041__B1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__2284__A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_output89_A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4047__B1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__2286__A1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_output90_A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__4051__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__2287__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_output91_A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__4054__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__2288__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_output92_A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__4056__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__2289__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_output93_A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__3969__A0 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout148_A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_output94_A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_output95_A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__4375__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_output96_A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__4377__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_output97_A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__4379__A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_output98_A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__4381__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_output101_A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__4387__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_output103_A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__4120__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__4117__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__4112__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__4109__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__4106__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__4001__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3986__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3975__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3972__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_output104_A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_output105_A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_output106_A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_output107_A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_output108_A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_output109_A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_output110_A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_output111_A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_output112_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_output113_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_output114_A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__2257__B (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_output115_A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__4171__A1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__3968__S (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__2364__A (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__2351__A1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__2318__A (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__2312__A2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__2254__S (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__2252__S (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__2250__S (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__2248__S (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__4588__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4580__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4576__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4645__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4679__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4574__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4677__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4641__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4642__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4680__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4638__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4566__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4678__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4986__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4894__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5007__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4643__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4644__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5006__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4999__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4989__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4586__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4991__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4582__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4584__CLK (.DIODE(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4589__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4984__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4985__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5025__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4753__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4757__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4668__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4758__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4754__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5024__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4982__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5022__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4672__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4891__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4578__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5037__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4575__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5036__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4577__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4579__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4983__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4581__CLK (.DIODE(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4585__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4609__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4698__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4705__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4685__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4709__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4716__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4699__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4707__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4708__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4898__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4700__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4732__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4670__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4637__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4667__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4666__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4897__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4706__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4730__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4729__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4682__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4686__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4608__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5041__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5040__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4710__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4714__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5043__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5045__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5042__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4616__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4620__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4602__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4606__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4604__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4603__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5039__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4615__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4713__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4681__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4697__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4617__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4607__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4605__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4621__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4653__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4622__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4731__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4688__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4684__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4712__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4687__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4650__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4646__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4952__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4950__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4954__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4711__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4715__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5038__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4683__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4955__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4965__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4956__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4949__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4913__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5044__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4951__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4656__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4652__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4624__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4912__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4941__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4648__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4647__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4953__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4657__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4654__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4625__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4651__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4975__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4979__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4980__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4968__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4920__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4967__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4914__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4981__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4963__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4958__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4905__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4910__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4628__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4649__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4623__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4909__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4908__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4907__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4974__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4915__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4917__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4978__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4919__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4936__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4918__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4901__CLK (.DIODE(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4674__CLK (.DIODE(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4556__CLK (.DIODE(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4972__CLK (.DIODE(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4595__CLK (.DIODE(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4971__CLK (.DIODE(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4973__CLK (.DIODE(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4960__CLK (.DIODE(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4929__CLK (.DIODE(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4928__CLK (.DIODE(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4931__CLK (.DIODE(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4927__CLK (.DIODE(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4930__CLK (.DIODE(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4976__CLK (.DIODE(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4969__CLK (.DIODE(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4970__CLK (.DIODE(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4977__CLK (.DIODE(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4959__CLK (.DIODE(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4957__CLK (.DIODE(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4391__CLK (.DIODE(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4921__CLK (.DIODE(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4469__CLK (.DIODE(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4494__CLK (.DIODE(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4467__CLK (.DIODE(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4468__CLK (.DIODE(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4636__CLK (.DIODE(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4635__CLK (.DIODE(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4760__CLK (.DIODE(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4759__CLK (.DIODE(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4669__CLK (.DIODE(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4634__CLK (.DIODE(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4466__CLK (.DIODE(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4627__CLK (.DIODE(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4631__CLK (.DIODE(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4655__CLK (.DIODE(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4632__CLK (.DIODE(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4626__CLK (.DIODE(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4630__CLK (.DIODE(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4629__CLK (.DIODE(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4633__CLK (.DIODE(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4902__CLK (.DIODE(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4903__CLK (.DIODE(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4596__CLK (.DIODE(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4900__CLK (.DIODE(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4673__CLK (.DIODE(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4899__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4597__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4601__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4455__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4471__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5017__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4554__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5014__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4456__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4443__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5003__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4472__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4444__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4445__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5011__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5002__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4442__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4457__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5010__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4768__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4764__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4997__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4454__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4470__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4995__CLK (.DIODE(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4846__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4848__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4502__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4856__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4852__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4503__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4498__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4851__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4501__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4847__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4855__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4505__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4436__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4437__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4509__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4500__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4504__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4506__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4435__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4507__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4525__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4520__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4524__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4508__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4884__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4834__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4806__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4774__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4833__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4805__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4880__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4452__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4451__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4473__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4881__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4876__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4879__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4878__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4513__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4434__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4512__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4875__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4850__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4882__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4849__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4853__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4822__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4854__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4823__CLK (.DIODE(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5026__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5030__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4832__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5027__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4762__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4761__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4763__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5013__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4829__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4767__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5012__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5005__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4830__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4453__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4450__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4808__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4765__CLK (.DIODE(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4827__CLK (.DIODE(clknet_leaf_21_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4446__CLK (.DIODE(clknet_leaf_21_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4865__CLK (.DIODE(clknet_leaf_21_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4447__CLK (.DIODE(clknet_leaf_21_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5033__CLK (.DIODE(clknet_leaf_21_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4866__CLK (.DIODE(clknet_leaf_21_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5031__CLK (.DIODE(clknet_leaf_21_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4886__CLK (.DIODE(clknet_leaf_21_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4885__CLK (.DIODE(clknet_leaf_21_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4751__CLK (.DIODE(clknet_leaf_21_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4862__CLK (.DIODE(clknet_leaf_21_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5032__CLK (.DIODE(clknet_leaf_21_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5020__CLK (.DIODE(clknet_leaf_21_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4766__CLK (.DIODE(clknet_leaf_21_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5018__CLK (.DIODE(clknet_leaf_21_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5021__CLK (.DIODE(clknet_leaf_21_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5019__CLK (.DIODE(clknet_leaf_21_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4449__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__5029__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4867__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4448__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4887__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4826__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4814__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4868__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4888__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4825__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4828__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4798__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4797__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4815__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4802__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4440__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4463__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4803__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4749__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4799__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4800__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4789__CLK (.DIODE(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4793__CLK (.DIODE(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4465__CLK (.DIODE(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4747__CLK (.DIODE(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4441__CLK (.DIODE(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4801__CLK (.DIODE(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4804__CLK (.DIODE(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4791__CLK (.DIODE(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4795__CLK (.DIODE(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4811__CLK (.DIODE(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4787__CLK (.DIODE(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4813__CLK (.DIODE(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4810__CLK (.DIODE(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4817__CLK (.DIODE(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4785__CLK (.DIODE(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4794__CLK (.DIODE(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4788__CLK (.DIODE(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4790__CLK (.DIODE(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4820__CLK (.DIODE(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4809__CLK (.DIODE(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4812__CLK (.DIODE(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4424__CLK (.DIODE(clknet_leaf_26_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4419__CLK (.DIODE(clknet_leaf_26_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4418__CLK (.DIODE(clknet_leaf_26_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4414__CLK (.DIODE(clknet_leaf_26_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4412__CLK (.DIODE(clknet_leaf_26_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4745__CLK (.DIODE(clknet_leaf_26_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4741__CLK (.DIODE(clknet_leaf_26_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4738__CLK (.DIODE(clknet_leaf_26_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4740__CLK (.DIODE(clknet_leaf_26_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4742__CLK (.DIODE(clknet_leaf_26_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4748__CLK (.DIODE(clknet_leaf_26_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4744__CLK (.DIODE(clknet_leaf_26_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4423__CLK (.DIODE(clknet_leaf_26_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4425__CLK (.DIODE(clknet_leaf_26_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4752__CLK (.DIODE(clknet_leaf_28_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4750__CLK (.DIODE(clknet_leaf_28_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4439__CLK (.DIODE(clknet_leaf_28_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4722__CLK (.DIODE(clknet_leaf_28_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4409__CLK (.DIODE(clknet_leaf_28_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4413__CLK (.DIODE(clknet_leaf_28_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4734__CLK (.DIODE(clknet_leaf_28_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4438__CLK (.DIODE(clknet_leaf_28_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4724__CLK (.DIODE(clknet_leaf_28_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4743__CLK (.DIODE(clknet_leaf_28_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4464__CLK (.DIODE(clknet_leaf_28_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4462__CLK (.DIODE(clknet_leaf_28_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4726__CLK (.DIODE(clknet_leaf_28_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4725__CLK (.DIODE(clknet_leaf_28_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4739__CLK (.DIODE(clknet_leaf_28_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4721__CLK (.DIODE(clknet_leaf_28_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4737__CLK (.DIODE(clknet_leaf_28_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4735__CLK (.DIODE(clknet_leaf_28_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4703__CLK (.DIODE(clknet_leaf_28_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4736__CLK (.DIODE(clknet_leaf_28_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4704__CLK (.DIODE(clknet_leaf_28_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4406__CLK (.DIODE(clknet_leaf_28_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4408__CLK (.DIODE(clknet_leaf_28_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4410__CLK (.DIODE(clknet_leaf_28_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4664__CLK (.DIODE(clknet_leaf_28_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4476__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4695__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4660__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4691__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4490__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4477__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4549__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4474__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4544__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4552__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4550__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4542__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4547__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4548__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4546__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4558__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4570__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4543__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4545__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4551__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4568__CLK (.DIODE(clknet_leaf_32_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4460__CLK (.DIODE(clknet_leaf_32_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4573__CLK (.DIODE(clknet_leaf_32_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4689__CLK (.DIODE(clknet_leaf_32_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4429__CLK (.DIODE(clknet_leaf_32_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4428__CLK (.DIODE(clknet_leaf_32_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4420__CLK (.DIODE(clknet_leaf_32_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4692__CLK (.DIODE(clknet_leaf_32_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4662__CLK (.DIODE(clknet_leaf_32_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4658__CLK (.DIODE(clknet_leaf_32_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4693__CLK (.DIODE(clknet_leaf_32_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4572__CLK (.DIODE(clknet_leaf_32_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4694__CLK (.DIODE(clknet_leaf_32_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4659__CLK (.DIODE(clknet_leaf_32_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4696__CLK (.DIODE(clknet_leaf_32_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_805 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_890 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_618 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_535 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_718 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_787 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_852 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_842 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_939 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_910 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_932 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_703 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_756 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_859 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_872 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_788 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_831 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_857 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_848 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_855 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_879 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_690 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_911 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_702 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_947 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_819 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_802 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_815 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_847 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_948 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_834 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_901 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_758 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_935 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_918 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_947 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_947 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_759 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_824 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_860 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_908 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_947 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_415 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_826 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_870 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_947 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_887 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_948 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_594 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_947 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_415 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_746 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_824 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_846 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_928 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_504 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_721 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_786 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_859 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_848 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_876 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_848 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_947 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_848 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_845 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_886 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_534 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_583 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_648 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_836 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_308 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_644 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_721 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_415 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_534 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_859 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_935 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_896 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_899 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_820 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_663 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_863 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_550 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_679 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_885 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_875 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_928 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_940 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_832 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_880 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_945 ();
 assign io_oeb[0] = net190;
 assign io_oeb[10] = net149;
 assign io_oeb[11] = net150;
 assign io_oeb[12] = net151;
 assign io_oeb[13] = net152;
 assign io_oeb[14] = net153;
 assign io_oeb[15] = net154;
 assign io_oeb[16] = net155;
 assign io_oeb[17] = net156;
 assign io_oeb[18] = net157;
 assign io_oeb[19] = net158;
 assign io_oeb[1] = net191;
 assign io_oeb[20] = net159;
 assign io_oeb[21] = net160;
 assign io_oeb[22] = net161;
 assign io_oeb[23] = net162;
 assign io_oeb[24] = net163;
 assign io_oeb[25] = net164;
 assign io_oeb[26] = net165;
 assign io_oeb[27] = net166;
 assign io_oeb[28] = net167;
 assign io_oeb[29] = net168;
 assign io_oeb[2] = net192;
 assign io_oeb[30] = net169;
 assign io_oeb[31] = net170;
 assign io_oeb[32] = net171;
 assign io_oeb[33] = net172;
 assign io_oeb[34] = net173;
 assign io_oeb[35] = net174;
 assign io_oeb[36] = net175;
 assign io_oeb[37] = net176;
 assign io_oeb[3] = net193;
 assign io_oeb[4] = net194;
 assign io_oeb[5] = net195;
 assign io_oeb[6] = net196;
 assign io_oeb[7] = net197;
 assign io_oeb[8] = net198;
 assign io_oeb[9] = net199;
 assign io_out[0] = net177;
 assign io_out[1] = net178;
 assign io_out[2] = net179;
 assign io_out[34] = net187;
 assign io_out[35] = net188;
 assign io_out[3] = net180;
 assign io_out[4] = net181;
 assign io_out[5] = net182;
 assign io_out[6] = net183;
 assign io_out[7] = net184;
 assign io_out[8] = net185;
 assign io_out[9] = net186;
 assign oram_addr[8] = net189;
endmodule

