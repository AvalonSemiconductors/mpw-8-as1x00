// This is the unpowered netlist.
module wrapped_tms1x00 (ram_we,
    rom_csb,
    wb_clk_i,
    wb_rom_csb,
    wb_rom_web,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    io_in,
    io_oeb,
    io_out,
    irq,
    ram_addr,
    ram_val_in,
    ram_val_out,
    rom_addr,
    rom_value,
    wb_rom_adrb,
    wb_rom_val,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o);
 output ram_we;
 output rom_csb;
 input wb_clk_i;
 output wb_rom_csb;
 output wb_rom_web;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 output [2:0] irq;
 output [6:0] ram_addr;
 input [3:0] ram_val_in;
 output [3:0] ram_val_out;
 output [8:0] rom_addr;
 input [31:0] rom_value;
 output [8:0] wb_rom_adrb;
 input [31:0] wb_rom_val;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;

 wire net1123;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1124;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1125;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1118;
 wire net1119;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1120;
 wire net1121;
 wire net1122;
 wire \K_override[0] ;
 wire \K_override[1] ;
 wire \K_override[2] ;
 wire \K_override[3] ;
 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire chip_sel_override;
 wire clknet_0_wb_clk_i;
 wire clknet_3_0_0_wb_clk_i;
 wire clknet_3_1_0_wb_clk_i;
 wire clknet_3_2_0_wb_clk_i;
 wire clknet_3_3_0_wb_clk_i;
 wire clknet_3_4_0_wb_clk_i;
 wire clknet_3_5_0_wb_clk_i;
 wire clknet_3_6_0_wb_clk_i;
 wire clknet_3_7_0_wb_clk_i;
 wire clknet_4_0__leaf_wb_clk_i;
 wire clknet_4_10__leaf_wb_clk_i;
 wire clknet_4_11__leaf_wb_clk_i;
 wire clknet_4_12__leaf_wb_clk_i;
 wire clknet_4_13__leaf_wb_clk_i;
 wire clknet_4_14__leaf_wb_clk_i;
 wire clknet_4_15__leaf_wb_clk_i;
 wire clknet_4_1__leaf_wb_clk_i;
 wire clknet_4_2__leaf_wb_clk_i;
 wire clknet_4_3__leaf_wb_clk_i;
 wire clknet_4_4__leaf_wb_clk_i;
 wire clknet_4_5__leaf_wb_clk_i;
 wire clknet_4_6__leaf_wb_clk_i;
 wire clknet_4_7__leaf_wb_clk_i;
 wire clknet_4_8__leaf_wb_clk_i;
 wire clknet_4_9__leaf_wb_clk_i;
 wire clknet_leaf_0_wb_clk_i;
 wire clknet_leaf_100_wb_clk_i;
 wire clknet_leaf_101_wb_clk_i;
 wire clknet_leaf_102_wb_clk_i;
 wire clknet_leaf_103_wb_clk_i;
 wire clknet_leaf_104_wb_clk_i;
 wire clknet_leaf_105_wb_clk_i;
 wire clknet_leaf_106_wb_clk_i;
 wire clknet_leaf_107_wb_clk_i;
 wire clknet_leaf_108_wb_clk_i;
 wire clknet_leaf_109_wb_clk_i;
 wire clknet_leaf_10_wb_clk_i;
 wire clknet_leaf_110_wb_clk_i;
 wire clknet_leaf_111_wb_clk_i;
 wire clknet_leaf_112_wb_clk_i;
 wire clknet_leaf_113_wb_clk_i;
 wire clknet_leaf_114_wb_clk_i;
 wire clknet_leaf_115_wb_clk_i;
 wire clknet_leaf_116_wb_clk_i;
 wire clknet_leaf_117_wb_clk_i;
 wire clknet_leaf_118_wb_clk_i;
 wire clknet_leaf_119_wb_clk_i;
 wire clknet_leaf_11_wb_clk_i;
 wire clknet_leaf_120_wb_clk_i;
 wire clknet_leaf_121_wb_clk_i;
 wire clknet_leaf_122_wb_clk_i;
 wire clknet_leaf_123_wb_clk_i;
 wire clknet_leaf_124_wb_clk_i;
 wire clknet_leaf_125_wb_clk_i;
 wire clknet_leaf_126_wb_clk_i;
 wire clknet_leaf_127_wb_clk_i;
 wire clknet_leaf_128_wb_clk_i;
 wire clknet_leaf_129_wb_clk_i;
 wire clknet_leaf_12_wb_clk_i;
 wire clknet_leaf_130_wb_clk_i;
 wire clknet_leaf_131_wb_clk_i;
 wire clknet_leaf_132_wb_clk_i;
 wire clknet_leaf_133_wb_clk_i;
 wire clknet_leaf_134_wb_clk_i;
 wire clknet_leaf_135_wb_clk_i;
 wire clknet_leaf_136_wb_clk_i;
 wire clknet_leaf_137_wb_clk_i;
 wire clknet_leaf_138_wb_clk_i;
 wire clknet_leaf_139_wb_clk_i;
 wire clknet_leaf_13_wb_clk_i;
 wire clknet_leaf_140_wb_clk_i;
 wire clknet_leaf_141_wb_clk_i;
 wire clknet_leaf_142_wb_clk_i;
 wire clknet_leaf_143_wb_clk_i;
 wire clknet_leaf_14_wb_clk_i;
 wire clknet_leaf_15_wb_clk_i;
 wire clknet_leaf_16_wb_clk_i;
 wire clknet_leaf_17_wb_clk_i;
 wire clknet_leaf_18_wb_clk_i;
 wire clknet_leaf_19_wb_clk_i;
 wire clknet_leaf_1_wb_clk_i;
 wire clknet_leaf_20_wb_clk_i;
 wire clknet_leaf_21_wb_clk_i;
 wire clknet_leaf_22_wb_clk_i;
 wire clknet_leaf_23_wb_clk_i;
 wire clknet_leaf_24_wb_clk_i;
 wire clknet_leaf_25_wb_clk_i;
 wire clknet_leaf_26_wb_clk_i;
 wire clknet_leaf_27_wb_clk_i;
 wire clknet_leaf_28_wb_clk_i;
 wire clknet_leaf_29_wb_clk_i;
 wire clknet_leaf_2_wb_clk_i;
 wire clknet_leaf_30_wb_clk_i;
 wire clknet_leaf_31_wb_clk_i;
 wire clknet_leaf_32_wb_clk_i;
 wire clknet_leaf_33_wb_clk_i;
 wire clknet_leaf_34_wb_clk_i;
 wire clknet_leaf_35_wb_clk_i;
 wire clknet_leaf_36_wb_clk_i;
 wire clknet_leaf_37_wb_clk_i;
 wire clknet_leaf_38_wb_clk_i;
 wire clknet_leaf_39_wb_clk_i;
 wire clknet_leaf_3_wb_clk_i;
 wire clknet_leaf_40_wb_clk_i;
 wire clknet_leaf_41_wb_clk_i;
 wire clknet_leaf_42_wb_clk_i;
 wire clknet_leaf_43_wb_clk_i;
 wire clknet_leaf_44_wb_clk_i;
 wire clknet_leaf_45_wb_clk_i;
 wire clknet_leaf_46_wb_clk_i;
 wire clknet_leaf_47_wb_clk_i;
 wire clknet_leaf_48_wb_clk_i;
 wire clknet_leaf_49_wb_clk_i;
 wire clknet_leaf_4_wb_clk_i;
 wire clknet_leaf_50_wb_clk_i;
 wire clknet_leaf_51_wb_clk_i;
 wire clknet_leaf_52_wb_clk_i;
 wire clknet_leaf_53_wb_clk_i;
 wire clknet_leaf_54_wb_clk_i;
 wire clknet_leaf_55_wb_clk_i;
 wire clknet_leaf_56_wb_clk_i;
 wire clknet_leaf_57_wb_clk_i;
 wire clknet_leaf_58_wb_clk_i;
 wire clknet_leaf_59_wb_clk_i;
 wire clknet_leaf_5_wb_clk_i;
 wire clknet_leaf_60_wb_clk_i;
 wire clknet_leaf_61_wb_clk_i;
 wire clknet_leaf_62_wb_clk_i;
 wire clknet_leaf_63_wb_clk_i;
 wire clknet_leaf_64_wb_clk_i;
 wire clknet_leaf_65_wb_clk_i;
 wire clknet_leaf_66_wb_clk_i;
 wire clknet_leaf_67_wb_clk_i;
 wire clknet_leaf_68_wb_clk_i;
 wire clknet_leaf_69_wb_clk_i;
 wire clknet_leaf_6_wb_clk_i;
 wire clknet_leaf_70_wb_clk_i;
 wire clknet_leaf_71_wb_clk_i;
 wire clknet_leaf_72_wb_clk_i;
 wire clknet_leaf_73_wb_clk_i;
 wire clknet_leaf_74_wb_clk_i;
 wire clknet_leaf_75_wb_clk_i;
 wire clknet_leaf_76_wb_clk_i;
 wire clknet_leaf_77_wb_clk_i;
 wire clknet_leaf_78_wb_clk_i;
 wire clknet_leaf_79_wb_clk_i;
 wire clknet_leaf_7_wb_clk_i;
 wire clknet_leaf_80_wb_clk_i;
 wire clknet_leaf_81_wb_clk_i;
 wire clknet_leaf_82_wb_clk_i;
 wire clknet_leaf_83_wb_clk_i;
 wire clknet_leaf_84_wb_clk_i;
 wire clknet_leaf_85_wb_clk_i;
 wire clknet_leaf_86_wb_clk_i;
 wire clknet_leaf_87_wb_clk_i;
 wire clknet_leaf_88_wb_clk_i;
 wire clknet_leaf_89_wb_clk_i;
 wire clknet_leaf_8_wb_clk_i;
 wire clknet_leaf_90_wb_clk_i;
 wire clknet_leaf_91_wb_clk_i;
 wire clknet_leaf_92_wb_clk_i;
 wire clknet_leaf_93_wb_clk_i;
 wire clknet_leaf_94_wb_clk_i;
 wire clknet_leaf_95_wb_clk_i;
 wire clknet_leaf_96_wb_clk_i;
 wire clknet_leaf_97_wb_clk_i;
 wire clknet_leaf_98_wb_clk_i;
 wire clknet_leaf_99_wb_clk_i;
 wire clknet_leaf_9_wb_clk_i;
 wire feedback_delay;
 wire net1;
 wire net10;
 wire net100;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net101;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net102;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net103;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net104;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net105;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net106;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net107;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net1133;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net87;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net88;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net89;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net9;
 wire net90;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net91;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net92;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net93;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net94;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net95;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net96;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net97;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net98;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net99;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire \tms1x00.A[0] ;
 wire \tms1x00.A[1] ;
 wire \tms1x00.A[2] ;
 wire \tms1x00.A[3] ;
 wire \tms1x00.B[0] ;
 wire \tms1x00.B[1] ;
 wire \tms1x00.CA ;
 wire \tms1x00.CB ;
 wire \tms1x00.CL ;
 wire \tms1x00.CS ;
 wire \tms1x00.K_in[0] ;
 wire \tms1x00.K_in[1] ;
 wire \tms1x00.K_in[2] ;
 wire \tms1x00.K_in[3] ;
 wire \tms1x00.K_latch[0] ;
 wire \tms1x00.K_latch[1] ;
 wire \tms1x00.K_latch[2] ;
 wire \tms1x00.K_latch[3] ;
 wire \tms1x00.N[0] ;
 wire \tms1x00.N[1] ;
 wire \tms1x00.N[2] ;
 wire \tms1x00.N[3] ;
 wire \tms1x00.O_latch[0] ;
 wire \tms1x00.O_latch[1] ;
 wire \tms1x00.O_latch[2] ;
 wire \tms1x00.O_latch[3] ;
 wire \tms1x00.O_latch[4] ;
 wire \tms1x00.O_pla_ands[0][0] ;
 wire \tms1x00.O_pla_ands[0][1] ;
 wire \tms1x00.O_pla_ands[0][2] ;
 wire \tms1x00.O_pla_ands[0][3] ;
 wire \tms1x00.O_pla_ands[0][4] ;
 wire \tms1x00.O_pla_ands[0][5] ;
 wire \tms1x00.O_pla_ands[0][6] ;
 wire \tms1x00.O_pla_ands[0][7] ;
 wire \tms1x00.O_pla_ands[0][8] ;
 wire \tms1x00.O_pla_ands[0][9] ;
 wire \tms1x00.O_pla_ands[10][0] ;
 wire \tms1x00.O_pla_ands[10][1] ;
 wire \tms1x00.O_pla_ands[10][2] ;
 wire \tms1x00.O_pla_ands[10][3] ;
 wire \tms1x00.O_pla_ands[10][4] ;
 wire \tms1x00.O_pla_ands[10][5] ;
 wire \tms1x00.O_pla_ands[10][6] ;
 wire \tms1x00.O_pla_ands[10][7] ;
 wire \tms1x00.O_pla_ands[10][8] ;
 wire \tms1x00.O_pla_ands[10][9] ;
 wire \tms1x00.O_pla_ands[11][0] ;
 wire \tms1x00.O_pla_ands[11][1] ;
 wire \tms1x00.O_pla_ands[11][2] ;
 wire \tms1x00.O_pla_ands[11][3] ;
 wire \tms1x00.O_pla_ands[11][4] ;
 wire \tms1x00.O_pla_ands[11][5] ;
 wire \tms1x00.O_pla_ands[11][6] ;
 wire \tms1x00.O_pla_ands[11][7] ;
 wire \tms1x00.O_pla_ands[11][8] ;
 wire \tms1x00.O_pla_ands[11][9] ;
 wire \tms1x00.O_pla_ands[12][0] ;
 wire \tms1x00.O_pla_ands[12][1] ;
 wire \tms1x00.O_pla_ands[12][2] ;
 wire \tms1x00.O_pla_ands[12][3] ;
 wire \tms1x00.O_pla_ands[12][4] ;
 wire \tms1x00.O_pla_ands[12][5] ;
 wire \tms1x00.O_pla_ands[12][6] ;
 wire \tms1x00.O_pla_ands[12][7] ;
 wire \tms1x00.O_pla_ands[12][8] ;
 wire \tms1x00.O_pla_ands[12][9] ;
 wire \tms1x00.O_pla_ands[13][0] ;
 wire \tms1x00.O_pla_ands[13][1] ;
 wire \tms1x00.O_pla_ands[13][2] ;
 wire \tms1x00.O_pla_ands[13][3] ;
 wire \tms1x00.O_pla_ands[13][4] ;
 wire \tms1x00.O_pla_ands[13][5] ;
 wire \tms1x00.O_pla_ands[13][6] ;
 wire \tms1x00.O_pla_ands[13][7] ;
 wire \tms1x00.O_pla_ands[13][8] ;
 wire \tms1x00.O_pla_ands[13][9] ;
 wire \tms1x00.O_pla_ands[14][0] ;
 wire \tms1x00.O_pla_ands[14][1] ;
 wire \tms1x00.O_pla_ands[14][2] ;
 wire \tms1x00.O_pla_ands[14][3] ;
 wire \tms1x00.O_pla_ands[14][4] ;
 wire \tms1x00.O_pla_ands[14][5] ;
 wire \tms1x00.O_pla_ands[14][6] ;
 wire \tms1x00.O_pla_ands[14][7] ;
 wire \tms1x00.O_pla_ands[14][8] ;
 wire \tms1x00.O_pla_ands[14][9] ;
 wire \tms1x00.O_pla_ands[15][0] ;
 wire \tms1x00.O_pla_ands[15][1] ;
 wire \tms1x00.O_pla_ands[15][2] ;
 wire \tms1x00.O_pla_ands[15][3] ;
 wire \tms1x00.O_pla_ands[15][4] ;
 wire \tms1x00.O_pla_ands[15][5] ;
 wire \tms1x00.O_pla_ands[15][6] ;
 wire \tms1x00.O_pla_ands[15][7] ;
 wire \tms1x00.O_pla_ands[15][8] ;
 wire \tms1x00.O_pla_ands[15][9] ;
 wire \tms1x00.O_pla_ands[16][0] ;
 wire \tms1x00.O_pla_ands[16][1] ;
 wire \tms1x00.O_pla_ands[16][2] ;
 wire \tms1x00.O_pla_ands[16][3] ;
 wire \tms1x00.O_pla_ands[16][4] ;
 wire \tms1x00.O_pla_ands[16][5] ;
 wire \tms1x00.O_pla_ands[16][6] ;
 wire \tms1x00.O_pla_ands[16][7] ;
 wire \tms1x00.O_pla_ands[16][8] ;
 wire \tms1x00.O_pla_ands[16][9] ;
 wire \tms1x00.O_pla_ands[17][0] ;
 wire \tms1x00.O_pla_ands[17][1] ;
 wire \tms1x00.O_pla_ands[17][2] ;
 wire \tms1x00.O_pla_ands[17][3] ;
 wire \tms1x00.O_pla_ands[17][4] ;
 wire \tms1x00.O_pla_ands[17][5] ;
 wire \tms1x00.O_pla_ands[17][6] ;
 wire \tms1x00.O_pla_ands[17][7] ;
 wire \tms1x00.O_pla_ands[17][8] ;
 wire \tms1x00.O_pla_ands[17][9] ;
 wire \tms1x00.O_pla_ands[18][0] ;
 wire \tms1x00.O_pla_ands[18][1] ;
 wire \tms1x00.O_pla_ands[18][2] ;
 wire \tms1x00.O_pla_ands[18][3] ;
 wire \tms1x00.O_pla_ands[18][4] ;
 wire \tms1x00.O_pla_ands[18][5] ;
 wire \tms1x00.O_pla_ands[18][6] ;
 wire \tms1x00.O_pla_ands[18][7] ;
 wire \tms1x00.O_pla_ands[18][8] ;
 wire \tms1x00.O_pla_ands[18][9] ;
 wire \tms1x00.O_pla_ands[19][0] ;
 wire \tms1x00.O_pla_ands[19][1] ;
 wire \tms1x00.O_pla_ands[19][2] ;
 wire \tms1x00.O_pla_ands[19][3] ;
 wire \tms1x00.O_pla_ands[19][4] ;
 wire \tms1x00.O_pla_ands[19][5] ;
 wire \tms1x00.O_pla_ands[19][6] ;
 wire \tms1x00.O_pla_ands[19][7] ;
 wire \tms1x00.O_pla_ands[19][8] ;
 wire \tms1x00.O_pla_ands[19][9] ;
 wire \tms1x00.O_pla_ands[1][0] ;
 wire \tms1x00.O_pla_ands[1][1] ;
 wire \tms1x00.O_pla_ands[1][2] ;
 wire \tms1x00.O_pla_ands[1][3] ;
 wire \tms1x00.O_pla_ands[1][4] ;
 wire \tms1x00.O_pla_ands[1][5] ;
 wire \tms1x00.O_pla_ands[1][6] ;
 wire \tms1x00.O_pla_ands[1][7] ;
 wire \tms1x00.O_pla_ands[1][8] ;
 wire \tms1x00.O_pla_ands[1][9] ;
 wire \tms1x00.O_pla_ands[20][0] ;
 wire \tms1x00.O_pla_ands[20][1] ;
 wire \tms1x00.O_pla_ands[20][2] ;
 wire \tms1x00.O_pla_ands[20][3] ;
 wire \tms1x00.O_pla_ands[20][4] ;
 wire \tms1x00.O_pla_ands[20][5] ;
 wire \tms1x00.O_pla_ands[20][6] ;
 wire \tms1x00.O_pla_ands[20][7] ;
 wire \tms1x00.O_pla_ands[20][8] ;
 wire \tms1x00.O_pla_ands[20][9] ;
 wire \tms1x00.O_pla_ands[21][0] ;
 wire \tms1x00.O_pla_ands[21][1] ;
 wire \tms1x00.O_pla_ands[21][2] ;
 wire \tms1x00.O_pla_ands[21][3] ;
 wire \tms1x00.O_pla_ands[21][4] ;
 wire \tms1x00.O_pla_ands[21][5] ;
 wire \tms1x00.O_pla_ands[21][6] ;
 wire \tms1x00.O_pla_ands[21][7] ;
 wire \tms1x00.O_pla_ands[21][8] ;
 wire \tms1x00.O_pla_ands[21][9] ;
 wire \tms1x00.O_pla_ands[22][0] ;
 wire \tms1x00.O_pla_ands[22][1] ;
 wire \tms1x00.O_pla_ands[22][2] ;
 wire \tms1x00.O_pla_ands[22][3] ;
 wire \tms1x00.O_pla_ands[22][4] ;
 wire \tms1x00.O_pla_ands[22][5] ;
 wire \tms1x00.O_pla_ands[22][6] ;
 wire \tms1x00.O_pla_ands[22][7] ;
 wire \tms1x00.O_pla_ands[22][8] ;
 wire \tms1x00.O_pla_ands[22][9] ;
 wire \tms1x00.O_pla_ands[23][0] ;
 wire \tms1x00.O_pla_ands[23][1] ;
 wire \tms1x00.O_pla_ands[23][2] ;
 wire \tms1x00.O_pla_ands[23][3] ;
 wire \tms1x00.O_pla_ands[23][4] ;
 wire \tms1x00.O_pla_ands[23][5] ;
 wire \tms1x00.O_pla_ands[23][6] ;
 wire \tms1x00.O_pla_ands[23][7] ;
 wire \tms1x00.O_pla_ands[23][8] ;
 wire \tms1x00.O_pla_ands[23][9] ;
 wire \tms1x00.O_pla_ands[24][0] ;
 wire \tms1x00.O_pla_ands[24][1] ;
 wire \tms1x00.O_pla_ands[24][2] ;
 wire \tms1x00.O_pla_ands[24][3] ;
 wire \tms1x00.O_pla_ands[24][4] ;
 wire \tms1x00.O_pla_ands[24][5] ;
 wire \tms1x00.O_pla_ands[24][6] ;
 wire \tms1x00.O_pla_ands[24][7] ;
 wire \tms1x00.O_pla_ands[24][8] ;
 wire \tms1x00.O_pla_ands[24][9] ;
 wire \tms1x00.O_pla_ands[25][0] ;
 wire \tms1x00.O_pla_ands[25][1] ;
 wire \tms1x00.O_pla_ands[25][2] ;
 wire \tms1x00.O_pla_ands[25][3] ;
 wire \tms1x00.O_pla_ands[25][4] ;
 wire \tms1x00.O_pla_ands[25][5] ;
 wire \tms1x00.O_pla_ands[25][6] ;
 wire \tms1x00.O_pla_ands[25][7] ;
 wire \tms1x00.O_pla_ands[25][8] ;
 wire \tms1x00.O_pla_ands[25][9] ;
 wire \tms1x00.O_pla_ands[26][0] ;
 wire \tms1x00.O_pla_ands[26][1] ;
 wire \tms1x00.O_pla_ands[26][2] ;
 wire \tms1x00.O_pla_ands[26][3] ;
 wire \tms1x00.O_pla_ands[26][4] ;
 wire \tms1x00.O_pla_ands[26][5] ;
 wire \tms1x00.O_pla_ands[26][6] ;
 wire \tms1x00.O_pla_ands[26][7] ;
 wire \tms1x00.O_pla_ands[26][8] ;
 wire \tms1x00.O_pla_ands[26][9] ;
 wire \tms1x00.O_pla_ands[27][0] ;
 wire \tms1x00.O_pla_ands[27][1] ;
 wire \tms1x00.O_pla_ands[27][2] ;
 wire \tms1x00.O_pla_ands[27][3] ;
 wire \tms1x00.O_pla_ands[27][4] ;
 wire \tms1x00.O_pla_ands[27][5] ;
 wire \tms1x00.O_pla_ands[27][6] ;
 wire \tms1x00.O_pla_ands[27][7] ;
 wire \tms1x00.O_pla_ands[27][8] ;
 wire \tms1x00.O_pla_ands[27][9] ;
 wire \tms1x00.O_pla_ands[28][0] ;
 wire \tms1x00.O_pla_ands[28][1] ;
 wire \tms1x00.O_pla_ands[28][2] ;
 wire \tms1x00.O_pla_ands[28][3] ;
 wire \tms1x00.O_pla_ands[28][4] ;
 wire \tms1x00.O_pla_ands[28][5] ;
 wire \tms1x00.O_pla_ands[28][6] ;
 wire \tms1x00.O_pla_ands[28][7] ;
 wire \tms1x00.O_pla_ands[28][8] ;
 wire \tms1x00.O_pla_ands[28][9] ;
 wire \tms1x00.O_pla_ands[29][0] ;
 wire \tms1x00.O_pla_ands[29][1] ;
 wire \tms1x00.O_pla_ands[29][2] ;
 wire \tms1x00.O_pla_ands[29][3] ;
 wire \tms1x00.O_pla_ands[29][4] ;
 wire \tms1x00.O_pla_ands[29][5] ;
 wire \tms1x00.O_pla_ands[29][6] ;
 wire \tms1x00.O_pla_ands[29][7] ;
 wire \tms1x00.O_pla_ands[29][8] ;
 wire \tms1x00.O_pla_ands[29][9] ;
 wire \tms1x00.O_pla_ands[2][0] ;
 wire \tms1x00.O_pla_ands[2][1] ;
 wire \tms1x00.O_pla_ands[2][2] ;
 wire \tms1x00.O_pla_ands[2][3] ;
 wire \tms1x00.O_pla_ands[2][4] ;
 wire \tms1x00.O_pla_ands[2][5] ;
 wire \tms1x00.O_pla_ands[2][6] ;
 wire \tms1x00.O_pla_ands[2][7] ;
 wire \tms1x00.O_pla_ands[2][8] ;
 wire \tms1x00.O_pla_ands[2][9] ;
 wire \tms1x00.O_pla_ands[30][0] ;
 wire \tms1x00.O_pla_ands[30][1] ;
 wire \tms1x00.O_pla_ands[30][2] ;
 wire \tms1x00.O_pla_ands[30][3] ;
 wire \tms1x00.O_pla_ands[30][4] ;
 wire \tms1x00.O_pla_ands[30][5] ;
 wire \tms1x00.O_pla_ands[30][6] ;
 wire \tms1x00.O_pla_ands[30][7] ;
 wire \tms1x00.O_pla_ands[30][8] ;
 wire \tms1x00.O_pla_ands[30][9] ;
 wire \tms1x00.O_pla_ands[31][0] ;
 wire \tms1x00.O_pla_ands[31][1] ;
 wire \tms1x00.O_pla_ands[31][2] ;
 wire \tms1x00.O_pla_ands[31][3] ;
 wire \tms1x00.O_pla_ands[31][4] ;
 wire \tms1x00.O_pla_ands[31][5] ;
 wire \tms1x00.O_pla_ands[31][6] ;
 wire \tms1x00.O_pla_ands[31][7] ;
 wire \tms1x00.O_pla_ands[31][8] ;
 wire \tms1x00.O_pla_ands[31][9] ;
 wire \tms1x00.O_pla_ands[3][0] ;
 wire \tms1x00.O_pla_ands[3][1] ;
 wire \tms1x00.O_pla_ands[3][2] ;
 wire \tms1x00.O_pla_ands[3][3] ;
 wire \tms1x00.O_pla_ands[3][4] ;
 wire \tms1x00.O_pla_ands[3][5] ;
 wire \tms1x00.O_pla_ands[3][6] ;
 wire \tms1x00.O_pla_ands[3][7] ;
 wire \tms1x00.O_pla_ands[3][8] ;
 wire \tms1x00.O_pla_ands[3][9] ;
 wire \tms1x00.O_pla_ands[4][0] ;
 wire \tms1x00.O_pla_ands[4][1] ;
 wire \tms1x00.O_pla_ands[4][2] ;
 wire \tms1x00.O_pla_ands[4][3] ;
 wire \tms1x00.O_pla_ands[4][4] ;
 wire \tms1x00.O_pla_ands[4][5] ;
 wire \tms1x00.O_pla_ands[4][6] ;
 wire \tms1x00.O_pla_ands[4][7] ;
 wire \tms1x00.O_pla_ands[4][8] ;
 wire \tms1x00.O_pla_ands[4][9] ;
 wire \tms1x00.O_pla_ands[5][0] ;
 wire \tms1x00.O_pla_ands[5][1] ;
 wire \tms1x00.O_pla_ands[5][2] ;
 wire \tms1x00.O_pla_ands[5][3] ;
 wire \tms1x00.O_pla_ands[5][4] ;
 wire \tms1x00.O_pla_ands[5][5] ;
 wire \tms1x00.O_pla_ands[5][6] ;
 wire \tms1x00.O_pla_ands[5][7] ;
 wire \tms1x00.O_pla_ands[5][8] ;
 wire \tms1x00.O_pla_ands[5][9] ;
 wire \tms1x00.O_pla_ands[6][0] ;
 wire \tms1x00.O_pla_ands[6][1] ;
 wire \tms1x00.O_pla_ands[6][2] ;
 wire \tms1x00.O_pla_ands[6][3] ;
 wire \tms1x00.O_pla_ands[6][4] ;
 wire \tms1x00.O_pla_ands[6][5] ;
 wire \tms1x00.O_pla_ands[6][6] ;
 wire \tms1x00.O_pla_ands[6][7] ;
 wire \tms1x00.O_pla_ands[6][8] ;
 wire \tms1x00.O_pla_ands[6][9] ;
 wire \tms1x00.O_pla_ands[7][0] ;
 wire \tms1x00.O_pla_ands[7][1] ;
 wire \tms1x00.O_pla_ands[7][2] ;
 wire \tms1x00.O_pla_ands[7][3] ;
 wire \tms1x00.O_pla_ands[7][4] ;
 wire \tms1x00.O_pla_ands[7][5] ;
 wire \tms1x00.O_pla_ands[7][6] ;
 wire \tms1x00.O_pla_ands[7][7] ;
 wire \tms1x00.O_pla_ands[7][8] ;
 wire \tms1x00.O_pla_ands[7][9] ;
 wire \tms1x00.O_pla_ands[8][0] ;
 wire \tms1x00.O_pla_ands[8][1] ;
 wire \tms1x00.O_pla_ands[8][2] ;
 wire \tms1x00.O_pla_ands[8][3] ;
 wire \tms1x00.O_pla_ands[8][4] ;
 wire \tms1x00.O_pla_ands[8][5] ;
 wire \tms1x00.O_pla_ands[8][6] ;
 wire \tms1x00.O_pla_ands[8][7] ;
 wire \tms1x00.O_pla_ands[8][8] ;
 wire \tms1x00.O_pla_ands[8][9] ;
 wire \tms1x00.O_pla_ands[9][0] ;
 wire \tms1x00.O_pla_ands[9][1] ;
 wire \tms1x00.O_pla_ands[9][2] ;
 wire \tms1x00.O_pla_ands[9][3] ;
 wire \tms1x00.O_pla_ands[9][4] ;
 wire \tms1x00.O_pla_ands[9][5] ;
 wire \tms1x00.O_pla_ands[9][6] ;
 wire \tms1x00.O_pla_ands[9][7] ;
 wire \tms1x00.O_pla_ands[9][8] ;
 wire \tms1x00.O_pla_ands[9][9] ;
 wire \tms1x00.O_pla_ors[0][0] ;
 wire \tms1x00.O_pla_ors[0][10] ;
 wire \tms1x00.O_pla_ors[0][11] ;
 wire \tms1x00.O_pla_ors[0][12] ;
 wire \tms1x00.O_pla_ors[0][13] ;
 wire \tms1x00.O_pla_ors[0][14] ;
 wire \tms1x00.O_pla_ors[0][15] ;
 wire \tms1x00.O_pla_ors[0][16] ;
 wire \tms1x00.O_pla_ors[0][17] ;
 wire \tms1x00.O_pla_ors[0][18] ;
 wire \tms1x00.O_pla_ors[0][19] ;
 wire \tms1x00.O_pla_ors[0][1] ;
 wire \tms1x00.O_pla_ors[0][2] ;
 wire \tms1x00.O_pla_ors[0][3] ;
 wire \tms1x00.O_pla_ors[0][4] ;
 wire \tms1x00.O_pla_ors[0][5] ;
 wire \tms1x00.O_pla_ors[0][6] ;
 wire \tms1x00.O_pla_ors[0][7] ;
 wire \tms1x00.O_pla_ors[0][8] ;
 wire \tms1x00.O_pla_ors[0][9] ;
 wire \tms1x00.O_pla_ors[1][0] ;
 wire \tms1x00.O_pla_ors[1][10] ;
 wire \tms1x00.O_pla_ors[1][11] ;
 wire \tms1x00.O_pla_ors[1][12] ;
 wire \tms1x00.O_pla_ors[1][13] ;
 wire \tms1x00.O_pla_ors[1][14] ;
 wire \tms1x00.O_pla_ors[1][15] ;
 wire \tms1x00.O_pla_ors[1][16] ;
 wire \tms1x00.O_pla_ors[1][17] ;
 wire \tms1x00.O_pla_ors[1][18] ;
 wire \tms1x00.O_pla_ors[1][19] ;
 wire \tms1x00.O_pla_ors[1][1] ;
 wire \tms1x00.O_pla_ors[1][2] ;
 wire \tms1x00.O_pla_ors[1][3] ;
 wire \tms1x00.O_pla_ors[1][4] ;
 wire \tms1x00.O_pla_ors[1][5] ;
 wire \tms1x00.O_pla_ors[1][6] ;
 wire \tms1x00.O_pla_ors[1][7] ;
 wire \tms1x00.O_pla_ors[1][8] ;
 wire \tms1x00.O_pla_ors[1][9] ;
 wire \tms1x00.O_pla_ors[2][0] ;
 wire \tms1x00.O_pla_ors[2][10] ;
 wire \tms1x00.O_pla_ors[2][11] ;
 wire \tms1x00.O_pla_ors[2][12] ;
 wire \tms1x00.O_pla_ors[2][13] ;
 wire \tms1x00.O_pla_ors[2][14] ;
 wire \tms1x00.O_pla_ors[2][15] ;
 wire \tms1x00.O_pla_ors[2][16] ;
 wire \tms1x00.O_pla_ors[2][17] ;
 wire \tms1x00.O_pla_ors[2][18] ;
 wire \tms1x00.O_pla_ors[2][19] ;
 wire \tms1x00.O_pla_ors[2][1] ;
 wire \tms1x00.O_pla_ors[2][2] ;
 wire \tms1x00.O_pla_ors[2][3] ;
 wire \tms1x00.O_pla_ors[2][4] ;
 wire \tms1x00.O_pla_ors[2][5] ;
 wire \tms1x00.O_pla_ors[2][6] ;
 wire \tms1x00.O_pla_ors[2][7] ;
 wire \tms1x00.O_pla_ors[2][8] ;
 wire \tms1x00.O_pla_ors[2][9] ;
 wire \tms1x00.O_pla_ors[3][0] ;
 wire \tms1x00.O_pla_ors[3][10] ;
 wire \tms1x00.O_pla_ors[3][11] ;
 wire \tms1x00.O_pla_ors[3][12] ;
 wire \tms1x00.O_pla_ors[3][13] ;
 wire \tms1x00.O_pla_ors[3][14] ;
 wire \tms1x00.O_pla_ors[3][15] ;
 wire \tms1x00.O_pla_ors[3][16] ;
 wire \tms1x00.O_pla_ors[3][17] ;
 wire \tms1x00.O_pla_ors[3][18] ;
 wire \tms1x00.O_pla_ors[3][19] ;
 wire \tms1x00.O_pla_ors[3][1] ;
 wire \tms1x00.O_pla_ors[3][2] ;
 wire \tms1x00.O_pla_ors[3][3] ;
 wire \tms1x00.O_pla_ors[3][4] ;
 wire \tms1x00.O_pla_ors[3][5] ;
 wire \tms1x00.O_pla_ors[3][6] ;
 wire \tms1x00.O_pla_ors[3][7] ;
 wire \tms1x00.O_pla_ors[3][8] ;
 wire \tms1x00.O_pla_ors[3][9] ;
 wire \tms1x00.O_pla_ors[4][0] ;
 wire \tms1x00.O_pla_ors[4][10] ;
 wire \tms1x00.O_pla_ors[4][11] ;
 wire \tms1x00.O_pla_ors[4][12] ;
 wire \tms1x00.O_pla_ors[4][13] ;
 wire \tms1x00.O_pla_ors[4][14] ;
 wire \tms1x00.O_pla_ors[4][15] ;
 wire \tms1x00.O_pla_ors[4][16] ;
 wire \tms1x00.O_pla_ors[4][17] ;
 wire \tms1x00.O_pla_ors[4][18] ;
 wire \tms1x00.O_pla_ors[4][19] ;
 wire \tms1x00.O_pla_ors[4][1] ;
 wire \tms1x00.O_pla_ors[4][2] ;
 wire \tms1x00.O_pla_ors[4][3] ;
 wire \tms1x00.O_pla_ors[4][4] ;
 wire \tms1x00.O_pla_ors[4][5] ;
 wire \tms1x00.O_pla_ors[4][6] ;
 wire \tms1x00.O_pla_ors[4][7] ;
 wire \tms1x00.O_pla_ors[4][8] ;
 wire \tms1x00.O_pla_ors[4][9] ;
 wire \tms1x00.O_pla_ors[5][0] ;
 wire \tms1x00.O_pla_ors[5][10] ;
 wire \tms1x00.O_pla_ors[5][11] ;
 wire \tms1x00.O_pla_ors[5][12] ;
 wire \tms1x00.O_pla_ors[5][13] ;
 wire \tms1x00.O_pla_ors[5][14] ;
 wire \tms1x00.O_pla_ors[5][15] ;
 wire \tms1x00.O_pla_ors[5][16] ;
 wire \tms1x00.O_pla_ors[5][17] ;
 wire \tms1x00.O_pla_ors[5][18] ;
 wire \tms1x00.O_pla_ors[5][19] ;
 wire \tms1x00.O_pla_ors[5][1] ;
 wire \tms1x00.O_pla_ors[5][2] ;
 wire \tms1x00.O_pla_ors[5][3] ;
 wire \tms1x00.O_pla_ors[5][4] ;
 wire \tms1x00.O_pla_ors[5][5] ;
 wire \tms1x00.O_pla_ors[5][6] ;
 wire \tms1x00.O_pla_ors[5][7] ;
 wire \tms1x00.O_pla_ors[5][8] ;
 wire \tms1x00.O_pla_ors[5][9] ;
 wire \tms1x00.O_pla_ors[6][0] ;
 wire \tms1x00.O_pla_ors[6][10] ;
 wire \tms1x00.O_pla_ors[6][11] ;
 wire \tms1x00.O_pla_ors[6][12] ;
 wire \tms1x00.O_pla_ors[6][13] ;
 wire \tms1x00.O_pla_ors[6][14] ;
 wire \tms1x00.O_pla_ors[6][15] ;
 wire \tms1x00.O_pla_ors[6][16] ;
 wire \tms1x00.O_pla_ors[6][17] ;
 wire \tms1x00.O_pla_ors[6][18] ;
 wire \tms1x00.O_pla_ors[6][19] ;
 wire \tms1x00.O_pla_ors[6][1] ;
 wire \tms1x00.O_pla_ors[6][2] ;
 wire \tms1x00.O_pla_ors[6][3] ;
 wire \tms1x00.O_pla_ors[6][4] ;
 wire \tms1x00.O_pla_ors[6][5] ;
 wire \tms1x00.O_pla_ors[6][6] ;
 wire \tms1x00.O_pla_ors[6][7] ;
 wire \tms1x00.O_pla_ors[6][8] ;
 wire \tms1x00.O_pla_ors[6][9] ;
 wire \tms1x00.O_pla_ors[7][0] ;
 wire \tms1x00.O_pla_ors[7][10] ;
 wire \tms1x00.O_pla_ors[7][11] ;
 wire \tms1x00.O_pla_ors[7][12] ;
 wire \tms1x00.O_pla_ors[7][13] ;
 wire \tms1x00.O_pla_ors[7][14] ;
 wire \tms1x00.O_pla_ors[7][15] ;
 wire \tms1x00.O_pla_ors[7][16] ;
 wire \tms1x00.O_pla_ors[7][17] ;
 wire \tms1x00.O_pla_ors[7][18] ;
 wire \tms1x00.O_pla_ors[7][19] ;
 wire \tms1x00.O_pla_ors[7][1] ;
 wire \tms1x00.O_pla_ors[7][2] ;
 wire \tms1x00.O_pla_ors[7][3] ;
 wire \tms1x00.O_pla_ors[7][4] ;
 wire \tms1x00.O_pla_ors[7][5] ;
 wire \tms1x00.O_pla_ors[7][6] ;
 wire \tms1x00.O_pla_ors[7][7] ;
 wire \tms1x00.O_pla_ors[7][8] ;
 wire \tms1x00.O_pla_ors[7][9] ;
 wire \tms1x00.PA[0] ;
 wire \tms1x00.PA[1] ;
 wire \tms1x00.PA[2] ;
 wire \tms1x00.PA[3] ;
 wire \tms1x00.PB[0] ;
 wire \tms1x00.PB[1] ;
 wire \tms1x00.PB[2] ;
 wire \tms1x00.PB[3] ;
 wire \tms1x00.PC[0] ;
 wire \tms1x00.PC[1] ;
 wire \tms1x00.PC[2] ;
 wire \tms1x00.PC[3] ;
 wire \tms1x00.PC[4] ;
 wire \tms1x00.PC[5] ;
 wire \tms1x00.P[0] ;
 wire \tms1x00.P[1] ;
 wire \tms1x00.P[2] ;
 wire \tms1x00.P[3] ;
 wire \tms1x00.SL ;
 wire \tms1x00.SR[0] ;
 wire \tms1x00.SR[1] ;
 wire \tms1x00.SR[2] ;
 wire \tms1x00.SR[3] ;
 wire \tms1x00.SR[4] ;
 wire \tms1x00.SR[5] ;
 wire \tms1x00.X[0] ;
 wire \tms1x00.X[1] ;
 wire \tms1x00.X[2] ;
 wire \tms1x00.Y[0] ;
 wire \tms1x00.Y[1] ;
 wire \tms1x00.Y[2] ;
 wire \tms1x00.Y[3] ;
 wire \tms1x00.cycle[0] ;
 wire \tms1x00.cycle[1] ;
 wire \tms1x00.cycle[2] ;
 wire \tms1x00.ins_arg[0] ;
 wire \tms1x00.ins_arg[1] ;
 wire \tms1x00.ins_arg[2] ;
 wire \tms1x00.ins_arg[3] ;
 wire \tms1x00.ins_arg[4] ;
 wire \tms1x00.ins_arg[5] ;
 wire \tms1x00.ins_pla_ands[0][0] ;
 wire \tms1x00.ins_pla_ands[0][10] ;
 wire \tms1x00.ins_pla_ands[0][11] ;
 wire \tms1x00.ins_pla_ands[0][12] ;
 wire \tms1x00.ins_pla_ands[0][13] ;
 wire \tms1x00.ins_pla_ands[0][14] ;
 wire \tms1x00.ins_pla_ands[0][15] ;
 wire \tms1x00.ins_pla_ands[0][1] ;
 wire \tms1x00.ins_pla_ands[0][2] ;
 wire \tms1x00.ins_pla_ands[0][3] ;
 wire \tms1x00.ins_pla_ands[0][4] ;
 wire \tms1x00.ins_pla_ands[0][5] ;
 wire \tms1x00.ins_pla_ands[0][6] ;
 wire \tms1x00.ins_pla_ands[0][7] ;
 wire \tms1x00.ins_pla_ands[0][8] ;
 wire \tms1x00.ins_pla_ands[0][9] ;
 wire \tms1x00.ins_pla_ands[10][0] ;
 wire \tms1x00.ins_pla_ands[10][10] ;
 wire \tms1x00.ins_pla_ands[10][11] ;
 wire \tms1x00.ins_pla_ands[10][12] ;
 wire \tms1x00.ins_pla_ands[10][13] ;
 wire \tms1x00.ins_pla_ands[10][14] ;
 wire \tms1x00.ins_pla_ands[10][15] ;
 wire \tms1x00.ins_pla_ands[10][1] ;
 wire \tms1x00.ins_pla_ands[10][2] ;
 wire \tms1x00.ins_pla_ands[10][3] ;
 wire \tms1x00.ins_pla_ands[10][4] ;
 wire \tms1x00.ins_pla_ands[10][5] ;
 wire \tms1x00.ins_pla_ands[10][6] ;
 wire \tms1x00.ins_pla_ands[10][7] ;
 wire \tms1x00.ins_pla_ands[10][8] ;
 wire \tms1x00.ins_pla_ands[10][9] ;
 wire \tms1x00.ins_pla_ands[11][0] ;
 wire \tms1x00.ins_pla_ands[11][10] ;
 wire \tms1x00.ins_pla_ands[11][11] ;
 wire \tms1x00.ins_pla_ands[11][12] ;
 wire \tms1x00.ins_pla_ands[11][13] ;
 wire \tms1x00.ins_pla_ands[11][14] ;
 wire \tms1x00.ins_pla_ands[11][15] ;
 wire \tms1x00.ins_pla_ands[11][1] ;
 wire \tms1x00.ins_pla_ands[11][2] ;
 wire \tms1x00.ins_pla_ands[11][3] ;
 wire \tms1x00.ins_pla_ands[11][4] ;
 wire \tms1x00.ins_pla_ands[11][5] ;
 wire \tms1x00.ins_pla_ands[11][6] ;
 wire \tms1x00.ins_pla_ands[11][7] ;
 wire \tms1x00.ins_pla_ands[11][8] ;
 wire \tms1x00.ins_pla_ands[11][9] ;
 wire \tms1x00.ins_pla_ands[12][0] ;
 wire \tms1x00.ins_pla_ands[12][10] ;
 wire \tms1x00.ins_pla_ands[12][11] ;
 wire \tms1x00.ins_pla_ands[12][12] ;
 wire \tms1x00.ins_pla_ands[12][13] ;
 wire \tms1x00.ins_pla_ands[12][14] ;
 wire \tms1x00.ins_pla_ands[12][15] ;
 wire \tms1x00.ins_pla_ands[12][1] ;
 wire \tms1x00.ins_pla_ands[12][2] ;
 wire \tms1x00.ins_pla_ands[12][3] ;
 wire \tms1x00.ins_pla_ands[12][4] ;
 wire \tms1x00.ins_pla_ands[12][5] ;
 wire \tms1x00.ins_pla_ands[12][6] ;
 wire \tms1x00.ins_pla_ands[12][7] ;
 wire \tms1x00.ins_pla_ands[12][8] ;
 wire \tms1x00.ins_pla_ands[12][9] ;
 wire \tms1x00.ins_pla_ands[13][0] ;
 wire \tms1x00.ins_pla_ands[13][10] ;
 wire \tms1x00.ins_pla_ands[13][11] ;
 wire \tms1x00.ins_pla_ands[13][12] ;
 wire \tms1x00.ins_pla_ands[13][13] ;
 wire \tms1x00.ins_pla_ands[13][14] ;
 wire \tms1x00.ins_pla_ands[13][15] ;
 wire \tms1x00.ins_pla_ands[13][1] ;
 wire \tms1x00.ins_pla_ands[13][2] ;
 wire \tms1x00.ins_pla_ands[13][3] ;
 wire \tms1x00.ins_pla_ands[13][4] ;
 wire \tms1x00.ins_pla_ands[13][5] ;
 wire \tms1x00.ins_pla_ands[13][6] ;
 wire \tms1x00.ins_pla_ands[13][7] ;
 wire \tms1x00.ins_pla_ands[13][8] ;
 wire \tms1x00.ins_pla_ands[13][9] ;
 wire \tms1x00.ins_pla_ands[14][0] ;
 wire \tms1x00.ins_pla_ands[14][10] ;
 wire \tms1x00.ins_pla_ands[14][11] ;
 wire \tms1x00.ins_pla_ands[14][12] ;
 wire \tms1x00.ins_pla_ands[14][13] ;
 wire \tms1x00.ins_pla_ands[14][14] ;
 wire \tms1x00.ins_pla_ands[14][15] ;
 wire \tms1x00.ins_pla_ands[14][1] ;
 wire \tms1x00.ins_pla_ands[14][2] ;
 wire \tms1x00.ins_pla_ands[14][3] ;
 wire \tms1x00.ins_pla_ands[14][4] ;
 wire \tms1x00.ins_pla_ands[14][5] ;
 wire \tms1x00.ins_pla_ands[14][6] ;
 wire \tms1x00.ins_pla_ands[14][7] ;
 wire \tms1x00.ins_pla_ands[14][8] ;
 wire \tms1x00.ins_pla_ands[14][9] ;
 wire \tms1x00.ins_pla_ands[15][0] ;
 wire \tms1x00.ins_pla_ands[15][10] ;
 wire \tms1x00.ins_pla_ands[15][11] ;
 wire \tms1x00.ins_pla_ands[15][12] ;
 wire \tms1x00.ins_pla_ands[15][13] ;
 wire \tms1x00.ins_pla_ands[15][14] ;
 wire \tms1x00.ins_pla_ands[15][15] ;
 wire \tms1x00.ins_pla_ands[15][1] ;
 wire \tms1x00.ins_pla_ands[15][2] ;
 wire \tms1x00.ins_pla_ands[15][3] ;
 wire \tms1x00.ins_pla_ands[15][4] ;
 wire \tms1x00.ins_pla_ands[15][5] ;
 wire \tms1x00.ins_pla_ands[15][6] ;
 wire \tms1x00.ins_pla_ands[15][7] ;
 wire \tms1x00.ins_pla_ands[15][8] ;
 wire \tms1x00.ins_pla_ands[15][9] ;
 wire \tms1x00.ins_pla_ands[16][0] ;
 wire \tms1x00.ins_pla_ands[16][10] ;
 wire \tms1x00.ins_pla_ands[16][11] ;
 wire \tms1x00.ins_pla_ands[16][12] ;
 wire \tms1x00.ins_pla_ands[16][13] ;
 wire \tms1x00.ins_pla_ands[16][14] ;
 wire \tms1x00.ins_pla_ands[16][15] ;
 wire \tms1x00.ins_pla_ands[16][1] ;
 wire \tms1x00.ins_pla_ands[16][2] ;
 wire \tms1x00.ins_pla_ands[16][3] ;
 wire \tms1x00.ins_pla_ands[16][4] ;
 wire \tms1x00.ins_pla_ands[16][5] ;
 wire \tms1x00.ins_pla_ands[16][6] ;
 wire \tms1x00.ins_pla_ands[16][7] ;
 wire \tms1x00.ins_pla_ands[16][8] ;
 wire \tms1x00.ins_pla_ands[16][9] ;
 wire \tms1x00.ins_pla_ands[17][0] ;
 wire \tms1x00.ins_pla_ands[17][10] ;
 wire \tms1x00.ins_pla_ands[17][11] ;
 wire \tms1x00.ins_pla_ands[17][12] ;
 wire \tms1x00.ins_pla_ands[17][13] ;
 wire \tms1x00.ins_pla_ands[17][14] ;
 wire \tms1x00.ins_pla_ands[17][15] ;
 wire \tms1x00.ins_pla_ands[17][1] ;
 wire \tms1x00.ins_pla_ands[17][2] ;
 wire \tms1x00.ins_pla_ands[17][3] ;
 wire \tms1x00.ins_pla_ands[17][4] ;
 wire \tms1x00.ins_pla_ands[17][5] ;
 wire \tms1x00.ins_pla_ands[17][6] ;
 wire \tms1x00.ins_pla_ands[17][7] ;
 wire \tms1x00.ins_pla_ands[17][8] ;
 wire \tms1x00.ins_pla_ands[17][9] ;
 wire \tms1x00.ins_pla_ands[18][0] ;
 wire \tms1x00.ins_pla_ands[18][10] ;
 wire \tms1x00.ins_pla_ands[18][11] ;
 wire \tms1x00.ins_pla_ands[18][12] ;
 wire \tms1x00.ins_pla_ands[18][13] ;
 wire \tms1x00.ins_pla_ands[18][14] ;
 wire \tms1x00.ins_pla_ands[18][15] ;
 wire \tms1x00.ins_pla_ands[18][1] ;
 wire \tms1x00.ins_pla_ands[18][2] ;
 wire \tms1x00.ins_pla_ands[18][3] ;
 wire \tms1x00.ins_pla_ands[18][4] ;
 wire \tms1x00.ins_pla_ands[18][5] ;
 wire \tms1x00.ins_pla_ands[18][6] ;
 wire \tms1x00.ins_pla_ands[18][7] ;
 wire \tms1x00.ins_pla_ands[18][8] ;
 wire \tms1x00.ins_pla_ands[18][9] ;
 wire \tms1x00.ins_pla_ands[19][0] ;
 wire \tms1x00.ins_pla_ands[19][10] ;
 wire \tms1x00.ins_pla_ands[19][11] ;
 wire \tms1x00.ins_pla_ands[19][12] ;
 wire \tms1x00.ins_pla_ands[19][13] ;
 wire \tms1x00.ins_pla_ands[19][14] ;
 wire \tms1x00.ins_pla_ands[19][15] ;
 wire \tms1x00.ins_pla_ands[19][1] ;
 wire \tms1x00.ins_pla_ands[19][2] ;
 wire \tms1x00.ins_pla_ands[19][3] ;
 wire \tms1x00.ins_pla_ands[19][4] ;
 wire \tms1x00.ins_pla_ands[19][5] ;
 wire \tms1x00.ins_pla_ands[19][6] ;
 wire \tms1x00.ins_pla_ands[19][7] ;
 wire \tms1x00.ins_pla_ands[19][8] ;
 wire \tms1x00.ins_pla_ands[19][9] ;
 wire \tms1x00.ins_pla_ands[1][0] ;
 wire \tms1x00.ins_pla_ands[1][10] ;
 wire \tms1x00.ins_pla_ands[1][11] ;
 wire \tms1x00.ins_pla_ands[1][12] ;
 wire \tms1x00.ins_pla_ands[1][13] ;
 wire \tms1x00.ins_pla_ands[1][14] ;
 wire \tms1x00.ins_pla_ands[1][15] ;
 wire \tms1x00.ins_pla_ands[1][1] ;
 wire \tms1x00.ins_pla_ands[1][2] ;
 wire \tms1x00.ins_pla_ands[1][3] ;
 wire \tms1x00.ins_pla_ands[1][4] ;
 wire \tms1x00.ins_pla_ands[1][5] ;
 wire \tms1x00.ins_pla_ands[1][6] ;
 wire \tms1x00.ins_pla_ands[1][7] ;
 wire \tms1x00.ins_pla_ands[1][8] ;
 wire \tms1x00.ins_pla_ands[1][9] ;
 wire \tms1x00.ins_pla_ands[20][0] ;
 wire \tms1x00.ins_pla_ands[20][10] ;
 wire \tms1x00.ins_pla_ands[20][11] ;
 wire \tms1x00.ins_pla_ands[20][12] ;
 wire \tms1x00.ins_pla_ands[20][13] ;
 wire \tms1x00.ins_pla_ands[20][14] ;
 wire \tms1x00.ins_pla_ands[20][15] ;
 wire \tms1x00.ins_pla_ands[20][1] ;
 wire \tms1x00.ins_pla_ands[20][2] ;
 wire \tms1x00.ins_pla_ands[20][3] ;
 wire \tms1x00.ins_pla_ands[20][4] ;
 wire \tms1x00.ins_pla_ands[20][5] ;
 wire \tms1x00.ins_pla_ands[20][6] ;
 wire \tms1x00.ins_pla_ands[20][7] ;
 wire \tms1x00.ins_pla_ands[20][8] ;
 wire \tms1x00.ins_pla_ands[20][9] ;
 wire \tms1x00.ins_pla_ands[21][0] ;
 wire \tms1x00.ins_pla_ands[21][10] ;
 wire \tms1x00.ins_pla_ands[21][11] ;
 wire \tms1x00.ins_pla_ands[21][12] ;
 wire \tms1x00.ins_pla_ands[21][13] ;
 wire \tms1x00.ins_pla_ands[21][14] ;
 wire \tms1x00.ins_pla_ands[21][15] ;
 wire \tms1x00.ins_pla_ands[21][1] ;
 wire \tms1x00.ins_pla_ands[21][2] ;
 wire \tms1x00.ins_pla_ands[21][3] ;
 wire \tms1x00.ins_pla_ands[21][4] ;
 wire \tms1x00.ins_pla_ands[21][5] ;
 wire \tms1x00.ins_pla_ands[21][6] ;
 wire \tms1x00.ins_pla_ands[21][7] ;
 wire \tms1x00.ins_pla_ands[21][8] ;
 wire \tms1x00.ins_pla_ands[21][9] ;
 wire \tms1x00.ins_pla_ands[22][0] ;
 wire \tms1x00.ins_pla_ands[22][10] ;
 wire \tms1x00.ins_pla_ands[22][11] ;
 wire \tms1x00.ins_pla_ands[22][12] ;
 wire \tms1x00.ins_pla_ands[22][13] ;
 wire \tms1x00.ins_pla_ands[22][14] ;
 wire \tms1x00.ins_pla_ands[22][15] ;
 wire \tms1x00.ins_pla_ands[22][1] ;
 wire \tms1x00.ins_pla_ands[22][2] ;
 wire \tms1x00.ins_pla_ands[22][3] ;
 wire \tms1x00.ins_pla_ands[22][4] ;
 wire \tms1x00.ins_pla_ands[22][5] ;
 wire \tms1x00.ins_pla_ands[22][6] ;
 wire \tms1x00.ins_pla_ands[22][7] ;
 wire \tms1x00.ins_pla_ands[22][8] ;
 wire \tms1x00.ins_pla_ands[22][9] ;
 wire \tms1x00.ins_pla_ands[23][0] ;
 wire \tms1x00.ins_pla_ands[23][10] ;
 wire \tms1x00.ins_pla_ands[23][11] ;
 wire \tms1x00.ins_pla_ands[23][12] ;
 wire \tms1x00.ins_pla_ands[23][13] ;
 wire \tms1x00.ins_pla_ands[23][14] ;
 wire \tms1x00.ins_pla_ands[23][15] ;
 wire \tms1x00.ins_pla_ands[23][1] ;
 wire \tms1x00.ins_pla_ands[23][2] ;
 wire \tms1x00.ins_pla_ands[23][3] ;
 wire \tms1x00.ins_pla_ands[23][4] ;
 wire \tms1x00.ins_pla_ands[23][5] ;
 wire \tms1x00.ins_pla_ands[23][6] ;
 wire \tms1x00.ins_pla_ands[23][7] ;
 wire \tms1x00.ins_pla_ands[23][8] ;
 wire \tms1x00.ins_pla_ands[23][9] ;
 wire \tms1x00.ins_pla_ands[24][0] ;
 wire \tms1x00.ins_pla_ands[24][10] ;
 wire \tms1x00.ins_pla_ands[24][11] ;
 wire \tms1x00.ins_pla_ands[24][12] ;
 wire \tms1x00.ins_pla_ands[24][13] ;
 wire \tms1x00.ins_pla_ands[24][14] ;
 wire \tms1x00.ins_pla_ands[24][15] ;
 wire \tms1x00.ins_pla_ands[24][1] ;
 wire \tms1x00.ins_pla_ands[24][2] ;
 wire \tms1x00.ins_pla_ands[24][3] ;
 wire \tms1x00.ins_pla_ands[24][4] ;
 wire \tms1x00.ins_pla_ands[24][5] ;
 wire \tms1x00.ins_pla_ands[24][6] ;
 wire \tms1x00.ins_pla_ands[24][7] ;
 wire \tms1x00.ins_pla_ands[24][8] ;
 wire \tms1x00.ins_pla_ands[24][9] ;
 wire \tms1x00.ins_pla_ands[25][0] ;
 wire \tms1x00.ins_pla_ands[25][10] ;
 wire \tms1x00.ins_pla_ands[25][11] ;
 wire \tms1x00.ins_pla_ands[25][12] ;
 wire \tms1x00.ins_pla_ands[25][13] ;
 wire \tms1x00.ins_pla_ands[25][14] ;
 wire \tms1x00.ins_pla_ands[25][15] ;
 wire \tms1x00.ins_pla_ands[25][1] ;
 wire \tms1x00.ins_pla_ands[25][2] ;
 wire \tms1x00.ins_pla_ands[25][3] ;
 wire \tms1x00.ins_pla_ands[25][4] ;
 wire \tms1x00.ins_pla_ands[25][5] ;
 wire \tms1x00.ins_pla_ands[25][6] ;
 wire \tms1x00.ins_pla_ands[25][7] ;
 wire \tms1x00.ins_pla_ands[25][8] ;
 wire \tms1x00.ins_pla_ands[25][9] ;
 wire \tms1x00.ins_pla_ands[26][0] ;
 wire \tms1x00.ins_pla_ands[26][10] ;
 wire \tms1x00.ins_pla_ands[26][11] ;
 wire \tms1x00.ins_pla_ands[26][12] ;
 wire \tms1x00.ins_pla_ands[26][13] ;
 wire \tms1x00.ins_pla_ands[26][14] ;
 wire \tms1x00.ins_pla_ands[26][15] ;
 wire \tms1x00.ins_pla_ands[26][1] ;
 wire \tms1x00.ins_pla_ands[26][2] ;
 wire \tms1x00.ins_pla_ands[26][3] ;
 wire \tms1x00.ins_pla_ands[26][4] ;
 wire \tms1x00.ins_pla_ands[26][5] ;
 wire \tms1x00.ins_pla_ands[26][6] ;
 wire \tms1x00.ins_pla_ands[26][7] ;
 wire \tms1x00.ins_pla_ands[26][8] ;
 wire \tms1x00.ins_pla_ands[26][9] ;
 wire \tms1x00.ins_pla_ands[27][0] ;
 wire \tms1x00.ins_pla_ands[27][10] ;
 wire \tms1x00.ins_pla_ands[27][11] ;
 wire \tms1x00.ins_pla_ands[27][12] ;
 wire \tms1x00.ins_pla_ands[27][13] ;
 wire \tms1x00.ins_pla_ands[27][14] ;
 wire \tms1x00.ins_pla_ands[27][15] ;
 wire \tms1x00.ins_pla_ands[27][1] ;
 wire \tms1x00.ins_pla_ands[27][2] ;
 wire \tms1x00.ins_pla_ands[27][3] ;
 wire \tms1x00.ins_pla_ands[27][4] ;
 wire \tms1x00.ins_pla_ands[27][5] ;
 wire \tms1x00.ins_pla_ands[27][6] ;
 wire \tms1x00.ins_pla_ands[27][7] ;
 wire \tms1x00.ins_pla_ands[27][8] ;
 wire \tms1x00.ins_pla_ands[27][9] ;
 wire \tms1x00.ins_pla_ands[28][0] ;
 wire \tms1x00.ins_pla_ands[28][10] ;
 wire \tms1x00.ins_pla_ands[28][11] ;
 wire \tms1x00.ins_pla_ands[28][12] ;
 wire \tms1x00.ins_pla_ands[28][13] ;
 wire \tms1x00.ins_pla_ands[28][14] ;
 wire \tms1x00.ins_pla_ands[28][15] ;
 wire \tms1x00.ins_pla_ands[28][1] ;
 wire \tms1x00.ins_pla_ands[28][2] ;
 wire \tms1x00.ins_pla_ands[28][3] ;
 wire \tms1x00.ins_pla_ands[28][4] ;
 wire \tms1x00.ins_pla_ands[28][5] ;
 wire \tms1x00.ins_pla_ands[28][6] ;
 wire \tms1x00.ins_pla_ands[28][7] ;
 wire \tms1x00.ins_pla_ands[28][8] ;
 wire \tms1x00.ins_pla_ands[28][9] ;
 wire \tms1x00.ins_pla_ands[29][0] ;
 wire \tms1x00.ins_pla_ands[29][10] ;
 wire \tms1x00.ins_pla_ands[29][11] ;
 wire \tms1x00.ins_pla_ands[29][12] ;
 wire \tms1x00.ins_pla_ands[29][13] ;
 wire \tms1x00.ins_pla_ands[29][14] ;
 wire \tms1x00.ins_pla_ands[29][15] ;
 wire \tms1x00.ins_pla_ands[29][1] ;
 wire \tms1x00.ins_pla_ands[29][2] ;
 wire \tms1x00.ins_pla_ands[29][3] ;
 wire \tms1x00.ins_pla_ands[29][4] ;
 wire \tms1x00.ins_pla_ands[29][5] ;
 wire \tms1x00.ins_pla_ands[29][6] ;
 wire \tms1x00.ins_pla_ands[29][7] ;
 wire \tms1x00.ins_pla_ands[29][8] ;
 wire \tms1x00.ins_pla_ands[29][9] ;
 wire \tms1x00.ins_pla_ands[2][0] ;
 wire \tms1x00.ins_pla_ands[2][10] ;
 wire \tms1x00.ins_pla_ands[2][11] ;
 wire \tms1x00.ins_pla_ands[2][12] ;
 wire \tms1x00.ins_pla_ands[2][13] ;
 wire \tms1x00.ins_pla_ands[2][14] ;
 wire \tms1x00.ins_pla_ands[2][15] ;
 wire \tms1x00.ins_pla_ands[2][1] ;
 wire \tms1x00.ins_pla_ands[2][2] ;
 wire \tms1x00.ins_pla_ands[2][3] ;
 wire \tms1x00.ins_pla_ands[2][4] ;
 wire \tms1x00.ins_pla_ands[2][5] ;
 wire \tms1x00.ins_pla_ands[2][6] ;
 wire \tms1x00.ins_pla_ands[2][7] ;
 wire \tms1x00.ins_pla_ands[2][8] ;
 wire \tms1x00.ins_pla_ands[2][9] ;
 wire \tms1x00.ins_pla_ands[30][0] ;
 wire \tms1x00.ins_pla_ands[30][10] ;
 wire \tms1x00.ins_pla_ands[30][11] ;
 wire \tms1x00.ins_pla_ands[30][12] ;
 wire \tms1x00.ins_pla_ands[30][13] ;
 wire \tms1x00.ins_pla_ands[30][14] ;
 wire \tms1x00.ins_pla_ands[30][15] ;
 wire \tms1x00.ins_pla_ands[30][1] ;
 wire \tms1x00.ins_pla_ands[30][2] ;
 wire \tms1x00.ins_pla_ands[30][3] ;
 wire \tms1x00.ins_pla_ands[30][4] ;
 wire \tms1x00.ins_pla_ands[30][5] ;
 wire \tms1x00.ins_pla_ands[30][6] ;
 wire \tms1x00.ins_pla_ands[30][7] ;
 wire \tms1x00.ins_pla_ands[30][8] ;
 wire \tms1x00.ins_pla_ands[30][9] ;
 wire \tms1x00.ins_pla_ands[31][0] ;
 wire \tms1x00.ins_pla_ands[31][10] ;
 wire \tms1x00.ins_pla_ands[31][11] ;
 wire \tms1x00.ins_pla_ands[31][12] ;
 wire \tms1x00.ins_pla_ands[31][13] ;
 wire \tms1x00.ins_pla_ands[31][14] ;
 wire \tms1x00.ins_pla_ands[31][15] ;
 wire \tms1x00.ins_pla_ands[31][1] ;
 wire \tms1x00.ins_pla_ands[31][2] ;
 wire \tms1x00.ins_pla_ands[31][3] ;
 wire \tms1x00.ins_pla_ands[31][4] ;
 wire \tms1x00.ins_pla_ands[31][5] ;
 wire \tms1x00.ins_pla_ands[31][6] ;
 wire \tms1x00.ins_pla_ands[31][7] ;
 wire \tms1x00.ins_pla_ands[31][8] ;
 wire \tms1x00.ins_pla_ands[31][9] ;
 wire \tms1x00.ins_pla_ands[3][0] ;
 wire \tms1x00.ins_pla_ands[3][10] ;
 wire \tms1x00.ins_pla_ands[3][11] ;
 wire \tms1x00.ins_pla_ands[3][12] ;
 wire \tms1x00.ins_pla_ands[3][13] ;
 wire \tms1x00.ins_pla_ands[3][14] ;
 wire \tms1x00.ins_pla_ands[3][15] ;
 wire \tms1x00.ins_pla_ands[3][1] ;
 wire \tms1x00.ins_pla_ands[3][2] ;
 wire \tms1x00.ins_pla_ands[3][3] ;
 wire \tms1x00.ins_pla_ands[3][4] ;
 wire \tms1x00.ins_pla_ands[3][5] ;
 wire \tms1x00.ins_pla_ands[3][6] ;
 wire \tms1x00.ins_pla_ands[3][7] ;
 wire \tms1x00.ins_pla_ands[3][8] ;
 wire \tms1x00.ins_pla_ands[3][9] ;
 wire \tms1x00.ins_pla_ands[4][0] ;
 wire \tms1x00.ins_pla_ands[4][10] ;
 wire \tms1x00.ins_pla_ands[4][11] ;
 wire \tms1x00.ins_pla_ands[4][12] ;
 wire \tms1x00.ins_pla_ands[4][13] ;
 wire \tms1x00.ins_pla_ands[4][14] ;
 wire \tms1x00.ins_pla_ands[4][15] ;
 wire \tms1x00.ins_pla_ands[4][1] ;
 wire \tms1x00.ins_pla_ands[4][2] ;
 wire \tms1x00.ins_pla_ands[4][3] ;
 wire \tms1x00.ins_pla_ands[4][4] ;
 wire \tms1x00.ins_pla_ands[4][5] ;
 wire \tms1x00.ins_pla_ands[4][6] ;
 wire \tms1x00.ins_pla_ands[4][7] ;
 wire \tms1x00.ins_pla_ands[4][8] ;
 wire \tms1x00.ins_pla_ands[4][9] ;
 wire \tms1x00.ins_pla_ands[5][0] ;
 wire \tms1x00.ins_pla_ands[5][10] ;
 wire \tms1x00.ins_pla_ands[5][11] ;
 wire \tms1x00.ins_pla_ands[5][12] ;
 wire \tms1x00.ins_pla_ands[5][13] ;
 wire \tms1x00.ins_pla_ands[5][14] ;
 wire \tms1x00.ins_pla_ands[5][15] ;
 wire \tms1x00.ins_pla_ands[5][1] ;
 wire \tms1x00.ins_pla_ands[5][2] ;
 wire \tms1x00.ins_pla_ands[5][3] ;
 wire \tms1x00.ins_pla_ands[5][4] ;
 wire \tms1x00.ins_pla_ands[5][5] ;
 wire \tms1x00.ins_pla_ands[5][6] ;
 wire \tms1x00.ins_pla_ands[5][7] ;
 wire \tms1x00.ins_pla_ands[5][8] ;
 wire \tms1x00.ins_pla_ands[5][9] ;
 wire \tms1x00.ins_pla_ands[6][0] ;
 wire \tms1x00.ins_pla_ands[6][10] ;
 wire \tms1x00.ins_pla_ands[6][11] ;
 wire \tms1x00.ins_pla_ands[6][12] ;
 wire \tms1x00.ins_pla_ands[6][13] ;
 wire \tms1x00.ins_pla_ands[6][14] ;
 wire \tms1x00.ins_pla_ands[6][15] ;
 wire \tms1x00.ins_pla_ands[6][1] ;
 wire \tms1x00.ins_pla_ands[6][2] ;
 wire \tms1x00.ins_pla_ands[6][3] ;
 wire \tms1x00.ins_pla_ands[6][4] ;
 wire \tms1x00.ins_pla_ands[6][5] ;
 wire \tms1x00.ins_pla_ands[6][6] ;
 wire \tms1x00.ins_pla_ands[6][7] ;
 wire \tms1x00.ins_pla_ands[6][8] ;
 wire \tms1x00.ins_pla_ands[6][9] ;
 wire \tms1x00.ins_pla_ands[7][0] ;
 wire \tms1x00.ins_pla_ands[7][10] ;
 wire \tms1x00.ins_pla_ands[7][11] ;
 wire \tms1x00.ins_pla_ands[7][12] ;
 wire \tms1x00.ins_pla_ands[7][13] ;
 wire \tms1x00.ins_pla_ands[7][14] ;
 wire \tms1x00.ins_pla_ands[7][15] ;
 wire \tms1x00.ins_pla_ands[7][1] ;
 wire \tms1x00.ins_pla_ands[7][2] ;
 wire \tms1x00.ins_pla_ands[7][3] ;
 wire \tms1x00.ins_pla_ands[7][4] ;
 wire \tms1x00.ins_pla_ands[7][5] ;
 wire \tms1x00.ins_pla_ands[7][6] ;
 wire \tms1x00.ins_pla_ands[7][7] ;
 wire \tms1x00.ins_pla_ands[7][8] ;
 wire \tms1x00.ins_pla_ands[7][9] ;
 wire \tms1x00.ins_pla_ands[8][0] ;
 wire \tms1x00.ins_pla_ands[8][10] ;
 wire \tms1x00.ins_pla_ands[8][11] ;
 wire \tms1x00.ins_pla_ands[8][12] ;
 wire \tms1x00.ins_pla_ands[8][13] ;
 wire \tms1x00.ins_pla_ands[8][14] ;
 wire \tms1x00.ins_pla_ands[8][15] ;
 wire \tms1x00.ins_pla_ands[8][1] ;
 wire \tms1x00.ins_pla_ands[8][2] ;
 wire \tms1x00.ins_pla_ands[8][3] ;
 wire \tms1x00.ins_pla_ands[8][4] ;
 wire \tms1x00.ins_pla_ands[8][5] ;
 wire \tms1x00.ins_pla_ands[8][6] ;
 wire \tms1x00.ins_pla_ands[8][7] ;
 wire \tms1x00.ins_pla_ands[8][8] ;
 wire \tms1x00.ins_pla_ands[8][9] ;
 wire \tms1x00.ins_pla_ands[9][0] ;
 wire \tms1x00.ins_pla_ands[9][10] ;
 wire \tms1x00.ins_pla_ands[9][11] ;
 wire \tms1x00.ins_pla_ands[9][12] ;
 wire \tms1x00.ins_pla_ands[9][13] ;
 wire \tms1x00.ins_pla_ands[9][14] ;
 wire \tms1x00.ins_pla_ands[9][15] ;
 wire \tms1x00.ins_pla_ands[9][1] ;
 wire \tms1x00.ins_pla_ands[9][2] ;
 wire \tms1x00.ins_pla_ands[9][3] ;
 wire \tms1x00.ins_pla_ands[9][4] ;
 wire \tms1x00.ins_pla_ands[9][5] ;
 wire \tms1x00.ins_pla_ands[9][6] ;
 wire \tms1x00.ins_pla_ands[9][7] ;
 wire \tms1x00.ins_pla_ands[9][8] ;
 wire \tms1x00.ins_pla_ands[9][9] ;
 wire \tms1x00.ins_pla_ors[0][0] ;
 wire \tms1x00.ins_pla_ors[0][10] ;
 wire \tms1x00.ins_pla_ors[0][11] ;
 wire \tms1x00.ins_pla_ors[0][12] ;
 wire \tms1x00.ins_pla_ors[0][13] ;
 wire \tms1x00.ins_pla_ors[0][14] ;
 wire \tms1x00.ins_pla_ors[0][15] ;
 wire \tms1x00.ins_pla_ors[0][16] ;
 wire \tms1x00.ins_pla_ors[0][17] ;
 wire \tms1x00.ins_pla_ors[0][18] ;
 wire \tms1x00.ins_pla_ors[0][19] ;
 wire \tms1x00.ins_pla_ors[0][1] ;
 wire \tms1x00.ins_pla_ors[0][20] ;
 wire \tms1x00.ins_pla_ors[0][21] ;
 wire \tms1x00.ins_pla_ors[0][22] ;
 wire \tms1x00.ins_pla_ors[0][23] ;
 wire \tms1x00.ins_pla_ors[0][24] ;
 wire \tms1x00.ins_pla_ors[0][25] ;
 wire \tms1x00.ins_pla_ors[0][26] ;
 wire \tms1x00.ins_pla_ors[0][27] ;
 wire \tms1x00.ins_pla_ors[0][28] ;
 wire \tms1x00.ins_pla_ors[0][29] ;
 wire \tms1x00.ins_pla_ors[0][2] ;
 wire \tms1x00.ins_pla_ors[0][3] ;
 wire \tms1x00.ins_pla_ors[0][4] ;
 wire \tms1x00.ins_pla_ors[0][5] ;
 wire \tms1x00.ins_pla_ors[0][6] ;
 wire \tms1x00.ins_pla_ors[0][7] ;
 wire \tms1x00.ins_pla_ors[0][8] ;
 wire \tms1x00.ins_pla_ors[0][9] ;
 wire \tms1x00.ins_pla_ors[10][0] ;
 wire \tms1x00.ins_pla_ors[10][10] ;
 wire \tms1x00.ins_pla_ors[10][11] ;
 wire \tms1x00.ins_pla_ors[10][12] ;
 wire \tms1x00.ins_pla_ors[10][13] ;
 wire \tms1x00.ins_pla_ors[10][14] ;
 wire \tms1x00.ins_pla_ors[10][15] ;
 wire \tms1x00.ins_pla_ors[10][16] ;
 wire \tms1x00.ins_pla_ors[10][17] ;
 wire \tms1x00.ins_pla_ors[10][18] ;
 wire \tms1x00.ins_pla_ors[10][19] ;
 wire \tms1x00.ins_pla_ors[10][1] ;
 wire \tms1x00.ins_pla_ors[10][20] ;
 wire \tms1x00.ins_pla_ors[10][21] ;
 wire \tms1x00.ins_pla_ors[10][22] ;
 wire \tms1x00.ins_pla_ors[10][23] ;
 wire \tms1x00.ins_pla_ors[10][24] ;
 wire \tms1x00.ins_pla_ors[10][25] ;
 wire \tms1x00.ins_pla_ors[10][26] ;
 wire \tms1x00.ins_pla_ors[10][27] ;
 wire \tms1x00.ins_pla_ors[10][28] ;
 wire \tms1x00.ins_pla_ors[10][29] ;
 wire \tms1x00.ins_pla_ors[10][2] ;
 wire \tms1x00.ins_pla_ors[10][3] ;
 wire \tms1x00.ins_pla_ors[10][4] ;
 wire \tms1x00.ins_pla_ors[10][5] ;
 wire \tms1x00.ins_pla_ors[10][6] ;
 wire \tms1x00.ins_pla_ors[10][7] ;
 wire \tms1x00.ins_pla_ors[10][8] ;
 wire \tms1x00.ins_pla_ors[10][9] ;
 wire \tms1x00.ins_pla_ors[11][0] ;
 wire \tms1x00.ins_pla_ors[11][10] ;
 wire \tms1x00.ins_pla_ors[11][11] ;
 wire \tms1x00.ins_pla_ors[11][12] ;
 wire \tms1x00.ins_pla_ors[11][13] ;
 wire \tms1x00.ins_pla_ors[11][14] ;
 wire \tms1x00.ins_pla_ors[11][15] ;
 wire \tms1x00.ins_pla_ors[11][16] ;
 wire \tms1x00.ins_pla_ors[11][17] ;
 wire \tms1x00.ins_pla_ors[11][18] ;
 wire \tms1x00.ins_pla_ors[11][19] ;
 wire \tms1x00.ins_pla_ors[11][1] ;
 wire \tms1x00.ins_pla_ors[11][20] ;
 wire \tms1x00.ins_pla_ors[11][21] ;
 wire \tms1x00.ins_pla_ors[11][22] ;
 wire \tms1x00.ins_pla_ors[11][23] ;
 wire \tms1x00.ins_pla_ors[11][24] ;
 wire \tms1x00.ins_pla_ors[11][25] ;
 wire \tms1x00.ins_pla_ors[11][26] ;
 wire \tms1x00.ins_pla_ors[11][27] ;
 wire \tms1x00.ins_pla_ors[11][28] ;
 wire \tms1x00.ins_pla_ors[11][29] ;
 wire \tms1x00.ins_pla_ors[11][2] ;
 wire \tms1x00.ins_pla_ors[11][3] ;
 wire \tms1x00.ins_pla_ors[11][4] ;
 wire \tms1x00.ins_pla_ors[11][5] ;
 wire \tms1x00.ins_pla_ors[11][6] ;
 wire \tms1x00.ins_pla_ors[11][7] ;
 wire \tms1x00.ins_pla_ors[11][8] ;
 wire \tms1x00.ins_pla_ors[11][9] ;
 wire \tms1x00.ins_pla_ors[12][0] ;
 wire \tms1x00.ins_pla_ors[12][10] ;
 wire \tms1x00.ins_pla_ors[12][11] ;
 wire \tms1x00.ins_pla_ors[12][12] ;
 wire \tms1x00.ins_pla_ors[12][13] ;
 wire \tms1x00.ins_pla_ors[12][14] ;
 wire \tms1x00.ins_pla_ors[12][15] ;
 wire \tms1x00.ins_pla_ors[12][16] ;
 wire \tms1x00.ins_pla_ors[12][17] ;
 wire \tms1x00.ins_pla_ors[12][18] ;
 wire \tms1x00.ins_pla_ors[12][19] ;
 wire \tms1x00.ins_pla_ors[12][1] ;
 wire \tms1x00.ins_pla_ors[12][20] ;
 wire \tms1x00.ins_pla_ors[12][21] ;
 wire \tms1x00.ins_pla_ors[12][22] ;
 wire \tms1x00.ins_pla_ors[12][23] ;
 wire \tms1x00.ins_pla_ors[12][24] ;
 wire \tms1x00.ins_pla_ors[12][25] ;
 wire \tms1x00.ins_pla_ors[12][26] ;
 wire \tms1x00.ins_pla_ors[12][27] ;
 wire \tms1x00.ins_pla_ors[12][28] ;
 wire \tms1x00.ins_pla_ors[12][29] ;
 wire \tms1x00.ins_pla_ors[12][2] ;
 wire \tms1x00.ins_pla_ors[12][3] ;
 wire \tms1x00.ins_pla_ors[12][4] ;
 wire \tms1x00.ins_pla_ors[12][5] ;
 wire \tms1x00.ins_pla_ors[12][6] ;
 wire \tms1x00.ins_pla_ors[12][7] ;
 wire \tms1x00.ins_pla_ors[12][8] ;
 wire \tms1x00.ins_pla_ors[12][9] ;
 wire \tms1x00.ins_pla_ors[13][0] ;
 wire \tms1x00.ins_pla_ors[13][10] ;
 wire \tms1x00.ins_pla_ors[13][11] ;
 wire \tms1x00.ins_pla_ors[13][12] ;
 wire \tms1x00.ins_pla_ors[13][13] ;
 wire \tms1x00.ins_pla_ors[13][14] ;
 wire \tms1x00.ins_pla_ors[13][15] ;
 wire \tms1x00.ins_pla_ors[13][16] ;
 wire \tms1x00.ins_pla_ors[13][17] ;
 wire \tms1x00.ins_pla_ors[13][18] ;
 wire \tms1x00.ins_pla_ors[13][19] ;
 wire \tms1x00.ins_pla_ors[13][1] ;
 wire \tms1x00.ins_pla_ors[13][20] ;
 wire \tms1x00.ins_pla_ors[13][21] ;
 wire \tms1x00.ins_pla_ors[13][22] ;
 wire \tms1x00.ins_pla_ors[13][23] ;
 wire \tms1x00.ins_pla_ors[13][24] ;
 wire \tms1x00.ins_pla_ors[13][25] ;
 wire \tms1x00.ins_pla_ors[13][26] ;
 wire \tms1x00.ins_pla_ors[13][27] ;
 wire \tms1x00.ins_pla_ors[13][28] ;
 wire \tms1x00.ins_pla_ors[13][29] ;
 wire \tms1x00.ins_pla_ors[13][2] ;
 wire \tms1x00.ins_pla_ors[13][3] ;
 wire \tms1x00.ins_pla_ors[13][4] ;
 wire \tms1x00.ins_pla_ors[13][5] ;
 wire \tms1x00.ins_pla_ors[13][6] ;
 wire \tms1x00.ins_pla_ors[13][7] ;
 wire \tms1x00.ins_pla_ors[13][8] ;
 wire \tms1x00.ins_pla_ors[13][9] ;
 wire \tms1x00.ins_pla_ors[14][0] ;
 wire \tms1x00.ins_pla_ors[14][10] ;
 wire \tms1x00.ins_pla_ors[14][11] ;
 wire \tms1x00.ins_pla_ors[14][12] ;
 wire \tms1x00.ins_pla_ors[14][13] ;
 wire \tms1x00.ins_pla_ors[14][14] ;
 wire \tms1x00.ins_pla_ors[14][15] ;
 wire \tms1x00.ins_pla_ors[14][16] ;
 wire \tms1x00.ins_pla_ors[14][17] ;
 wire \tms1x00.ins_pla_ors[14][18] ;
 wire \tms1x00.ins_pla_ors[14][19] ;
 wire \tms1x00.ins_pla_ors[14][1] ;
 wire \tms1x00.ins_pla_ors[14][20] ;
 wire \tms1x00.ins_pla_ors[14][21] ;
 wire \tms1x00.ins_pla_ors[14][22] ;
 wire \tms1x00.ins_pla_ors[14][23] ;
 wire \tms1x00.ins_pla_ors[14][24] ;
 wire \tms1x00.ins_pla_ors[14][25] ;
 wire \tms1x00.ins_pla_ors[14][26] ;
 wire \tms1x00.ins_pla_ors[14][27] ;
 wire \tms1x00.ins_pla_ors[14][28] ;
 wire \tms1x00.ins_pla_ors[14][29] ;
 wire \tms1x00.ins_pla_ors[14][2] ;
 wire \tms1x00.ins_pla_ors[14][3] ;
 wire \tms1x00.ins_pla_ors[14][4] ;
 wire \tms1x00.ins_pla_ors[14][5] ;
 wire \tms1x00.ins_pla_ors[14][6] ;
 wire \tms1x00.ins_pla_ors[14][7] ;
 wire \tms1x00.ins_pla_ors[14][8] ;
 wire \tms1x00.ins_pla_ors[14][9] ;
 wire \tms1x00.ins_pla_ors[15][0] ;
 wire \tms1x00.ins_pla_ors[15][10] ;
 wire \tms1x00.ins_pla_ors[15][11] ;
 wire \tms1x00.ins_pla_ors[15][12] ;
 wire \tms1x00.ins_pla_ors[15][13] ;
 wire \tms1x00.ins_pla_ors[15][14] ;
 wire \tms1x00.ins_pla_ors[15][15] ;
 wire \tms1x00.ins_pla_ors[15][16] ;
 wire \tms1x00.ins_pla_ors[15][17] ;
 wire \tms1x00.ins_pla_ors[15][18] ;
 wire \tms1x00.ins_pla_ors[15][19] ;
 wire \tms1x00.ins_pla_ors[15][1] ;
 wire \tms1x00.ins_pla_ors[15][20] ;
 wire \tms1x00.ins_pla_ors[15][21] ;
 wire \tms1x00.ins_pla_ors[15][22] ;
 wire \tms1x00.ins_pla_ors[15][23] ;
 wire \tms1x00.ins_pla_ors[15][24] ;
 wire \tms1x00.ins_pla_ors[15][25] ;
 wire \tms1x00.ins_pla_ors[15][26] ;
 wire \tms1x00.ins_pla_ors[15][27] ;
 wire \tms1x00.ins_pla_ors[15][28] ;
 wire \tms1x00.ins_pla_ors[15][29] ;
 wire \tms1x00.ins_pla_ors[15][2] ;
 wire \tms1x00.ins_pla_ors[15][3] ;
 wire \tms1x00.ins_pla_ors[15][4] ;
 wire \tms1x00.ins_pla_ors[15][5] ;
 wire \tms1x00.ins_pla_ors[15][6] ;
 wire \tms1x00.ins_pla_ors[15][7] ;
 wire \tms1x00.ins_pla_ors[15][8] ;
 wire \tms1x00.ins_pla_ors[15][9] ;
 wire \tms1x00.ins_pla_ors[1][0] ;
 wire \tms1x00.ins_pla_ors[1][10] ;
 wire \tms1x00.ins_pla_ors[1][11] ;
 wire \tms1x00.ins_pla_ors[1][12] ;
 wire \tms1x00.ins_pla_ors[1][13] ;
 wire \tms1x00.ins_pla_ors[1][14] ;
 wire \tms1x00.ins_pla_ors[1][15] ;
 wire \tms1x00.ins_pla_ors[1][16] ;
 wire \tms1x00.ins_pla_ors[1][17] ;
 wire \tms1x00.ins_pla_ors[1][18] ;
 wire \tms1x00.ins_pla_ors[1][19] ;
 wire \tms1x00.ins_pla_ors[1][1] ;
 wire \tms1x00.ins_pla_ors[1][20] ;
 wire \tms1x00.ins_pla_ors[1][21] ;
 wire \tms1x00.ins_pla_ors[1][22] ;
 wire \tms1x00.ins_pla_ors[1][23] ;
 wire \tms1x00.ins_pla_ors[1][24] ;
 wire \tms1x00.ins_pla_ors[1][25] ;
 wire \tms1x00.ins_pla_ors[1][26] ;
 wire \tms1x00.ins_pla_ors[1][27] ;
 wire \tms1x00.ins_pla_ors[1][28] ;
 wire \tms1x00.ins_pla_ors[1][29] ;
 wire \tms1x00.ins_pla_ors[1][2] ;
 wire \tms1x00.ins_pla_ors[1][3] ;
 wire \tms1x00.ins_pla_ors[1][4] ;
 wire \tms1x00.ins_pla_ors[1][5] ;
 wire \tms1x00.ins_pla_ors[1][6] ;
 wire \tms1x00.ins_pla_ors[1][7] ;
 wire \tms1x00.ins_pla_ors[1][8] ;
 wire \tms1x00.ins_pla_ors[1][9] ;
 wire \tms1x00.ins_pla_ors[2][0] ;
 wire \tms1x00.ins_pla_ors[2][10] ;
 wire \tms1x00.ins_pla_ors[2][11] ;
 wire \tms1x00.ins_pla_ors[2][12] ;
 wire \tms1x00.ins_pla_ors[2][13] ;
 wire \tms1x00.ins_pla_ors[2][14] ;
 wire \tms1x00.ins_pla_ors[2][15] ;
 wire \tms1x00.ins_pla_ors[2][16] ;
 wire \tms1x00.ins_pla_ors[2][17] ;
 wire \tms1x00.ins_pla_ors[2][18] ;
 wire \tms1x00.ins_pla_ors[2][19] ;
 wire \tms1x00.ins_pla_ors[2][1] ;
 wire \tms1x00.ins_pla_ors[2][20] ;
 wire \tms1x00.ins_pla_ors[2][21] ;
 wire \tms1x00.ins_pla_ors[2][22] ;
 wire \tms1x00.ins_pla_ors[2][23] ;
 wire \tms1x00.ins_pla_ors[2][24] ;
 wire \tms1x00.ins_pla_ors[2][25] ;
 wire \tms1x00.ins_pla_ors[2][26] ;
 wire \tms1x00.ins_pla_ors[2][27] ;
 wire \tms1x00.ins_pla_ors[2][28] ;
 wire \tms1x00.ins_pla_ors[2][29] ;
 wire \tms1x00.ins_pla_ors[2][2] ;
 wire \tms1x00.ins_pla_ors[2][3] ;
 wire \tms1x00.ins_pla_ors[2][4] ;
 wire \tms1x00.ins_pla_ors[2][5] ;
 wire \tms1x00.ins_pla_ors[2][6] ;
 wire \tms1x00.ins_pla_ors[2][7] ;
 wire \tms1x00.ins_pla_ors[2][8] ;
 wire \tms1x00.ins_pla_ors[2][9] ;
 wire \tms1x00.ins_pla_ors[3][0] ;
 wire \tms1x00.ins_pla_ors[3][10] ;
 wire \tms1x00.ins_pla_ors[3][11] ;
 wire \tms1x00.ins_pla_ors[3][12] ;
 wire \tms1x00.ins_pla_ors[3][13] ;
 wire \tms1x00.ins_pla_ors[3][14] ;
 wire \tms1x00.ins_pla_ors[3][15] ;
 wire \tms1x00.ins_pla_ors[3][16] ;
 wire \tms1x00.ins_pla_ors[3][17] ;
 wire \tms1x00.ins_pla_ors[3][18] ;
 wire \tms1x00.ins_pla_ors[3][19] ;
 wire \tms1x00.ins_pla_ors[3][1] ;
 wire \tms1x00.ins_pla_ors[3][20] ;
 wire \tms1x00.ins_pla_ors[3][21] ;
 wire \tms1x00.ins_pla_ors[3][22] ;
 wire \tms1x00.ins_pla_ors[3][23] ;
 wire \tms1x00.ins_pla_ors[3][24] ;
 wire \tms1x00.ins_pla_ors[3][25] ;
 wire \tms1x00.ins_pla_ors[3][26] ;
 wire \tms1x00.ins_pla_ors[3][27] ;
 wire \tms1x00.ins_pla_ors[3][28] ;
 wire \tms1x00.ins_pla_ors[3][29] ;
 wire \tms1x00.ins_pla_ors[3][2] ;
 wire \tms1x00.ins_pla_ors[3][3] ;
 wire \tms1x00.ins_pla_ors[3][4] ;
 wire \tms1x00.ins_pla_ors[3][5] ;
 wire \tms1x00.ins_pla_ors[3][6] ;
 wire \tms1x00.ins_pla_ors[3][7] ;
 wire \tms1x00.ins_pla_ors[3][8] ;
 wire \tms1x00.ins_pla_ors[3][9] ;
 wire \tms1x00.ins_pla_ors[4][0] ;
 wire \tms1x00.ins_pla_ors[4][10] ;
 wire \tms1x00.ins_pla_ors[4][11] ;
 wire \tms1x00.ins_pla_ors[4][12] ;
 wire \tms1x00.ins_pla_ors[4][13] ;
 wire \tms1x00.ins_pla_ors[4][14] ;
 wire \tms1x00.ins_pla_ors[4][15] ;
 wire \tms1x00.ins_pla_ors[4][16] ;
 wire \tms1x00.ins_pla_ors[4][17] ;
 wire \tms1x00.ins_pla_ors[4][18] ;
 wire \tms1x00.ins_pla_ors[4][19] ;
 wire \tms1x00.ins_pla_ors[4][1] ;
 wire \tms1x00.ins_pla_ors[4][20] ;
 wire \tms1x00.ins_pla_ors[4][21] ;
 wire \tms1x00.ins_pla_ors[4][22] ;
 wire \tms1x00.ins_pla_ors[4][23] ;
 wire \tms1x00.ins_pla_ors[4][24] ;
 wire \tms1x00.ins_pla_ors[4][25] ;
 wire \tms1x00.ins_pla_ors[4][26] ;
 wire \tms1x00.ins_pla_ors[4][27] ;
 wire \tms1x00.ins_pla_ors[4][28] ;
 wire \tms1x00.ins_pla_ors[4][29] ;
 wire \tms1x00.ins_pla_ors[4][2] ;
 wire \tms1x00.ins_pla_ors[4][3] ;
 wire \tms1x00.ins_pla_ors[4][4] ;
 wire \tms1x00.ins_pla_ors[4][5] ;
 wire \tms1x00.ins_pla_ors[4][6] ;
 wire \tms1x00.ins_pla_ors[4][7] ;
 wire \tms1x00.ins_pla_ors[4][8] ;
 wire \tms1x00.ins_pla_ors[4][9] ;
 wire \tms1x00.ins_pla_ors[5][0] ;
 wire \tms1x00.ins_pla_ors[5][10] ;
 wire \tms1x00.ins_pla_ors[5][11] ;
 wire \tms1x00.ins_pla_ors[5][12] ;
 wire \tms1x00.ins_pla_ors[5][13] ;
 wire \tms1x00.ins_pla_ors[5][14] ;
 wire \tms1x00.ins_pla_ors[5][15] ;
 wire \tms1x00.ins_pla_ors[5][16] ;
 wire \tms1x00.ins_pla_ors[5][17] ;
 wire \tms1x00.ins_pla_ors[5][18] ;
 wire \tms1x00.ins_pla_ors[5][19] ;
 wire \tms1x00.ins_pla_ors[5][1] ;
 wire \tms1x00.ins_pla_ors[5][20] ;
 wire \tms1x00.ins_pla_ors[5][21] ;
 wire \tms1x00.ins_pla_ors[5][22] ;
 wire \tms1x00.ins_pla_ors[5][23] ;
 wire \tms1x00.ins_pla_ors[5][24] ;
 wire \tms1x00.ins_pla_ors[5][25] ;
 wire \tms1x00.ins_pla_ors[5][26] ;
 wire \tms1x00.ins_pla_ors[5][27] ;
 wire \tms1x00.ins_pla_ors[5][28] ;
 wire \tms1x00.ins_pla_ors[5][29] ;
 wire \tms1x00.ins_pla_ors[5][2] ;
 wire \tms1x00.ins_pla_ors[5][3] ;
 wire \tms1x00.ins_pla_ors[5][4] ;
 wire \tms1x00.ins_pla_ors[5][5] ;
 wire \tms1x00.ins_pla_ors[5][6] ;
 wire \tms1x00.ins_pla_ors[5][7] ;
 wire \tms1x00.ins_pla_ors[5][8] ;
 wire \tms1x00.ins_pla_ors[5][9] ;
 wire \tms1x00.ins_pla_ors[6][0] ;
 wire \tms1x00.ins_pla_ors[6][10] ;
 wire \tms1x00.ins_pla_ors[6][11] ;
 wire \tms1x00.ins_pla_ors[6][12] ;
 wire \tms1x00.ins_pla_ors[6][13] ;
 wire \tms1x00.ins_pla_ors[6][14] ;
 wire \tms1x00.ins_pla_ors[6][15] ;
 wire \tms1x00.ins_pla_ors[6][16] ;
 wire \tms1x00.ins_pla_ors[6][17] ;
 wire \tms1x00.ins_pla_ors[6][18] ;
 wire \tms1x00.ins_pla_ors[6][19] ;
 wire \tms1x00.ins_pla_ors[6][1] ;
 wire \tms1x00.ins_pla_ors[6][20] ;
 wire \tms1x00.ins_pla_ors[6][21] ;
 wire \tms1x00.ins_pla_ors[6][22] ;
 wire \tms1x00.ins_pla_ors[6][23] ;
 wire \tms1x00.ins_pla_ors[6][24] ;
 wire \tms1x00.ins_pla_ors[6][25] ;
 wire \tms1x00.ins_pla_ors[6][26] ;
 wire \tms1x00.ins_pla_ors[6][27] ;
 wire \tms1x00.ins_pla_ors[6][28] ;
 wire \tms1x00.ins_pla_ors[6][29] ;
 wire \tms1x00.ins_pla_ors[6][2] ;
 wire \tms1x00.ins_pla_ors[6][3] ;
 wire \tms1x00.ins_pla_ors[6][4] ;
 wire \tms1x00.ins_pla_ors[6][5] ;
 wire \tms1x00.ins_pla_ors[6][6] ;
 wire \tms1x00.ins_pla_ors[6][7] ;
 wire \tms1x00.ins_pla_ors[6][8] ;
 wire \tms1x00.ins_pla_ors[6][9] ;
 wire \tms1x00.ins_pla_ors[7][0] ;
 wire \tms1x00.ins_pla_ors[7][10] ;
 wire \tms1x00.ins_pla_ors[7][11] ;
 wire \tms1x00.ins_pla_ors[7][12] ;
 wire \tms1x00.ins_pla_ors[7][13] ;
 wire \tms1x00.ins_pla_ors[7][14] ;
 wire \tms1x00.ins_pla_ors[7][15] ;
 wire \tms1x00.ins_pla_ors[7][16] ;
 wire \tms1x00.ins_pla_ors[7][17] ;
 wire \tms1x00.ins_pla_ors[7][18] ;
 wire \tms1x00.ins_pla_ors[7][19] ;
 wire \tms1x00.ins_pla_ors[7][1] ;
 wire \tms1x00.ins_pla_ors[7][20] ;
 wire \tms1x00.ins_pla_ors[7][21] ;
 wire \tms1x00.ins_pla_ors[7][22] ;
 wire \tms1x00.ins_pla_ors[7][23] ;
 wire \tms1x00.ins_pla_ors[7][24] ;
 wire \tms1x00.ins_pla_ors[7][25] ;
 wire \tms1x00.ins_pla_ors[7][26] ;
 wire \tms1x00.ins_pla_ors[7][27] ;
 wire \tms1x00.ins_pla_ors[7][28] ;
 wire \tms1x00.ins_pla_ors[7][29] ;
 wire \tms1x00.ins_pla_ors[7][2] ;
 wire \tms1x00.ins_pla_ors[7][3] ;
 wire \tms1x00.ins_pla_ors[7][4] ;
 wire \tms1x00.ins_pla_ors[7][5] ;
 wire \tms1x00.ins_pla_ors[7][6] ;
 wire \tms1x00.ins_pla_ors[7][7] ;
 wire \tms1x00.ins_pla_ors[7][8] ;
 wire \tms1x00.ins_pla_ors[7][9] ;
 wire \tms1x00.ins_pla_ors[8][0] ;
 wire \tms1x00.ins_pla_ors[8][10] ;
 wire \tms1x00.ins_pla_ors[8][11] ;
 wire \tms1x00.ins_pla_ors[8][12] ;
 wire \tms1x00.ins_pla_ors[8][13] ;
 wire \tms1x00.ins_pla_ors[8][14] ;
 wire \tms1x00.ins_pla_ors[8][15] ;
 wire \tms1x00.ins_pla_ors[8][16] ;
 wire \tms1x00.ins_pla_ors[8][17] ;
 wire \tms1x00.ins_pla_ors[8][18] ;
 wire \tms1x00.ins_pla_ors[8][19] ;
 wire \tms1x00.ins_pla_ors[8][1] ;
 wire \tms1x00.ins_pla_ors[8][20] ;
 wire \tms1x00.ins_pla_ors[8][21] ;
 wire \tms1x00.ins_pla_ors[8][22] ;
 wire \tms1x00.ins_pla_ors[8][23] ;
 wire \tms1x00.ins_pla_ors[8][24] ;
 wire \tms1x00.ins_pla_ors[8][25] ;
 wire \tms1x00.ins_pla_ors[8][26] ;
 wire \tms1x00.ins_pla_ors[8][27] ;
 wire \tms1x00.ins_pla_ors[8][28] ;
 wire \tms1x00.ins_pla_ors[8][29] ;
 wire \tms1x00.ins_pla_ors[8][2] ;
 wire \tms1x00.ins_pla_ors[8][3] ;
 wire \tms1x00.ins_pla_ors[8][4] ;
 wire \tms1x00.ins_pla_ors[8][5] ;
 wire \tms1x00.ins_pla_ors[8][6] ;
 wire \tms1x00.ins_pla_ors[8][7] ;
 wire \tms1x00.ins_pla_ors[8][8] ;
 wire \tms1x00.ins_pla_ors[8][9] ;
 wire \tms1x00.ins_pla_ors[9][0] ;
 wire \tms1x00.ins_pla_ors[9][10] ;
 wire \tms1x00.ins_pla_ors[9][11] ;
 wire \tms1x00.ins_pla_ors[9][12] ;
 wire \tms1x00.ins_pla_ors[9][13] ;
 wire \tms1x00.ins_pla_ors[9][14] ;
 wire \tms1x00.ins_pla_ors[9][15] ;
 wire \tms1x00.ins_pla_ors[9][16] ;
 wire \tms1x00.ins_pla_ors[9][17] ;
 wire \tms1x00.ins_pla_ors[9][18] ;
 wire \tms1x00.ins_pla_ors[9][19] ;
 wire \tms1x00.ins_pla_ors[9][1] ;
 wire \tms1x00.ins_pla_ors[9][20] ;
 wire \tms1x00.ins_pla_ors[9][21] ;
 wire \tms1x00.ins_pla_ors[9][22] ;
 wire \tms1x00.ins_pla_ors[9][23] ;
 wire \tms1x00.ins_pla_ors[9][24] ;
 wire \tms1x00.ins_pla_ors[9][25] ;
 wire \tms1x00.ins_pla_ors[9][26] ;
 wire \tms1x00.ins_pla_ors[9][27] ;
 wire \tms1x00.ins_pla_ors[9][28] ;
 wire \tms1x00.ins_pla_ors[9][29] ;
 wire \tms1x00.ins_pla_ors[9][2] ;
 wire \tms1x00.ins_pla_ors[9][3] ;
 wire \tms1x00.ins_pla_ors[9][4] ;
 wire \tms1x00.ins_pla_ors[9][5] ;
 wire \tms1x00.ins_pla_ors[9][6] ;
 wire \tms1x00.ins_pla_ors[9][7] ;
 wire \tms1x00.ins_pla_ors[9][8] ;
 wire \tms1x00.ins_pla_ors[9][9] ;
 wire \tms1x00.pla_override ;
 wire \tms1x00.rom_addr[0] ;
 wire \tms1x00.rom_addr[1] ;
 wire \tms1x00.status ;
 wire \tms1x00.wb_step ;
 wire \tms1x00.wb_step_state ;
 wire valid;
 wire wb_rst_override;
 wire \wbs_o_buff[0] ;
 wire \wbs_o_buff[10] ;
 wire \wbs_o_buff[11] ;
 wire \wbs_o_buff[12] ;
 wire \wbs_o_buff[13] ;
 wire \wbs_o_buff[14] ;
 wire \wbs_o_buff[15] ;
 wire \wbs_o_buff[16] ;
 wire \wbs_o_buff[17] ;
 wire \wbs_o_buff[18] ;
 wire \wbs_o_buff[19] ;
 wire \wbs_o_buff[1] ;
 wire \wbs_o_buff[20] ;
 wire \wbs_o_buff[21] ;
 wire \wbs_o_buff[22] ;
 wire \wbs_o_buff[23] ;
 wire \wbs_o_buff[24] ;
 wire \wbs_o_buff[25] ;
 wire \wbs_o_buff[26] ;
 wire \wbs_o_buff[27] ;
 wire \wbs_o_buff[28] ;
 wire \wbs_o_buff[29] ;
 wire \wbs_o_buff[2] ;
 wire \wbs_o_buff[30] ;
 wire \wbs_o_buff[31] ;
 wire \wbs_o_buff[3] ;
 wire \wbs_o_buff[4] ;
 wire \wbs_o_buff[5] ;
 wire \wbs_o_buff[6] ;
 wire \wbs_o_buff[7] ;
 wire \wbs_o_buff[8] ;
 wire \wbs_o_buff[9] ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_01763_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_02228_));
 sky130_fd_sc_hd__diode_2 ANTENNA_100 (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_101 (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA_102 (.DIODE(net594));
 sky130_fd_sc_hd__diode_2 ANTENNA_103 (.DIODE(net594));
 sky130_fd_sc_hd__diode_2 ANTENNA_104 (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA_105 (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA_106 (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_107 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_108 (.DIODE(net755));
 sky130_fd_sc_hd__diode_2 ANTENNA_109 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_02230_));
 sky130_fd_sc_hd__diode_2 ANTENNA_110 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_111 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_112 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_113 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_114 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_115 (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_116 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_117 (.DIODE(net893));
 sky130_fd_sc_hd__diode_2 ANTENNA_118 (.DIODE(net904));
 sky130_fd_sc_hd__diode_2 ANTENNA_119 (.DIODE(net943));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_02231_));
 sky130_fd_sc_hd__diode_2 ANTENNA_120 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_121 (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_122 (.DIODE(net958));
 sky130_fd_sc_hd__diode_2 ANTENNA_123 (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_124 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_125 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_126 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_127 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_128 (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_129 (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_02459_));
 sky130_fd_sc_hd__diode_2 ANTENNA_130 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_131 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_132 (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA_133 (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_134 (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_135 (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA_136 (.DIODE(net1066));
 sky130_fd_sc_hd__diode_2 ANTENNA_137 (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_138 (.DIODE(_01674_));
 sky130_fd_sc_hd__diode_2 ANTENNA_139 (.DIODE(_01718_));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_02490_));
 sky130_fd_sc_hd__diode_2 ANTENNA_140 (.DIODE(_01951_));
 sky130_fd_sc_hd__diode_2 ANTENNA_141 (.DIODE(_01973_));
 sky130_fd_sc_hd__diode_2 ANTENNA_142 (.DIODE(_01973_));
 sky130_fd_sc_hd__diode_2 ANTENNA_143 (.DIODE(_01984_));
 sky130_fd_sc_hd__diode_2 ANTENNA_144 (.DIODE(_02224_));
 sky130_fd_sc_hd__diode_2 ANTENNA_145 (.DIODE(_02231_));
 sky130_fd_sc_hd__diode_2 ANTENNA_146 (.DIODE(_02400_));
 sky130_fd_sc_hd__diode_2 ANTENNA_147 (.DIODE(_02437_));
 sky130_fd_sc_hd__diode_2 ANTENNA_148 (.DIODE(_02452_));
 sky130_fd_sc_hd__diode_2 ANTENNA_149 (.DIODE(_02564_));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_02636_));
 sky130_fd_sc_hd__diode_2 ANTENNA_150 (.DIODE(_03260_));
 sky130_fd_sc_hd__diode_2 ANTENNA_151 (.DIODE(_03356_));
 sky130_fd_sc_hd__diode_2 ANTENNA_152 (.DIODE(_03457_));
 sky130_fd_sc_hd__diode_2 ANTENNA_153 (.DIODE(_03457_));
 sky130_fd_sc_hd__diode_2 ANTENNA_154 (.DIODE(_03457_));
 sky130_fd_sc_hd__diode_2 ANTENNA_155 (.DIODE(_03485_));
 sky130_fd_sc_hd__diode_2 ANTENNA_156 (.DIODE(_03485_));
 sky130_fd_sc_hd__diode_2 ANTENNA_157 (.DIODE(_04002_));
 sky130_fd_sc_hd__diode_2 ANTENNA_158 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_159 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(_02688_));
 sky130_fd_sc_hd__diode_2 ANTENNA_160 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_161 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_162 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_163 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_164 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_165 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_166 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_167 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_168 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_169 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(_02693_));
 sky130_fd_sc_hd__diode_2 ANTENNA_170 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_171 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_172 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA_173 (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA_174 (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA_175 (.DIODE(net738));
 sky130_fd_sc_hd__diode_2 ANTENNA_176 (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_177 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_178 (.DIODE(net761));
 sky130_fd_sc_hd__diode_2 ANTENNA_179 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(_02869_));
 sky130_fd_sc_hd__diode_2 ANTENNA_180 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_181 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_182 (.DIODE(net876));
 sky130_fd_sc_hd__diode_2 ANTENNA_183 (.DIODE(net934));
 sky130_fd_sc_hd__diode_2 ANTENNA_184 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_185 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_186 (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_187 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_188 (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_189 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(_02915_));
 sky130_fd_sc_hd__diode_2 ANTENNA_190 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_191 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_192 (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_193 (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_194 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_195 (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA_196 (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_197 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_198 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_199 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_01798_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(_03039_));
 sky130_fd_sc_hd__diode_2 ANTENNA_200 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_201 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_202 (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_203 (.DIODE(_01940_));
 sky130_fd_sc_hd__diode_2 ANTENNA_204 (.DIODE(_01940_));
 sky130_fd_sc_hd__diode_2 ANTENNA_205 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_206 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_207 (.DIODE(net849));
 sky130_fd_sc_hd__diode_2 ANTENNA_208 (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(_03049_));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(_03123_));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(_03234_));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(_03321_));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(_03321_));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(_03357_));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(_03429_));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(_03429_));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(_03429_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_01798_));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(_03434_));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(_03439_));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(_03439_));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(_03574_));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(_04090_));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(_04167_));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(_04532_));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(_04848_));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(\tms1x00.CA ));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(\tms1x00.ins_pla_ors[9][23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_01852_));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(\wbs_o_buff[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_01896_));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_01918_));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_01918_));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_02228_));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_89 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_02228_));
 sky130_fd_sc_hd__diode_2 ANTENNA_90 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_91 (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_92 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_93 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_94 (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_95 (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_96 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA_97 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA_98 (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA_99 (.DIODE(net436));
 sky130_fd_sc_hd__decap_6 FILLER_0_1002 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1073 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1228 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_855 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1090 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1125 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1225 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1279 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1297 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1328 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1349 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1353 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1359 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1385 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1020 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1101 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1139 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1152 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1251 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1262 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1286 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1297 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1304 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1324 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1336 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1363 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1375 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1383 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_690 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1080 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1172 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1214 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1297 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1356 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1368 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_891 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_916 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1036 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1106 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1139 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1196 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1215 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1257 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1267 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_1285 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1305 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1356 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1368 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1380 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_704 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_963 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_974 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1066 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1226 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1235 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1247 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1287 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1294 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1317 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1348 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1360 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1377 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1384 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_887 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_904 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1023 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1092 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1101 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_1201 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1220 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1287 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1304 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1328 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1340 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_971 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1221 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1272 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_1280 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1288 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1349 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1353 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_992 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1030 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1092 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1152 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1164 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1257 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1265 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1299 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1316 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1326 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_1335 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1343 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1358 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1382 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_871 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1030 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1160 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1223 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_1235 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1269 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_1281 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1300 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1312 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_1317 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1325 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1355 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1048 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1080 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1108 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1132 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1271 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1287 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1297 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1308 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1320 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1369 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_926 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1172 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1188 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1242 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1103 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1114 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1142 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1164 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1179 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1215 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1240 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1283 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1295 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1303 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1315 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1335 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1347 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1359 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1385 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_771 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1094 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1135 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1218 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1254 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1267 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1286 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1297 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1307 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1327 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1339 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1356 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1368 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1380 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_871 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1055 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1120 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1173 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_1212 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1220 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1237 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1246 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1270 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_1282 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1290 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1301 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1353 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_799 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1050 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1086 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1104 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1139 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1151 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1163 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1270 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1282 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1289 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1322 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1352 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1364 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_1376 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1384 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1153 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1171 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_1183 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_1215 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_1279 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1287 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1305 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1385 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_882 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_954 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1027 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1084 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1199 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1268 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1307 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1328 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1357 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1369 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1384 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_812 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_863 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_875 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_915 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_927 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_971 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1064 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1167 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1178 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1190 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1236 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_1248 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1293 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_1305 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_674 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_880 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1195 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1277 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_998 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1087 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1163 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1172 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1186 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1202 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1238 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1261 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1296 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1308 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1365 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1385 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_955 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1075 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1142 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1152 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1206 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1228 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1239 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1265 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1297 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1309 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1321 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1333 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1385 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_971 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1247 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1271 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_870 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_995 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1104 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1180 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1223 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1232 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_1240 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1293 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1305 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1385 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_718 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1040 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1083 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1152 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1262 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1274 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1308 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1320 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1332 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1385 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_704 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_970 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1163 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_1172 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1247 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1261 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1279 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1298 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1310 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_935 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_956 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1042 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1132 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1199 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1260 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1272 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1385 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_647 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_815 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1013 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1178 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1187 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1200 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1292 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1304 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_723 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_887 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1134 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1168 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1231 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1267 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1369 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1377 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1384 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1106 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1167 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1236 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_619 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_723 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_860 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_882 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_900 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1207 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1263 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_871 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_915 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_971 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1012 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1163 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1179 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1385 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1154 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1243 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1267 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_532 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_758 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1014 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1052 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1104 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1116 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1168 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1180 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1216 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1228 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1371 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1377 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1384 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_850 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_882 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_891 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_943 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_970 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1179 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1187 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1234 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1023 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1058 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1076 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1140 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1168 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1243 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1267 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1337 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1369 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1243 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1285 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1365 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1385 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_999 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1151 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1243 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1267 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1385 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_759 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_823 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_880 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_959 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1024 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_831 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_885 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_959 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1036 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1377 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1384 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_639 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_759 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1019 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1027 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1071 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1079 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1131 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1155 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1228 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1251 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1263 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1269 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1301 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_816 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_874 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1377 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1384 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1167 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1176 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1226 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1238 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1242 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1252 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1283 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1292 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1304 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1353 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1385 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_899 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1377 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1384 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1241 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1256 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1268 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1289 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1294 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1304 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1328 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1334 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1357 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1364 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1385 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1029 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1042 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1168 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1190 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1226 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1253 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1265 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1056 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1171 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1192 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1215 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1235 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1244 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1254 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1292 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1304 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1365 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1385 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_616 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1125 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1209 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1242 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1250 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1267 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1275 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1066 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1080 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1163 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1191 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1236 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1248 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1310 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1385 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_835 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_935 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_954 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1024 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1083 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1103 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1156 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1202 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1244 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1256 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1262 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1270 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1299 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1324 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1336 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1385 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_859 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_926 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_985 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1166 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_807 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_827 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_964 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1059 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1153 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1212 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1254 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1276 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1294 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1304 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1324 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1336 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1348 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1360 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1385 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_675 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_907 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_955 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_999 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1098 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1153 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1187 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1267 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1369 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1385 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_690 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_812 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_927 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1050 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1104 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1116 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1268 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1301 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1317 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1328 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1334 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1356 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1368 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1377 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1384 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_779 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_964 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_994 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1052 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1248 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1269 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1289 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1301 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1316 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1324 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1342 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1353 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1363 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1375 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_1383 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_756 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_930 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1125 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1191 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1270 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1279 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1297 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1338 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1350 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_730 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1000 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1056 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1139 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1175 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1204 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1262 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1289 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1324 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1336 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1366 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1378 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_814 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_962 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1018 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1059 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1180 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1213 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_1225 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1236 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1240 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1261 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1297 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1315 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1328 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1337 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1385 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_674 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1174 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1251 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1260 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1268 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1296 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1308 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1327 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1364 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1376 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1384 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_932 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1159 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1171 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1179 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1215 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1227 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1239 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1281 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1293 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1305 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1324 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1332 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1354 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1360 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1366 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1385 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_992 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_1061 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1097 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1286 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1312 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_1324 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1336 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1353 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1359 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_648 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_826 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_970 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1048 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_1361 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1366 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1377 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1384 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1014 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1123 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1140 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1179 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1270 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1279 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1291 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1313 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1340 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1352 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1385 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_992 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1040 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1087 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1095 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1156 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1195 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1260 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1299 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1324 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1333 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1362 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1371 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_1383 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1050 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1060 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1068 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1120 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1174 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_1186 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1218 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1281 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1299 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1315 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1335 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1348 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1352 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1385 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_945 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_952 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_958 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1183 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1240 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1262 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1321 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1333 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1364 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1376 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1384 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_816 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_966 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1084 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1126 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_1134 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1159 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1238 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1296 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1348 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1356 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_619 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_688 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1079 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1104 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1140 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1264 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1276 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1321 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1330 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1374 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_908 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1192 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1222 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1234 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1271 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1282 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1294 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1301 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1314 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1317 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1325 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1343 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1355 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1364 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1385 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_504 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1086 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1231 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1243 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1270 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1274 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1299 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_1307 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1318 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1330 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1345 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1376 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1384 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1171 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1212 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1239 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1258 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1261 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_1269 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1292 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1312 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1335 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1344 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_1352 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1357 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1368 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1373 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1380 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_618 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1266 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1278 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1284 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1289 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_1297 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1309 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1318 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_1330 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1342 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1345 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_1353 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1372 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1384 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_758 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_906 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1104 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1188 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1285 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_1293 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1349 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1353 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1364 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1385 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_618 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_878 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_886 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_938 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1125 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1142 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1210 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1220 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1263 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1289 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1309 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1321 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1333 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1076 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1190 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1258 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1265 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1274 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1282 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1299 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1317 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1333 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1344 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1355 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1364 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_887 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1110 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_1173 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1224 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1242 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1263 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1267 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1289 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1297 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1303 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1342 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1358 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1384 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_919 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1103 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1122 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1180 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1247 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1256 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1265 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1271 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_1279 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1287 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1300 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1338 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1366 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1385 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1050 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1097 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1197 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1215 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1231 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1267 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1286 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1297 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1315 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1327 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1335 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1342 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1382 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_940 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1162 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1174 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1186 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1200 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1227 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_1281 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1300 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_1341 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1366 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1019 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1230 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1239 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1248 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1265 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1295 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1307 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1328 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1336 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1342 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1353 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1374 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_929 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1022 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1030 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1114 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1124 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1191 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1238 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1270 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1282 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1288 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1294 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1324 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_1332 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1351 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1364 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1384 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_784 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_968 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1022 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1096 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1139 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1150 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1156 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1164 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1245 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1268 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1280 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1289 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_1297 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1320 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1332 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1336 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1356 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1360 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_926 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_938 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_975 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1022 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_999 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1032 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1167 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1178 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1202 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1240 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1261 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1284 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1296 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1304 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1335 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1343 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1361 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1385 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1148 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1162 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1260 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1264 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1286 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1295 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1301 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1309 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1328 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1340 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1362 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1374 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_805 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_818 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1104 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1122 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1218 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1270 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1274 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1278 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1295 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1329 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1341 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1349 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1385 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_823 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_899 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_990 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_998 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1026 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1058 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1197 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1270 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1319 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1331 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1338 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1345 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1350 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1361 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1384 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1044 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1120 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1123 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1135 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1238 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_1285 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1293 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1305 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_1313 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1317 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_1325 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1348 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1361 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1385 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_665 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_883 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_999 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1031 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1132 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1230 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1239 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1296 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1316 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1324 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1342 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1345 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1353 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1372 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1384 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_702 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_815 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1124 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1144 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1163 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1227 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1239 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1272 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1280 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1298 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1304 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1335 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1343 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1349 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1360 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1385 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_891 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_944 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1132 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1199 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1210 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1246 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1266 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1299 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_1307 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1327 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1339 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1372 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1384 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1048 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1153 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1170 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_1178 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1239 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1248 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1271 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1283 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1300 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_1337 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1349 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1385 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_616 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_844 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_860 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_907 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1039 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1131 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1200 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1208 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1251 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1266 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1289 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1296 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1302 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1319 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1331 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1354 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1358 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_871 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_969 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1042 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_702 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_855 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1055 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1214 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1218 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1242 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1284 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1304 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1359 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1385 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_665 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1015 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1038 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1092 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1188 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1219 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1253 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1265 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1286 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1297 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1311 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1323 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1335 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1385 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_646 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_910 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_1169 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1222 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1232 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1261 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1268 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1274 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1280 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1292 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1304 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1317 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_1325 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1337 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1346 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1358 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1385 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1082 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1268 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1280 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1313 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1325 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1363 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_1375 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1384 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_622 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_855 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_975 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1024 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1050 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1088 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1123 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1192 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1234 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1281 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1315 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1321 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1355 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_450 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_672 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_784 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_875 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_910 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1029 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1079 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1142 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1151 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1200 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1265 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1285 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1298 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1310 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1316 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1324 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1331 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1343 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1345 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1353 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1364 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1376 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1384 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_639 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_886 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1032 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1124 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1232 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1250 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1277 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1305 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1335 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1353 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_891 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1000 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1188 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1218 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1269 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1300 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1312 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1319 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1339 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1345 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1375 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_1383 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_695 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_805 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_924 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1125 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1159 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1183 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1225 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1234 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1238 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1272 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1284 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1302 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1312 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1321 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1331 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1351 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1385 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_844 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_900 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_957 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1075 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1199 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_1207 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1296 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1385 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_892 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_942 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1079 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1026 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1167 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1268 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1282 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1294 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1300 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1310 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1385 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_840 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1135 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1195 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1204 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1210 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1216 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1228 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1313 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1327 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1339 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1385 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1228 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_1240 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1248 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1288 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1300 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1312 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1335 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1347 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1359 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_1086 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1188 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1215 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1268 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1280 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1385 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_824 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_975 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1086 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1106 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1110 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1122 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1168 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1371 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1377 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1384 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1039 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1385 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_647 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_928 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_974 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1135 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1038 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1184 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1267 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_420 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_532 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_874 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1000 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1070 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1220 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_1228 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1240 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1280 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1292 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1304 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1385 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_896 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_940 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_957 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1036 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1051 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1086 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1098 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1207 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1266 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1357 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_907 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1039 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_824 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1076 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1136 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1176 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1211 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1309 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1100 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1215 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1245 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1263 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1272 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_760 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_816 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_851 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1068 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1110 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1126 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1159 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1240 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1279 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1291 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1385 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_939 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_968 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1026 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1038 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1215 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1253 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1313 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1385 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_812 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_940 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1055 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1104 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1160 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1296 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1308 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1323 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1352 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1364 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1377 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1384 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_972 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1164 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1187 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_1199 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1207 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1245 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1299 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1311 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1323 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_1335 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_939 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_995 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1055 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1159 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1171 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1202 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1219 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1268 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1276 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1287 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1365 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1385 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_991 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1263 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1275 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1311 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_704 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_812 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_883 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_927 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1012 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1058 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1270 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1282 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1294 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1298 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1315 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1336 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1348 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1360 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1385 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_663 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_843 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1094 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1250 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1262 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1272 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1318 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1327 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1339 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1385 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_820 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1044 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1056 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1079 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_1201 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1215 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1238 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1287 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1294 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1324 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1337 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1349 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1361 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_796 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_827 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_956 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1101 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1197 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1240 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1252 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1269 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1280 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1356 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1368 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1380 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_818 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_871 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_974 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1051 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1159 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1172 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1192 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1239 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1270 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1281 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1293 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1300 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1306 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_1313 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1317 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1333 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1355 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1385 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_955 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1208 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1212 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1256 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1262 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1270 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1282 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1293 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1310 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1322 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1352 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1364 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1376 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1384 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1003 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1103 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1160 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1216 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1274 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1293 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1303 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1352 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1364 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1377 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1384 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_956 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1019 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1041 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1094 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1198 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1248 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1287 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1305 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1325 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1333 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1340 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1363 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1375 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_1383 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_926 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_970 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1156 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1176 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_1201 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1238 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1297 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1324 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1328 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1349 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1385 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_1173 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1240 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1252 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1276 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1289 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1356 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1023 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1047 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_1059 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1071 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1146 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1176 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1238 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1258 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1285 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1297 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1301 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1310 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1329 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1341 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1358 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_875 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_990 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1027 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1052 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1128 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1207 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1249 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1257 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1270 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1282 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1298 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1318 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1330 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1342 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1345 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1353 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1371 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_1383 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_644 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_918 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1039 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_814 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_826 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_864 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_994 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__inv_2 _05072_ (.A(net651),
    .Y(_01614_));
 sky130_fd_sc_hd__inv_2 _05073_ (.A(\tms1x00.PC[4] ),
    .Y(_01615_));
 sky130_fd_sc_hd__inv_2 _05074_ (.A(\tms1x00.CL ),
    .Y(_01616_));
 sky130_fd_sc_hd__clkinv_2 _05075_ (.A(\tms1x00.O_latch[4] ),
    .Y(_01617_));
 sky130_fd_sc_hd__inv_2 _05076_ (.A(net660),
    .Y(_01618_));
 sky130_fd_sc_hd__clkinv_2 _05077_ (.A(net661),
    .Y(_01619_));
 sky130_fd_sc_hd__clkinv_2 _05078_ (.A(net664),
    .Y(_01620_));
 sky130_fd_sc_hd__inv_2 _05079_ (.A(net665),
    .Y(_01621_));
 sky130_fd_sc_hd__clkinv_2 _05080_ (.A(\tms1x00.cycle[0] ),
    .Y(_01622_));
 sky130_fd_sc_hd__inv_2 _05081_ (.A(net668),
    .Y(_01623_));
 sky130_fd_sc_hd__clkinv_4 _05082_ (.A(net672),
    .Y(_01624_));
 sky130_fd_sc_hd__inv_6 _05083_ (.A(net679),
    .Y(_01625_));
 sky130_fd_sc_hd__clkinv_4 _05084_ (.A(net681),
    .Y(_01626_));
 sky130_fd_sc_hd__inv_4 _05085_ (.A(net690),
    .Y(_01627_));
 sky130_fd_sc_hd__clkinv_2 _05086_ (.A(net693),
    .Y(_01628_));
 sky130_fd_sc_hd__inv_6 _05087_ (.A(net698),
    .Y(_01629_));
 sky130_fd_sc_hd__inv_4 _05088_ (.A(net701),
    .Y(_01630_));
 sky130_fd_sc_hd__inv_2 _05089_ (.A(\tms1x00.ins_pla_ands[0][15] ),
    .Y(_01631_));
 sky130_fd_sc_hd__inv_2 _05090_ (.A(\tms1x00.ins_pla_ands[1][15] ),
    .Y(_01632_));
 sky130_fd_sc_hd__clkinv_2 _05091_ (.A(net989),
    .Y(_01633_));
 sky130_fd_sc_hd__inv_2 _05092_ (.A(net994),
    .Y(_01634_));
 sky130_fd_sc_hd__inv_6 _05093_ (.A(net74),
    .Y(_01635_));
 sky130_fd_sc_hd__inv_12 _05094_ (.A(net119),
    .Y(net178));
 sky130_fd_sc_hd__inv_2 _05095_ (.A(net985),
    .Y(_01636_));
 sky130_fd_sc_hd__inv_8 _05096_ (.A(net984),
    .Y(_01637_));
 sky130_fd_sc_hd__clkinv_4 _05097_ (.A(net705),
    .Y(_01638_));
 sky130_fd_sc_hd__inv_2 _05098_ (.A(\tms1x00.rom_addr[0] ),
    .Y(_01639_));
 sky130_fd_sc_hd__inv_2 _05099_ (.A(\tms1x00.rom_addr[1] ),
    .Y(_01640_));
 sky130_fd_sc_hd__nor2_1 _05100_ (.A(wb_rst_override),
    .B(net74),
    .Y(_01641_));
 sky130_fd_sc_hd__inv_2 _05101_ (.A(net631),
    .Y(net167));
 sky130_fd_sc_hd__and2_4 _05102_ (.A(net118),
    .B(net87),
    .X(valid));
 sky130_fd_sc_hd__mux2_1 _05103_ (.A0(\tms1x00.ins_pla_ands[24][1] ),
    .A1(\tms1x00.ins_pla_ands[24][0] ),
    .S(net700),
    .X(_01642_));
 sky130_fd_sc_hd__mux2_1 _05104_ (.A0(\tms1x00.ins_pla_ands[24][7] ),
    .A1(\tms1x00.ins_pla_ands[24][6] ),
    .S(net687),
    .X(_01643_));
 sky130_fd_sc_hd__mux2_1 _05105_ (.A0(\tms1x00.ins_pla_ands[24][5] ),
    .A1(\tms1x00.ins_pla_ands[24][4] ),
    .S(net691),
    .X(_01644_));
 sky130_fd_sc_hd__mux2_1 _05106_ (.A0(\tms1x00.ins_pla_ands[24][9] ),
    .A1(\tms1x00.ins_pla_ands[24][8] ),
    .S(net683),
    .X(_01645_));
 sky130_fd_sc_hd__or4_4 _05107_ (.A(_01642_),
    .B(_01643_),
    .C(_01644_),
    .D(_01645_),
    .X(_01646_));
 sky130_fd_sc_hd__mux2_1 _05108_ (.A0(\tms1x00.ins_pla_ands[24][3] ),
    .A1(\tms1x00.ins_pla_ands[24][2] ),
    .S(net697),
    .X(_01647_));
 sky130_fd_sc_hd__mux2_1 _05109_ (.A0(\tms1x00.ins_pla_ands[24][13] ),
    .A1(\tms1x00.ins_pla_ands[24][12] ),
    .S(net673),
    .X(_01648_));
 sky130_fd_sc_hd__mux2_1 _05110_ (.A0(\tms1x00.ins_pla_ands[24][11] ),
    .A1(\tms1x00.ins_pla_ands[24][10] ),
    .S(net678),
    .X(_01649_));
 sky130_fd_sc_hd__mux2_1 _05111_ (.A0(\tms1x00.ins_pla_ands[24][15] ),
    .A1(\tms1x00.ins_pla_ands[24][14] ),
    .S(net669),
    .X(_01650_));
 sky130_fd_sc_hd__or4_4 _05112_ (.A(_01647_),
    .B(_01648_),
    .C(_01649_),
    .D(_01650_),
    .X(_01651_));
 sky130_fd_sc_hd__nor2_8 _05113_ (.A(_01646_),
    .B(_01651_),
    .Y(_01652_));
 sky130_fd_sc_hd__mux2_1 _05114_ (.A0(\tms1x00.ins_pla_ands[26][11] ),
    .A1(\tms1x00.ins_pla_ands[26][10] ),
    .S(net677),
    .X(_01653_));
 sky130_fd_sc_hd__mux2_1 _05115_ (.A0(\tms1x00.ins_pla_ands[26][7] ),
    .A1(\tms1x00.ins_pla_ands[26][6] ),
    .S(net687),
    .X(_01654_));
 sky130_fd_sc_hd__mux2_1 _05116_ (.A0(\tms1x00.ins_pla_ands[26][3] ),
    .A1(\tms1x00.ins_pla_ands[26][2] ),
    .S(net696),
    .X(_01655_));
 sky130_fd_sc_hd__mux2_1 _05117_ (.A0(\tms1x00.ins_pla_ands[26][5] ),
    .A1(\tms1x00.ins_pla_ands[26][4] ),
    .S(net691),
    .X(_01656_));
 sky130_fd_sc_hd__or4_4 _05118_ (.A(_01653_),
    .B(_01654_),
    .C(_01655_),
    .D(_01656_),
    .X(_01657_));
 sky130_fd_sc_hd__mux2_1 _05119_ (.A0(\tms1x00.ins_pla_ands[26][1] ),
    .A1(\tms1x00.ins_pla_ands[26][0] ),
    .S(net704),
    .X(_01658_));
 sky130_fd_sc_hd__mux2_1 _05120_ (.A0(\tms1x00.ins_pla_ands[26][13] ),
    .A1(\tms1x00.ins_pla_ands[26][12] ),
    .S(net675),
    .X(_01659_));
 sky130_fd_sc_hd__mux2_1 _05121_ (.A0(\tms1x00.ins_pla_ands[26][15] ),
    .A1(\tms1x00.ins_pla_ands[26][14] ),
    .S(net667),
    .X(_01660_));
 sky130_fd_sc_hd__mux2_1 _05122_ (.A0(\tms1x00.ins_pla_ands[26][9] ),
    .A1(\tms1x00.ins_pla_ands[26][8] ),
    .S(net685),
    .X(_01661_));
 sky130_fd_sc_hd__or4_2 _05123_ (.A(_01658_),
    .B(_01659_),
    .C(_01660_),
    .D(_01661_),
    .X(_01662_));
 sky130_fd_sc_hd__nor2_4 _05124_ (.A(_01657_),
    .B(_01662_),
    .Y(_01663_));
 sky130_fd_sc_hd__mux2_1 _05125_ (.A0(\tms1x00.ins_pla_ands[20][11] ),
    .A1(\tms1x00.ins_pla_ands[20][10] ),
    .S(net678),
    .X(_01664_));
 sky130_fd_sc_hd__mux2_1 _05126_ (.A0(\tms1x00.ins_pla_ands[20][7] ),
    .A1(\tms1x00.ins_pla_ands[20][6] ),
    .S(net687),
    .X(_01665_));
 sky130_fd_sc_hd__mux2_1 _05127_ (.A0(\tms1x00.ins_pla_ands[20][3] ),
    .A1(\tms1x00.ins_pla_ands[20][2] ),
    .S(net696),
    .X(_01666_));
 sky130_fd_sc_hd__mux2_1 _05128_ (.A0(\tms1x00.ins_pla_ands[20][5] ),
    .A1(\tms1x00.ins_pla_ands[20][4] ),
    .S(net691),
    .X(_01667_));
 sky130_fd_sc_hd__or4_4 _05129_ (.A(_01664_),
    .B(_01665_),
    .C(_01666_),
    .D(_01667_),
    .X(_01668_));
 sky130_fd_sc_hd__mux2_1 _05130_ (.A0(\tms1x00.ins_pla_ands[20][1] ),
    .A1(\tms1x00.ins_pla_ands[20][0] ),
    .S(net700),
    .X(_01669_));
 sky130_fd_sc_hd__mux2_1 _05131_ (.A0(\tms1x00.ins_pla_ands[20][13] ),
    .A1(\tms1x00.ins_pla_ands[20][12] ),
    .S(net673),
    .X(_01670_));
 sky130_fd_sc_hd__mux2_1 _05132_ (.A0(\tms1x00.ins_pla_ands[20][15] ),
    .A1(\tms1x00.ins_pla_ands[20][14] ),
    .S(net667),
    .X(_01671_));
 sky130_fd_sc_hd__mux2_1 _05133_ (.A0(\tms1x00.ins_pla_ands[20][9] ),
    .A1(\tms1x00.ins_pla_ands[20][8] ),
    .S(net683),
    .X(_01672_));
 sky130_fd_sc_hd__or4_4 _05134_ (.A(_01669_),
    .B(_01670_),
    .C(_01671_),
    .D(_01672_),
    .X(_01673_));
 sky130_fd_sc_hd__nor2_8 _05135_ (.A(_01668_),
    .B(_01673_),
    .Y(_01674_));
 sky130_fd_sc_hd__mux2_1 _05136_ (.A0(\tms1x00.ins_pla_ands[7][11] ),
    .A1(\tms1x00.ins_pla_ands[7][10] ),
    .S(net680),
    .X(_01675_));
 sky130_fd_sc_hd__mux2_1 _05137_ (.A0(\tms1x00.ins_pla_ands[7][7] ),
    .A1(\tms1x00.ins_pla_ands[7][6] ),
    .S(net689),
    .X(_01676_));
 sky130_fd_sc_hd__mux2_1 _05138_ (.A0(\tms1x00.ins_pla_ands[7][3] ),
    .A1(\tms1x00.ins_pla_ands[7][2] ),
    .S(net698),
    .X(_01677_));
 sky130_fd_sc_hd__mux2_1 _05139_ (.A0(\tms1x00.ins_pla_ands[7][5] ),
    .A1(\tms1x00.ins_pla_ands[7][4] ),
    .S(net694),
    .X(_01678_));
 sky130_fd_sc_hd__or4_4 _05140_ (.A(_01675_),
    .B(_01676_),
    .C(_01677_),
    .D(_01678_),
    .X(_01679_));
 sky130_fd_sc_hd__mux2_1 _05141_ (.A0(\tms1x00.ins_pla_ands[7][1] ),
    .A1(\tms1x00.ins_pla_ands[7][0] ),
    .S(net703),
    .X(_01680_));
 sky130_fd_sc_hd__mux2_1 _05142_ (.A0(\tms1x00.ins_pla_ands[7][13] ),
    .A1(\tms1x00.ins_pla_ands[7][12] ),
    .S(net674),
    .X(_01681_));
 sky130_fd_sc_hd__mux2_1 _05143_ (.A0(\tms1x00.ins_pla_ands[7][15] ),
    .A1(\tms1x00.ins_pla_ands[7][14] ),
    .S(net670),
    .X(_01682_));
 sky130_fd_sc_hd__mux2_1 _05144_ (.A0(\tms1x00.ins_pla_ands[7][9] ),
    .A1(\tms1x00.ins_pla_ands[7][8] ),
    .S(net684),
    .X(_01683_));
 sky130_fd_sc_hd__or4_4 _05145_ (.A(_01680_),
    .B(_01681_),
    .C(_01682_),
    .D(_01683_),
    .X(_01684_));
 sky130_fd_sc_hd__nor2_8 _05146_ (.A(_01679_),
    .B(_01684_),
    .Y(_01685_));
 sky130_fd_sc_hd__mux2_1 _05147_ (.A0(\tms1x00.ins_pla_ands[11][11] ),
    .A1(\tms1x00.ins_pla_ands[11][10] ),
    .S(net679),
    .X(_01686_));
 sky130_fd_sc_hd__mux2_1 _05148_ (.A0(\tms1x00.ins_pla_ands[11][7] ),
    .A1(\tms1x00.ins_pla_ands[11][6] ),
    .S(net686),
    .X(_01687_));
 sky130_fd_sc_hd__mux2_1 _05149_ (.A0(\tms1x00.ins_pla_ands[11][3] ),
    .A1(\tms1x00.ins_pla_ands[11][2] ),
    .S(net697),
    .X(_01688_));
 sky130_fd_sc_hd__mux2_1 _05150_ (.A0(\tms1x00.ins_pla_ands[11][5] ),
    .A1(\tms1x00.ins_pla_ands[11][4] ),
    .S(net692),
    .X(_01689_));
 sky130_fd_sc_hd__or4_4 _05151_ (.A(_01686_),
    .B(_01687_),
    .C(_01688_),
    .D(_01689_),
    .X(_01690_));
 sky130_fd_sc_hd__mux2_1 _05152_ (.A0(\tms1x00.ins_pla_ands[11][1] ),
    .A1(\tms1x00.ins_pla_ands[11][0] ),
    .S(net701),
    .X(_01691_));
 sky130_fd_sc_hd__mux2_1 _05153_ (.A0(\tms1x00.ins_pla_ands[11][13] ),
    .A1(\tms1x00.ins_pla_ands[11][12] ),
    .S(net672),
    .X(_01692_));
 sky130_fd_sc_hd__mux2_1 _05154_ (.A0(\tms1x00.ins_pla_ands[11][15] ),
    .A1(\tms1x00.ins_pla_ands[11][14] ),
    .S(net668),
    .X(_01693_));
 sky130_fd_sc_hd__mux2_1 _05155_ (.A0(\tms1x00.ins_pla_ands[11][9] ),
    .A1(\tms1x00.ins_pla_ands[11][8] ),
    .S(net681),
    .X(_01694_));
 sky130_fd_sc_hd__or4_4 _05156_ (.A(_01691_),
    .B(_01692_),
    .C(_01693_),
    .D(_01694_),
    .X(_01695_));
 sky130_fd_sc_hd__nor2_8 _05157_ (.A(_01690_),
    .B(_01695_),
    .Y(_01696_));
 sky130_fd_sc_hd__mux2_1 _05158_ (.A0(\tms1x00.ins_pla_ands[28][7] ),
    .A1(\tms1x00.ins_pla_ands[28][6] ),
    .S(net687),
    .X(_01697_));
 sky130_fd_sc_hd__mux2_1 _05159_ (.A0(\tms1x00.ins_pla_ands[28][15] ),
    .A1(\tms1x00.ins_pla_ands[28][14] ),
    .S(net667),
    .X(_01698_));
 sky130_fd_sc_hd__mux2_1 _05160_ (.A0(\tms1x00.ins_pla_ands[28][13] ),
    .A1(\tms1x00.ins_pla_ands[28][12] ),
    .S(net673),
    .X(_01699_));
 sky130_fd_sc_hd__mux2_1 _05161_ (.A0(\tms1x00.ins_pla_ands[28][3] ),
    .A1(\tms1x00.ins_pla_ands[28][2] ),
    .S(net697),
    .X(_01700_));
 sky130_fd_sc_hd__or4_2 _05162_ (.A(_01697_),
    .B(_01698_),
    .C(_01699_),
    .D(_01700_),
    .X(_01701_));
 sky130_fd_sc_hd__mux2_1 _05163_ (.A0(\tms1x00.ins_pla_ands[28][1] ),
    .A1(\tms1x00.ins_pla_ands[28][0] ),
    .S(net700),
    .X(_01702_));
 sky130_fd_sc_hd__mux2_1 _05164_ (.A0(\tms1x00.ins_pla_ands[28][9] ),
    .A1(\tms1x00.ins_pla_ands[28][8] ),
    .S(net683),
    .X(_01703_));
 sky130_fd_sc_hd__mux2_1 _05165_ (.A0(\tms1x00.ins_pla_ands[28][5] ),
    .A1(\tms1x00.ins_pla_ands[28][4] ),
    .S(net691),
    .X(_01704_));
 sky130_fd_sc_hd__mux2_1 _05166_ (.A0(\tms1x00.ins_pla_ands[28][11] ),
    .A1(\tms1x00.ins_pla_ands[28][10] ),
    .S(net677),
    .X(_01705_));
 sky130_fd_sc_hd__or4_1 _05167_ (.A(_01702_),
    .B(_01703_),
    .C(_01704_),
    .D(_01705_),
    .X(_01706_));
 sky130_fd_sc_hd__nor2_2 _05168_ (.A(_01701_),
    .B(_01706_),
    .Y(_01707_));
 sky130_fd_sc_hd__mux2_1 _05169_ (.A0(\tms1x00.ins_pla_ands[16][5] ),
    .A1(\tms1x00.ins_pla_ands[16][4] ),
    .S(net691),
    .X(_01708_));
 sky130_fd_sc_hd__mux2_1 _05170_ (.A0(\tms1x00.ins_pla_ands[16][7] ),
    .A1(\tms1x00.ins_pla_ands[16][6] ),
    .S(net690),
    .X(_01709_));
 sky130_fd_sc_hd__mux2_1 _05171_ (.A0(\tms1x00.ins_pla_ands[16][13] ),
    .A1(\tms1x00.ins_pla_ands[16][12] ),
    .S(net676),
    .X(_01710_));
 sky130_fd_sc_hd__mux2_2 _05172_ (.A0(\tms1x00.ins_pla_ands[16][15] ),
    .A1(\tms1x00.ins_pla_ands[16][14] ),
    .S(net668),
    .X(_01711_));
 sky130_fd_sc_hd__mux2_1 _05173_ (.A0(\tms1x00.ins_pla_ands[16][11] ),
    .A1(\tms1x00.ins_pla_ands[16][10] ),
    .S(net678),
    .X(_01712_));
 sky130_fd_sc_hd__mux2_1 _05174_ (.A0(\tms1x00.ins_pla_ands[16][9] ),
    .A1(\tms1x00.ins_pla_ands[16][8] ),
    .S(net681),
    .X(_01713_));
 sky130_fd_sc_hd__mux2_1 _05175_ (.A0(\tms1x00.ins_pla_ands[16][3] ),
    .A1(\tms1x00.ins_pla_ands[16][2] ),
    .S(net696),
    .X(_01714_));
 sky130_fd_sc_hd__or4_4 _05176_ (.A(_01708_),
    .B(_01709_),
    .C(_01713_),
    .D(_01714_),
    .X(_01715_));
 sky130_fd_sc_hd__mux2_1 _05177_ (.A0(\tms1x00.ins_pla_ands[16][1] ),
    .A1(\tms1x00.ins_pla_ands[16][0] ),
    .S(net701),
    .X(_01716_));
 sky130_fd_sc_hd__or4_4 _05178_ (.A(_01710_),
    .B(_01711_),
    .C(_01712_),
    .D(_01716_),
    .X(_01717_));
 sky130_fd_sc_hd__nor2_8 _05179_ (.A(_01715_),
    .B(_01717_),
    .Y(_01718_));
 sky130_fd_sc_hd__mux2_1 _05180_ (.A0(\tms1x00.ins_pla_ands[4][11] ),
    .A1(\tms1x00.ins_pla_ands[4][10] ),
    .S(net680),
    .X(_01719_));
 sky130_fd_sc_hd__mux2_1 _05181_ (.A0(\tms1x00.ins_pla_ands[4][7] ),
    .A1(\tms1x00.ins_pla_ands[4][6] ),
    .S(net688),
    .X(_01720_));
 sky130_fd_sc_hd__mux2_1 _05182_ (.A0(\tms1x00.ins_pla_ands[4][3] ),
    .A1(\tms1x00.ins_pla_ands[4][2] ),
    .S(net698),
    .X(_01721_));
 sky130_fd_sc_hd__mux2_1 _05183_ (.A0(\tms1x00.ins_pla_ands[4][5] ),
    .A1(\tms1x00.ins_pla_ands[4][4] ),
    .S(net693),
    .X(_01722_));
 sky130_fd_sc_hd__or4_2 _05184_ (.A(_01719_),
    .B(_01720_),
    .C(_01721_),
    .D(_01722_),
    .X(_01723_));
 sky130_fd_sc_hd__mux2_1 _05185_ (.A0(\tms1x00.ins_pla_ands[4][1] ),
    .A1(\tms1x00.ins_pla_ands[4][0] ),
    .S(net702),
    .X(_01724_));
 sky130_fd_sc_hd__mux2_1 _05186_ (.A0(\tms1x00.ins_pla_ands[4][13] ),
    .A1(\tms1x00.ins_pla_ands[4][12] ),
    .S(net674),
    .X(_01725_));
 sky130_fd_sc_hd__mux2_1 _05187_ (.A0(\tms1x00.ins_pla_ands[4][15] ),
    .A1(\tms1x00.ins_pla_ands[4][14] ),
    .S(net670),
    .X(_01726_));
 sky130_fd_sc_hd__mux2_1 _05188_ (.A0(\tms1x00.ins_pla_ands[4][9] ),
    .A1(\tms1x00.ins_pla_ands[4][8] ),
    .S(net684),
    .X(_01727_));
 sky130_fd_sc_hd__or4_4 _05189_ (.A(_01724_),
    .B(_01725_),
    .C(_01726_),
    .D(_01727_),
    .X(_01728_));
 sky130_fd_sc_hd__nor2_4 _05190_ (.A(_01723_),
    .B(_01728_),
    .Y(_01729_));
 sky130_fd_sc_hd__and2_1 _05191_ (.A(net680),
    .B(\tms1x00.ins_pla_ands[0][10] ),
    .X(_01730_));
 sky130_fd_sc_hd__mux2_1 _05192_ (.A0(\tms1x00.ins_pla_ands[0][5] ),
    .A1(\tms1x00.ins_pla_ands[0][4] ),
    .S(net694),
    .X(_01731_));
 sky130_fd_sc_hd__mux2_1 _05193_ (.A0(\tms1x00.ins_pla_ands[0][9] ),
    .A1(\tms1x00.ins_pla_ands[0][8] ),
    .S(net684),
    .X(_01732_));
 sky130_fd_sc_hd__and2b_1 _05194_ (.A_N(net674),
    .B(\tms1x00.ins_pla_ands[0][13] ),
    .X(_01733_));
 sky130_fd_sc_hd__and2_1 _05195_ (.A(net698),
    .B(\tms1x00.ins_pla_ands[0][2] ),
    .X(_01734_));
 sky130_fd_sc_hd__mux2_1 _05196_ (.A0(\tms1x00.ins_pla_ands[0][7] ),
    .A1(\tms1x00.ins_pla_ands[0][6] ),
    .S(net689),
    .X(_01735_));
 sky130_fd_sc_hd__nand2b_1 _05197_ (.A_N(net703),
    .B(\tms1x00.ins_pla_ands[0][1] ),
    .Y(_01736_));
 sky130_fd_sc_hd__nand2_1 _05198_ (.A(net703),
    .B(\tms1x00.ins_pla_ands[0][0] ),
    .Y(_01737_));
 sky130_fd_sc_hd__a2111o_1 _05199_ (.A1(_01629_),
    .A2(\tms1x00.ins_pla_ands[0][3] ),
    .B1(_01730_),
    .C1(_01733_),
    .D1(_01734_),
    .X(_01738_));
 sky130_fd_sc_hd__nand2_1 _05200_ (.A(net670),
    .B(\tms1x00.ins_pla_ands[0][14] ),
    .Y(_01739_));
 sky130_fd_sc_hd__o2111a_1 _05201_ (.A1(net670),
    .A2(_01631_),
    .B1(_01736_),
    .C1(_01737_),
    .D1(_01739_),
    .X(_01740_));
 sky130_fd_sc_hd__a221oi_2 _05202_ (.A1(net674),
    .A2(\tms1x00.ins_pla_ands[0][12] ),
    .B1(\tms1x00.ins_pla_ands[0][11] ),
    .B2(_01625_),
    .C1(_01735_),
    .Y(_01741_));
 sky130_fd_sc_hd__nor2_1 _05203_ (.A(_01731_),
    .B(_01732_),
    .Y(_01742_));
 sky130_fd_sc_hd__and4b_4 _05204_ (.A_N(_01738_),
    .B(_01740_),
    .C(_01741_),
    .D(_01742_),
    .X(_01743_));
 sky130_fd_sc_hd__mux2_1 _05205_ (.A0(\tms1x00.ins_pla_ands[2][3] ),
    .A1(\tms1x00.ins_pla_ands[2][2] ),
    .S(net698),
    .X(_01744_));
 sky130_fd_sc_hd__a221o_2 _05206_ (.A1(_01630_),
    .A2(\tms1x00.ins_pla_ands[2][1] ),
    .B1(\tms1x00.ins_pla_ands[2][7] ),
    .B2(_01627_),
    .C1(_01744_),
    .X(_01745_));
 sky130_fd_sc_hd__mux2_2 _05207_ (.A0(\tms1x00.ins_pla_ands[2][11] ),
    .A1(\tms1x00.ins_pla_ands[2][10] ),
    .S(net680),
    .X(_01746_));
 sky130_fd_sc_hd__mux2_2 _05208_ (.A0(\tms1x00.ins_pla_ands[2][13] ),
    .A1(\tms1x00.ins_pla_ands[2][12] ),
    .S(net674),
    .X(_01747_));
 sky130_fd_sc_hd__a22o_1 _05209_ (.A1(net688),
    .A2(\tms1x00.ins_pla_ands[2][6] ),
    .B1(\tms1x00.ins_pla_ands[2][0] ),
    .B2(net702),
    .X(_01748_));
 sky130_fd_sc_hd__mux2_1 _05210_ (.A0(\tms1x00.ins_pla_ands[2][9] ),
    .A1(\tms1x00.ins_pla_ands[2][8] ),
    .S(net684),
    .X(_01749_));
 sky130_fd_sc_hd__mux2_1 _05211_ (.A0(\tms1x00.ins_pla_ands[2][5] ),
    .A1(\tms1x00.ins_pla_ands[2][4] ),
    .S(net693),
    .X(_01750_));
 sky130_fd_sc_hd__mux2_1 _05212_ (.A0(\tms1x00.ins_pla_ands[2][15] ),
    .A1(\tms1x00.ins_pla_ands[2][14] ),
    .S(net670),
    .X(_01751_));
 sky130_fd_sc_hd__or4_2 _05213_ (.A(_01748_),
    .B(_01749_),
    .C(_01750_),
    .D(_01751_),
    .X(_01752_));
 sky130_fd_sc_hd__nor4_4 _05214_ (.A(_01745_),
    .B(_01746_),
    .C(_01747_),
    .D(_01752_),
    .Y(_01753_));
 sky130_fd_sc_hd__mux2_1 _05215_ (.A0(\tms1x00.ins_pla_ands[13][11] ),
    .A1(\tms1x00.ins_pla_ands[13][10] ),
    .S(net679),
    .X(_01754_));
 sky130_fd_sc_hd__a221o_2 _05216_ (.A1(net686),
    .A2(\tms1x00.ins_pla_ands[13][6] ),
    .B1(\tms1x00.ins_pla_ands[13][9] ),
    .B2(_01626_),
    .C1(_01754_),
    .X(_01755_));
 sky130_fd_sc_hd__mux2_1 _05217_ (.A0(\tms1x00.ins_pla_ands[13][13] ),
    .A1(\tms1x00.ins_pla_ands[13][12] ),
    .S(net672),
    .X(_01756_));
 sky130_fd_sc_hd__mux2_1 _05218_ (.A0(\tms1x00.ins_pla_ands[13][3] ),
    .A1(\tms1x00.ins_pla_ands[13][2] ),
    .S(\tms1x00.B[0] ),
    .X(_01757_));
 sky130_fd_sc_hd__a22o_2 _05219_ (.A1(_01623_),
    .A2(\tms1x00.ins_pla_ands[13][15] ),
    .B1(\tms1x00.ins_pla_ands[13][8] ),
    .B2(net681),
    .X(_01758_));
 sky130_fd_sc_hd__a22o_1 _05220_ (.A1(_01627_),
    .A2(\tms1x00.ins_pla_ands[13][7] ),
    .B1(\tms1x00.ins_pla_ands[13][14] ),
    .B2(net669),
    .X(_01759_));
 sky130_fd_sc_hd__mux2_1 _05221_ (.A0(\tms1x00.ins_pla_ands[13][5] ),
    .A1(\tms1x00.ins_pla_ands[13][4] ),
    .S(\tms1x00.ins_arg[5] ),
    .X(_01760_));
 sky130_fd_sc_hd__mux2_1 _05222_ (.A0(\tms1x00.ins_pla_ands[13][1] ),
    .A1(\tms1x00.ins_pla_ands[13][0] ),
    .S(net701),
    .X(_01761_));
 sky130_fd_sc_hd__or4_2 _05223_ (.A(_01756_),
    .B(_01757_),
    .C(_01760_),
    .D(_01761_),
    .X(_01762_));
 sky130_fd_sc_hd__nor4_4 _05224_ (.A(_01755_),
    .B(_01758_),
    .C(_01759_),
    .D(_01762_),
    .Y(_01763_));
 sky130_fd_sc_hd__and2_1 _05225_ (.A(net680),
    .B(\tms1x00.ins_pla_ands[1][10] ),
    .X(_01764_));
 sky130_fd_sc_hd__mux2_1 _05226_ (.A0(\tms1x00.ins_pla_ands[1][5] ),
    .A1(\tms1x00.ins_pla_ands[1][4] ),
    .S(net694),
    .X(_01765_));
 sky130_fd_sc_hd__mux2_1 _05227_ (.A0(\tms1x00.ins_pla_ands[1][9] ),
    .A1(\tms1x00.ins_pla_ands[1][8] ),
    .S(net685),
    .X(_01766_));
 sky130_fd_sc_hd__and2b_1 _05228_ (.A_N(net674),
    .B(\tms1x00.ins_pla_ands[1][13] ),
    .X(_01767_));
 sky130_fd_sc_hd__and2_1 _05229_ (.A(net699),
    .B(\tms1x00.ins_pla_ands[1][2] ),
    .X(_01768_));
 sky130_fd_sc_hd__mux2_1 _05230_ (.A0(\tms1x00.ins_pla_ands[1][7] ),
    .A1(\tms1x00.ins_pla_ands[1][6] ),
    .S(net689),
    .X(_01769_));
 sky130_fd_sc_hd__nand2b_1 _05231_ (.A_N(net703),
    .B(\tms1x00.ins_pla_ands[1][1] ),
    .Y(_01770_));
 sky130_fd_sc_hd__nand2_1 _05232_ (.A(net703),
    .B(\tms1x00.ins_pla_ands[1][0] ),
    .Y(_01771_));
 sky130_fd_sc_hd__a2111o_1 _05233_ (.A1(_01629_),
    .A2(\tms1x00.ins_pla_ands[1][3] ),
    .B1(_01764_),
    .C1(_01767_),
    .D1(_01768_),
    .X(_01772_));
 sky130_fd_sc_hd__nand2_1 _05234_ (.A(net670),
    .B(\tms1x00.ins_pla_ands[1][14] ),
    .Y(_01773_));
 sky130_fd_sc_hd__o2111a_1 _05235_ (.A1(net670),
    .A2(_01632_),
    .B1(_01770_),
    .C1(_01771_),
    .D1(_01773_),
    .X(_01774_));
 sky130_fd_sc_hd__a221oi_2 _05236_ (.A1(net674),
    .A2(\tms1x00.ins_pla_ands[1][12] ),
    .B1(\tms1x00.ins_pla_ands[1][11] ),
    .B2(_01625_),
    .C1(_01769_),
    .Y(_01775_));
 sky130_fd_sc_hd__nor2_1 _05237_ (.A(_01765_),
    .B(_01766_),
    .Y(_01776_));
 sky130_fd_sc_hd__and4b_4 _05238_ (.A_N(_01772_),
    .B(_01774_),
    .C(_01775_),
    .D(_01776_),
    .X(_01777_));
 sky130_fd_sc_hd__mux2_1 _05239_ (.A0(\tms1x00.ins_pla_ands[3][3] ),
    .A1(\tms1x00.ins_pla_ands[3][2] ),
    .S(net698),
    .X(_01778_));
 sky130_fd_sc_hd__a221o_2 _05240_ (.A1(_01627_),
    .A2(\tms1x00.ins_pla_ands[3][7] ),
    .B1(\tms1x00.ins_pla_ands[3][1] ),
    .B2(_01630_),
    .C1(_01778_),
    .X(_01779_));
 sky130_fd_sc_hd__mux2_2 _05241_ (.A0(\tms1x00.ins_pla_ands[3][11] ),
    .A1(\tms1x00.ins_pla_ands[3][10] ),
    .S(net680),
    .X(_01780_));
 sky130_fd_sc_hd__mux2_2 _05242_ (.A0(\tms1x00.ins_pla_ands[3][13] ),
    .A1(\tms1x00.ins_pla_ands[3][12] ),
    .S(net674),
    .X(_01781_));
 sky130_fd_sc_hd__a22o_1 _05243_ (.A1(net702),
    .A2(\tms1x00.ins_pla_ands[3][0] ),
    .B1(\tms1x00.ins_pla_ands[3][6] ),
    .B2(net689),
    .X(_01782_));
 sky130_fd_sc_hd__mux2_1 _05244_ (.A0(\tms1x00.ins_pla_ands[3][9] ),
    .A1(\tms1x00.ins_pla_ands[3][8] ),
    .S(net684),
    .X(_01783_));
 sky130_fd_sc_hd__mux2_1 _05245_ (.A0(\tms1x00.ins_pla_ands[3][5] ),
    .A1(\tms1x00.ins_pla_ands[3][4] ),
    .S(net693),
    .X(_01784_));
 sky130_fd_sc_hd__mux2_1 _05246_ (.A0(\tms1x00.ins_pla_ands[3][15] ),
    .A1(\tms1x00.ins_pla_ands[3][14] ),
    .S(net671),
    .X(_01785_));
 sky130_fd_sc_hd__or4_2 _05247_ (.A(_01782_),
    .B(_01783_),
    .C(_01784_),
    .D(_01785_),
    .X(_01786_));
 sky130_fd_sc_hd__nor4_4 _05248_ (.A(_01779_),
    .B(_01780_),
    .C(_01781_),
    .D(_01786_),
    .Y(_01787_));
 sky130_fd_sc_hd__mux2_1 _05249_ (.A0(\tms1x00.ins_pla_ands[18][1] ),
    .A1(\tms1x00.ins_pla_ands[18][0] ),
    .S(net704),
    .X(_01788_));
 sky130_fd_sc_hd__mux2_1 _05250_ (.A0(\tms1x00.ins_pla_ands[18][7] ),
    .A1(\tms1x00.ins_pla_ands[18][6] ),
    .S(net689),
    .X(_01789_));
 sky130_fd_sc_hd__mux2_1 _05251_ (.A0(\tms1x00.ins_pla_ands[18][5] ),
    .A1(\tms1x00.ins_pla_ands[18][4] ),
    .S(net695),
    .X(_01790_));
 sky130_fd_sc_hd__mux2_2 _05252_ (.A0(\tms1x00.ins_pla_ands[18][9] ),
    .A1(\tms1x00.ins_pla_ands[18][8] ),
    .S(net681),
    .X(_01791_));
 sky130_fd_sc_hd__or4_4 _05253_ (.A(_01788_),
    .B(_01789_),
    .C(_01790_),
    .D(_01791_),
    .X(_01792_));
 sky130_fd_sc_hd__mux2_1 _05254_ (.A0(\tms1x00.ins_pla_ands[18][11] ),
    .A1(\tms1x00.ins_pla_ands[18][10] ),
    .S(net677),
    .X(_01793_));
 sky130_fd_sc_hd__mux2_1 _05255_ (.A0(\tms1x00.ins_pla_ands[18][13] ),
    .A1(\tms1x00.ins_pla_ands[18][12] ),
    .S(net673),
    .X(_01794_));
 sky130_fd_sc_hd__mux2_1 _05256_ (.A0(\tms1x00.ins_pla_ands[18][3] ),
    .A1(\tms1x00.ins_pla_ands[18][2] ),
    .S(net697),
    .X(_01795_));
 sky130_fd_sc_hd__mux2_2 _05257_ (.A0(\tms1x00.ins_pla_ands[18][15] ),
    .A1(\tms1x00.ins_pla_ands[18][14] ),
    .S(net667),
    .X(_01796_));
 sky130_fd_sc_hd__or4_4 _05258_ (.A(_01793_),
    .B(_01794_),
    .C(_01795_),
    .D(_01796_),
    .X(_01797_));
 sky130_fd_sc_hd__nor2_8 _05259_ (.A(_01792_),
    .B(_01797_),
    .Y(_01798_));
 sky130_fd_sc_hd__mux2_1 _05260_ (.A0(\tms1x00.ins_pla_ands[29][7] ),
    .A1(\tms1x00.ins_pla_ands[29][6] ),
    .S(net687),
    .X(_01799_));
 sky130_fd_sc_hd__mux2_1 _05261_ (.A0(\tms1x00.ins_pla_ands[29][15] ),
    .A1(\tms1x00.ins_pla_ands[29][14] ),
    .S(net667),
    .X(_01800_));
 sky130_fd_sc_hd__mux2_1 _05262_ (.A0(\tms1x00.ins_pla_ands[29][13] ),
    .A1(\tms1x00.ins_pla_ands[29][12] ),
    .S(net673),
    .X(_01801_));
 sky130_fd_sc_hd__mux2_1 _05263_ (.A0(\tms1x00.ins_pla_ands[29][3] ),
    .A1(\tms1x00.ins_pla_ands[29][2] ),
    .S(net696),
    .X(_01802_));
 sky130_fd_sc_hd__or4_1 _05264_ (.A(_01799_),
    .B(_01800_),
    .C(_01801_),
    .D(_01802_),
    .X(_01803_));
 sky130_fd_sc_hd__mux2_1 _05265_ (.A0(\tms1x00.ins_pla_ands[29][1] ),
    .A1(\tms1x00.ins_pla_ands[29][0] ),
    .S(net700),
    .X(_01804_));
 sky130_fd_sc_hd__mux2_1 _05266_ (.A0(\tms1x00.ins_pla_ands[29][9] ),
    .A1(\tms1x00.ins_pla_ands[29][8] ),
    .S(net683),
    .X(_01805_));
 sky130_fd_sc_hd__mux2_1 _05267_ (.A0(\tms1x00.ins_pla_ands[29][5] ),
    .A1(\tms1x00.ins_pla_ands[29][4] ),
    .S(net691),
    .X(_01806_));
 sky130_fd_sc_hd__mux2_1 _05268_ (.A0(\tms1x00.ins_pla_ands[29][11] ),
    .A1(\tms1x00.ins_pla_ands[29][10] ),
    .S(net677),
    .X(_01807_));
 sky130_fd_sc_hd__or4_1 _05269_ (.A(_01804_),
    .B(_01805_),
    .C(_01806_),
    .D(_01807_),
    .X(_01808_));
 sky130_fd_sc_hd__nor2_2 _05270_ (.A(_01803_),
    .B(_01808_),
    .Y(_01809_));
 sky130_fd_sc_hd__mux2_1 _05271_ (.A0(\tms1x00.ins_pla_ands[23][11] ),
    .A1(\tms1x00.ins_pla_ands[23][10] ),
    .S(net677),
    .X(_01810_));
 sky130_fd_sc_hd__mux2_1 _05272_ (.A0(\tms1x00.ins_pla_ands[23][7] ),
    .A1(\tms1x00.ins_pla_ands[23][6] ),
    .S(net687),
    .X(_01811_));
 sky130_fd_sc_hd__mux2_1 _05273_ (.A0(\tms1x00.ins_pla_ands[23][3] ),
    .A1(\tms1x00.ins_pla_ands[23][2] ),
    .S(net699),
    .X(_01812_));
 sky130_fd_sc_hd__mux2_1 _05274_ (.A0(\tms1x00.ins_pla_ands[23][5] ),
    .A1(\tms1x00.ins_pla_ands[23][4] ),
    .S(net692),
    .X(_01813_));
 sky130_fd_sc_hd__or4_4 _05275_ (.A(_01810_),
    .B(_01811_),
    .C(_01812_),
    .D(_01813_),
    .X(_01814_));
 sky130_fd_sc_hd__mux2_1 _05276_ (.A0(\tms1x00.ins_pla_ands[23][1] ),
    .A1(\tms1x00.ins_pla_ands[23][0] ),
    .S(net700),
    .X(_01815_));
 sky130_fd_sc_hd__mux2_1 _05277_ (.A0(\tms1x00.ins_pla_ands[23][13] ),
    .A1(\tms1x00.ins_pla_ands[23][12] ),
    .S(net673),
    .X(_01816_));
 sky130_fd_sc_hd__mux2_1 _05278_ (.A0(\tms1x00.ins_pla_ands[23][15] ),
    .A1(\tms1x00.ins_pla_ands[23][14] ),
    .S(net667),
    .X(_01817_));
 sky130_fd_sc_hd__mux2_1 _05279_ (.A0(\tms1x00.ins_pla_ands[23][9] ),
    .A1(\tms1x00.ins_pla_ands[23][8] ),
    .S(net683),
    .X(_01818_));
 sky130_fd_sc_hd__or4_4 _05280_ (.A(_01815_),
    .B(_01816_),
    .C(_01817_),
    .D(_01818_),
    .X(_01819_));
 sky130_fd_sc_hd__nor2_8 _05281_ (.A(_01814_),
    .B(_01819_),
    .Y(_01820_));
 sky130_fd_sc_hd__mux2_1 _05282_ (.A0(\tms1x00.ins_pla_ands[12][11] ),
    .A1(\tms1x00.ins_pla_ands[12][10] ),
    .S(net679),
    .X(_01821_));
 sky130_fd_sc_hd__a221o_2 _05283_ (.A1(net686),
    .A2(\tms1x00.ins_pla_ands[12][6] ),
    .B1(\tms1x00.ins_pla_ands[12][9] ),
    .B2(_01626_),
    .C1(_01821_),
    .X(_01822_));
 sky130_fd_sc_hd__mux2_1 _05284_ (.A0(\tms1x00.ins_pla_ands[12][13] ),
    .A1(\tms1x00.ins_pla_ands[12][12] ),
    .S(net672),
    .X(_01823_));
 sky130_fd_sc_hd__mux2_1 _05285_ (.A0(\tms1x00.ins_pla_ands[12][3] ),
    .A1(\tms1x00.ins_pla_ands[12][2] ),
    .S(net697),
    .X(_01824_));
 sky130_fd_sc_hd__a22o_2 _05286_ (.A1(_01623_),
    .A2(\tms1x00.ins_pla_ands[12][15] ),
    .B1(\tms1x00.ins_pla_ands[12][8] ),
    .B2(net681),
    .X(_01825_));
 sky130_fd_sc_hd__a22o_1 _05287_ (.A1(_01627_),
    .A2(\tms1x00.ins_pla_ands[12][7] ),
    .B1(\tms1x00.ins_pla_ands[12][14] ),
    .B2(net668),
    .X(_01826_));
 sky130_fd_sc_hd__mux2_1 _05288_ (.A0(\tms1x00.ins_pla_ands[12][5] ),
    .A1(\tms1x00.ins_pla_ands[12][4] ),
    .S(net692),
    .X(_01827_));
 sky130_fd_sc_hd__mux2_1 _05289_ (.A0(\tms1x00.ins_pla_ands[12][1] ),
    .A1(\tms1x00.ins_pla_ands[12][0] ),
    .S(\tms1x00.B[1] ),
    .X(_01828_));
 sky130_fd_sc_hd__or4_2 _05290_ (.A(_01823_),
    .B(_01824_),
    .C(_01827_),
    .D(_01828_),
    .X(_01829_));
 sky130_fd_sc_hd__nor4_4 _05291_ (.A(_01822_),
    .B(_01825_),
    .C(_01826_),
    .D(_01829_),
    .Y(_01830_));
 sky130_fd_sc_hd__mux2_1 _05292_ (.A0(\tms1x00.ins_pla_ands[27][11] ),
    .A1(\tms1x00.ins_pla_ands[27][10] ),
    .S(net677),
    .X(_01831_));
 sky130_fd_sc_hd__mux2_1 _05293_ (.A0(\tms1x00.ins_pla_ands[27][7] ),
    .A1(\tms1x00.ins_pla_ands[27][6] ),
    .S(net687),
    .X(_01832_));
 sky130_fd_sc_hd__mux2_1 _05294_ (.A0(\tms1x00.ins_pla_ands[27][3] ),
    .A1(\tms1x00.ins_pla_ands[27][2] ),
    .S(net696),
    .X(_01833_));
 sky130_fd_sc_hd__mux2_1 _05295_ (.A0(\tms1x00.ins_pla_ands[27][5] ),
    .A1(\tms1x00.ins_pla_ands[27][4] ),
    .S(net691),
    .X(_01834_));
 sky130_fd_sc_hd__or4_4 _05296_ (.A(_01831_),
    .B(_01832_),
    .C(_01833_),
    .D(_01834_),
    .X(_01835_));
 sky130_fd_sc_hd__mux2_1 _05297_ (.A0(\tms1x00.ins_pla_ands[27][1] ),
    .A1(\tms1x00.ins_pla_ands[27][0] ),
    .S(net704),
    .X(_01836_));
 sky130_fd_sc_hd__mux2_1 _05298_ (.A0(\tms1x00.ins_pla_ands[27][13] ),
    .A1(\tms1x00.ins_pla_ands[27][12] ),
    .S(net675),
    .X(_01837_));
 sky130_fd_sc_hd__mux2_1 _05299_ (.A0(\tms1x00.ins_pla_ands[27][15] ),
    .A1(\tms1x00.ins_pla_ands[27][14] ),
    .S(net671),
    .X(_01838_));
 sky130_fd_sc_hd__mux2_1 _05300_ (.A0(\tms1x00.ins_pla_ands[27][9] ),
    .A1(\tms1x00.ins_pla_ands[27][8] ),
    .S(net685),
    .X(_01839_));
 sky130_fd_sc_hd__or4_2 _05301_ (.A(_01836_),
    .B(_01837_),
    .C(_01838_),
    .D(_01839_),
    .X(_01840_));
 sky130_fd_sc_hd__nor2_4 _05302_ (.A(_01835_),
    .B(_01840_),
    .Y(_01841_));
 sky130_fd_sc_hd__mux2_1 _05303_ (.A0(\tms1x00.ins_pla_ands[10][11] ),
    .A1(\tms1x00.ins_pla_ands[10][10] ),
    .S(net680),
    .X(_01842_));
 sky130_fd_sc_hd__mux2_1 _05304_ (.A0(\tms1x00.ins_pla_ands[10][7] ),
    .A1(\tms1x00.ins_pla_ands[10][6] ),
    .S(net690),
    .X(_01843_));
 sky130_fd_sc_hd__mux2_1 _05305_ (.A0(\tms1x00.ins_pla_ands[10][3] ),
    .A1(\tms1x00.ins_pla_ands[10][2] ),
    .S(\tms1x00.B[0] ),
    .X(_01844_));
 sky130_fd_sc_hd__mux2_1 _05306_ (.A0(\tms1x00.ins_pla_ands[10][5] ),
    .A1(\tms1x00.ins_pla_ands[10][4] ),
    .S(net692),
    .X(_01845_));
 sky130_fd_sc_hd__or4_4 _05307_ (.A(_01842_),
    .B(_01843_),
    .C(_01844_),
    .D(_01845_),
    .X(_01846_));
 sky130_fd_sc_hd__mux2_1 _05308_ (.A0(\tms1x00.ins_pla_ands[10][1] ),
    .A1(\tms1x00.ins_pla_ands[10][0] ),
    .S(\tms1x00.B[1] ),
    .X(_01847_));
 sky130_fd_sc_hd__mux2_1 _05309_ (.A0(\tms1x00.ins_pla_ands[10][13] ),
    .A1(\tms1x00.ins_pla_ands[10][12] ),
    .S(net672),
    .X(_01848_));
 sky130_fd_sc_hd__mux2_1 _05310_ (.A0(\tms1x00.ins_pla_ands[10][15] ),
    .A1(\tms1x00.ins_pla_ands[10][14] ),
    .S(net668),
    .X(_01849_));
 sky130_fd_sc_hd__mux2_1 _05311_ (.A0(\tms1x00.ins_pla_ands[10][9] ),
    .A1(\tms1x00.ins_pla_ands[10][8] ),
    .S(net681),
    .X(_01850_));
 sky130_fd_sc_hd__or4_4 _05312_ (.A(_01847_),
    .B(_01848_),
    .C(_01849_),
    .D(_01850_),
    .X(_01851_));
 sky130_fd_sc_hd__nor2_8 _05313_ (.A(_01846_),
    .B(_01851_),
    .Y(_01852_));
 sky130_fd_sc_hd__mux2_1 _05314_ (.A0(\tms1x00.ins_pla_ands[21][11] ),
    .A1(\tms1x00.ins_pla_ands[21][10] ),
    .S(net677),
    .X(_01853_));
 sky130_fd_sc_hd__mux2_1 _05315_ (.A0(\tms1x00.ins_pla_ands[21][7] ),
    .A1(\tms1x00.ins_pla_ands[21][6] ),
    .S(net687),
    .X(_01854_));
 sky130_fd_sc_hd__mux2_1 _05316_ (.A0(\tms1x00.ins_pla_ands[21][3] ),
    .A1(\tms1x00.ins_pla_ands[21][2] ),
    .S(net696),
    .X(_01855_));
 sky130_fd_sc_hd__mux2_1 _05317_ (.A0(\tms1x00.ins_pla_ands[21][5] ),
    .A1(\tms1x00.ins_pla_ands[21][4] ),
    .S(net691),
    .X(_01856_));
 sky130_fd_sc_hd__or4_4 _05318_ (.A(_01853_),
    .B(_01854_),
    .C(_01855_),
    .D(_01856_),
    .X(_01857_));
 sky130_fd_sc_hd__mux2_1 _05319_ (.A0(\tms1x00.ins_pla_ands[21][1] ),
    .A1(\tms1x00.ins_pla_ands[21][0] ),
    .S(net700),
    .X(_01858_));
 sky130_fd_sc_hd__mux2_1 _05320_ (.A0(\tms1x00.ins_pla_ands[21][13] ),
    .A1(\tms1x00.ins_pla_ands[21][12] ),
    .S(net673),
    .X(_01859_));
 sky130_fd_sc_hd__mux2_1 _05321_ (.A0(\tms1x00.ins_pla_ands[21][15] ),
    .A1(\tms1x00.ins_pla_ands[21][14] ),
    .S(net667),
    .X(_01860_));
 sky130_fd_sc_hd__mux2_1 _05322_ (.A0(\tms1x00.ins_pla_ands[21][9] ),
    .A1(\tms1x00.ins_pla_ands[21][8] ),
    .S(net683),
    .X(_01861_));
 sky130_fd_sc_hd__or4_4 _05323_ (.A(_01858_),
    .B(_01859_),
    .C(_01860_),
    .D(_01861_),
    .X(_01862_));
 sky130_fd_sc_hd__nor2_8 _05324_ (.A(_01857_),
    .B(_01862_),
    .Y(_01863_));
 sky130_fd_sc_hd__mux2_1 _05325_ (.A0(\tms1x00.ins_pla_ands[22][11] ),
    .A1(\tms1x00.ins_pla_ands[22][10] ),
    .S(net677),
    .X(_01864_));
 sky130_fd_sc_hd__mux2_1 _05326_ (.A0(\tms1x00.ins_pla_ands[22][7] ),
    .A1(\tms1x00.ins_pla_ands[22][6] ),
    .S(net690),
    .X(_01865_));
 sky130_fd_sc_hd__mux2_1 _05327_ (.A0(\tms1x00.ins_pla_ands[22][3] ),
    .A1(\tms1x00.ins_pla_ands[22][2] ),
    .S(net699),
    .X(_01866_));
 sky130_fd_sc_hd__mux2_1 _05328_ (.A0(\tms1x00.ins_pla_ands[22][5] ),
    .A1(\tms1x00.ins_pla_ands[22][4] ),
    .S(net695),
    .X(_01867_));
 sky130_fd_sc_hd__or4_4 _05329_ (.A(_01864_),
    .B(_01865_),
    .C(_01866_),
    .D(_01867_),
    .X(_01868_));
 sky130_fd_sc_hd__mux2_1 _05330_ (.A0(\tms1x00.ins_pla_ands[22][1] ),
    .A1(\tms1x00.ins_pla_ands[22][0] ),
    .S(net700),
    .X(_01869_));
 sky130_fd_sc_hd__mux2_1 _05331_ (.A0(\tms1x00.ins_pla_ands[22][13] ),
    .A1(\tms1x00.ins_pla_ands[22][12] ),
    .S(net673),
    .X(_01870_));
 sky130_fd_sc_hd__mux2_1 _05332_ (.A0(\tms1x00.ins_pla_ands[22][15] ),
    .A1(\tms1x00.ins_pla_ands[22][14] ),
    .S(net667),
    .X(_01871_));
 sky130_fd_sc_hd__mux2_1 _05333_ (.A0(\tms1x00.ins_pla_ands[22][9] ),
    .A1(\tms1x00.ins_pla_ands[22][8] ),
    .S(net683),
    .X(_01872_));
 sky130_fd_sc_hd__or4_4 _05334_ (.A(_01869_),
    .B(_01870_),
    .C(_01871_),
    .D(_01872_),
    .X(_01873_));
 sky130_fd_sc_hd__nor2_8 _05335_ (.A(_01868_),
    .B(_01873_),
    .Y(_01874_));
 sky130_fd_sc_hd__mux2_1 _05336_ (.A0(\tms1x00.ins_pla_ands[9][5] ),
    .A1(\tms1x00.ins_pla_ands[9][4] ),
    .S(net692),
    .X(_01875_));
 sky130_fd_sc_hd__mux2_1 _05337_ (.A0(\tms1x00.ins_pla_ands[9][13] ),
    .A1(\tms1x00.ins_pla_ands[9][12] ),
    .S(net676),
    .X(_01876_));
 sky130_fd_sc_hd__mux2_1 _05338_ (.A0(\tms1x00.ins_pla_ands[9][7] ),
    .A1(\tms1x00.ins_pla_ands[9][6] ),
    .S(net686),
    .X(_01877_));
 sky130_fd_sc_hd__mux2_1 _05339_ (.A0(\tms1x00.ins_pla_ands[9][1] ),
    .A1(\tms1x00.ins_pla_ands[9][0] ),
    .S(net701),
    .X(_01878_));
 sky130_fd_sc_hd__or4_4 _05340_ (.A(_01875_),
    .B(_01876_),
    .C(_01877_),
    .D(_01878_),
    .X(_01879_));
 sky130_fd_sc_hd__mux2_1 _05341_ (.A0(\tms1x00.ins_pla_ands[9][3] ),
    .A1(\tms1x00.ins_pla_ands[9][2] ),
    .S(net698),
    .X(_01880_));
 sky130_fd_sc_hd__mux2_1 _05342_ (.A0(\tms1x00.ins_pla_ands[9][11] ),
    .A1(\tms1x00.ins_pla_ands[9][10] ),
    .S(net679),
    .X(_01881_));
 sky130_fd_sc_hd__mux2_1 _05343_ (.A0(\tms1x00.ins_pla_ands[9][15] ),
    .A1(\tms1x00.ins_pla_ands[9][14] ),
    .S(net670),
    .X(_01882_));
 sky130_fd_sc_hd__mux2_1 _05344_ (.A0(\tms1x00.ins_pla_ands[9][9] ),
    .A1(\tms1x00.ins_pla_ands[9][8] ),
    .S(net682),
    .X(_01883_));
 sky130_fd_sc_hd__or4_4 _05345_ (.A(_01880_),
    .B(_01881_),
    .C(_01882_),
    .D(_01883_),
    .X(_01884_));
 sky130_fd_sc_hd__nor2_8 _05346_ (.A(_01879_),
    .B(_01884_),
    .Y(_01885_));
 sky130_fd_sc_hd__mux2_1 _05347_ (.A0(\tms1x00.ins_pla_ands[17][5] ),
    .A1(\tms1x00.ins_pla_ands[17][4] ),
    .S(net695),
    .X(_01886_));
 sky130_fd_sc_hd__mux2_1 _05348_ (.A0(\tms1x00.ins_pla_ands[17][7] ),
    .A1(\tms1x00.ins_pla_ands[17][6] ),
    .S(net687),
    .X(_01887_));
 sky130_fd_sc_hd__mux2_1 _05349_ (.A0(\tms1x00.ins_pla_ands[17][13] ),
    .A1(\tms1x00.ins_pla_ands[17][12] ),
    .S(net676),
    .X(_01888_));
 sky130_fd_sc_hd__mux2_2 _05350_ (.A0(\tms1x00.ins_pla_ands[17][15] ),
    .A1(\tms1x00.ins_pla_ands[17][14] ),
    .S(net668),
    .X(_01889_));
 sky130_fd_sc_hd__mux2_1 _05351_ (.A0(\tms1x00.ins_pla_ands[17][11] ),
    .A1(\tms1x00.ins_pla_ands[17][10] ),
    .S(net677),
    .X(_01890_));
 sky130_fd_sc_hd__mux2_2 _05352_ (.A0(\tms1x00.ins_pla_ands[17][9] ),
    .A1(\tms1x00.ins_pla_ands[17][8] ),
    .S(net681),
    .X(_01891_));
 sky130_fd_sc_hd__mux2_1 _05353_ (.A0(\tms1x00.ins_pla_ands[17][3] ),
    .A1(\tms1x00.ins_pla_ands[17][2] ),
    .S(net696),
    .X(_01892_));
 sky130_fd_sc_hd__or4_4 _05354_ (.A(_01886_),
    .B(_01887_),
    .C(_01891_),
    .D(_01892_),
    .X(_01893_));
 sky130_fd_sc_hd__mux2_1 _05355_ (.A0(\tms1x00.ins_pla_ands[17][1] ),
    .A1(\tms1x00.ins_pla_ands[17][0] ),
    .S(net700),
    .X(_01894_));
 sky130_fd_sc_hd__or4_4 _05356_ (.A(_01888_),
    .B(_01889_),
    .C(_01890_),
    .D(_01894_),
    .X(_01895_));
 sky130_fd_sc_hd__nor2_8 _05357_ (.A(_01893_),
    .B(_01895_),
    .Y(_01896_));
 sky130_fd_sc_hd__mux2_1 _05358_ (.A0(\tms1x00.ins_pla_ands[15][11] ),
    .A1(\tms1x00.ins_pla_ands[15][10] ),
    .S(net679),
    .X(_01897_));
 sky130_fd_sc_hd__mux2_1 _05359_ (.A0(\tms1x00.ins_pla_ands[15][7] ),
    .A1(\tms1x00.ins_pla_ands[15][6] ),
    .S(net686),
    .X(_01898_));
 sky130_fd_sc_hd__mux2_1 _05360_ (.A0(\tms1x00.ins_pla_ands[15][3] ),
    .A1(\tms1x00.ins_pla_ands[15][2] ),
    .S(net697),
    .X(_01899_));
 sky130_fd_sc_hd__mux2_1 _05361_ (.A0(\tms1x00.ins_pla_ands[15][5] ),
    .A1(\tms1x00.ins_pla_ands[15][4] ),
    .S(net692),
    .X(_01900_));
 sky130_fd_sc_hd__or4_4 _05362_ (.A(_01897_),
    .B(_01898_),
    .C(_01899_),
    .D(_01900_),
    .X(_01901_));
 sky130_fd_sc_hd__mux2_2 _05363_ (.A0(\tms1x00.ins_pla_ands[15][1] ),
    .A1(\tms1x00.ins_pla_ands[15][0] ),
    .S(net701),
    .X(_01902_));
 sky130_fd_sc_hd__mux2_1 _05364_ (.A0(\tms1x00.ins_pla_ands[15][13] ),
    .A1(\tms1x00.ins_pla_ands[15][12] ),
    .S(net672),
    .X(_01903_));
 sky130_fd_sc_hd__mux2_1 _05365_ (.A0(\tms1x00.ins_pla_ands[15][15] ),
    .A1(\tms1x00.ins_pla_ands[15][14] ),
    .S(net668),
    .X(_01904_));
 sky130_fd_sc_hd__mux2_1 _05366_ (.A0(\tms1x00.ins_pla_ands[15][9] ),
    .A1(\tms1x00.ins_pla_ands[15][8] ),
    .S(net682),
    .X(_01905_));
 sky130_fd_sc_hd__or4_4 _05367_ (.A(_01902_),
    .B(_01903_),
    .C(_01904_),
    .D(_01905_),
    .X(_01906_));
 sky130_fd_sc_hd__nor2_8 _05368_ (.A(_01901_),
    .B(_01906_),
    .Y(_01907_));
 sky130_fd_sc_hd__mux2_1 _05369_ (.A0(\tms1x00.ins_pla_ands[14][11] ),
    .A1(\tms1x00.ins_pla_ands[14][10] ),
    .S(net679),
    .X(_01908_));
 sky130_fd_sc_hd__mux2_1 _05370_ (.A0(\tms1x00.ins_pla_ands[14][7] ),
    .A1(\tms1x00.ins_pla_ands[14][6] ),
    .S(net686),
    .X(_01909_));
 sky130_fd_sc_hd__mux2_1 _05371_ (.A0(\tms1x00.ins_pla_ands[14][3] ),
    .A1(\tms1x00.ins_pla_ands[14][2] ),
    .S(net697),
    .X(_01910_));
 sky130_fd_sc_hd__mux2_1 _05372_ (.A0(\tms1x00.ins_pla_ands[14][5] ),
    .A1(\tms1x00.ins_pla_ands[14][4] ),
    .S(net692),
    .X(_01911_));
 sky130_fd_sc_hd__or4_4 _05373_ (.A(_01908_),
    .B(_01909_),
    .C(_01910_),
    .D(_01911_),
    .X(_01912_));
 sky130_fd_sc_hd__mux2_1 _05374_ (.A0(\tms1x00.ins_pla_ands[14][1] ),
    .A1(\tms1x00.ins_pla_ands[14][0] ),
    .S(net701),
    .X(_01913_));
 sky130_fd_sc_hd__mux2_2 _05375_ (.A0(\tms1x00.ins_pla_ands[14][13] ),
    .A1(\tms1x00.ins_pla_ands[14][12] ),
    .S(net672),
    .X(_01914_));
 sky130_fd_sc_hd__mux2_1 _05376_ (.A0(\tms1x00.ins_pla_ands[14][15] ),
    .A1(\tms1x00.ins_pla_ands[14][14] ),
    .S(net668),
    .X(_01915_));
 sky130_fd_sc_hd__mux2_2 _05377_ (.A0(\tms1x00.ins_pla_ands[14][9] ),
    .A1(\tms1x00.ins_pla_ands[14][8] ),
    .S(net681),
    .X(_01916_));
 sky130_fd_sc_hd__or4_4 _05378_ (.A(_01913_),
    .B(_01914_),
    .C(_01915_),
    .D(_01916_),
    .X(_01917_));
 sky130_fd_sc_hd__nor2_8 _05379_ (.A(_01912_),
    .B(_01917_),
    .Y(_01918_));
 sky130_fd_sc_hd__mux2_1 _05380_ (.A0(\tms1x00.ins_pla_ands[19][1] ),
    .A1(\tms1x00.ins_pla_ands[19][0] ),
    .S(net704),
    .X(_01919_));
 sky130_fd_sc_hd__mux2_1 _05381_ (.A0(\tms1x00.ins_pla_ands[19][7] ),
    .A1(\tms1x00.ins_pla_ands[19][6] ),
    .S(net689),
    .X(_01920_));
 sky130_fd_sc_hd__mux2_1 _05382_ (.A0(\tms1x00.ins_pla_ands[19][5] ),
    .A1(\tms1x00.ins_pla_ands[19][4] ),
    .S(net695),
    .X(_01921_));
 sky130_fd_sc_hd__mux2_2 _05383_ (.A0(\tms1x00.ins_pla_ands[19][9] ),
    .A1(\tms1x00.ins_pla_ands[19][8] ),
    .S(net682),
    .X(_01922_));
 sky130_fd_sc_hd__or4_4 _05384_ (.A(_01919_),
    .B(_01920_),
    .C(_01921_),
    .D(_01922_),
    .X(_01923_));
 sky130_fd_sc_hd__mux2_1 _05385_ (.A0(\tms1x00.ins_pla_ands[19][11] ),
    .A1(\tms1x00.ins_pla_ands[19][10] ),
    .S(net677),
    .X(_01924_));
 sky130_fd_sc_hd__mux2_1 _05386_ (.A0(\tms1x00.ins_pla_ands[19][13] ),
    .A1(\tms1x00.ins_pla_ands[19][12] ),
    .S(net673),
    .X(_01925_));
 sky130_fd_sc_hd__mux2_1 _05387_ (.A0(\tms1x00.ins_pla_ands[19][3] ),
    .A1(\tms1x00.ins_pla_ands[19][2] ),
    .S(net696),
    .X(_01926_));
 sky130_fd_sc_hd__mux2_1 _05388_ (.A0(\tms1x00.ins_pla_ands[19][15] ),
    .A1(\tms1x00.ins_pla_ands[19][14] ),
    .S(net667),
    .X(_01927_));
 sky130_fd_sc_hd__or4_4 _05389_ (.A(_01924_),
    .B(_01925_),
    .C(_01926_),
    .D(_01927_),
    .X(_01928_));
 sky130_fd_sc_hd__nor2_8 _05390_ (.A(_01923_),
    .B(_01928_),
    .Y(_01929_));
 sky130_fd_sc_hd__mux2_1 _05391_ (.A0(\tms1x00.ins_pla_ands[25][1] ),
    .A1(\tms1x00.ins_pla_ands[25][0] ),
    .S(net700),
    .X(_01930_));
 sky130_fd_sc_hd__mux2_1 _05392_ (.A0(\tms1x00.ins_pla_ands[25][7] ),
    .A1(\tms1x00.ins_pla_ands[25][6] ),
    .S(net687),
    .X(_01931_));
 sky130_fd_sc_hd__mux2_1 _05393_ (.A0(\tms1x00.ins_pla_ands[25][5] ),
    .A1(\tms1x00.ins_pla_ands[25][4] ),
    .S(net691),
    .X(_01932_));
 sky130_fd_sc_hd__mux2_1 _05394_ (.A0(\tms1x00.ins_pla_ands[25][9] ),
    .A1(\tms1x00.ins_pla_ands[25][8] ),
    .S(net683),
    .X(_01933_));
 sky130_fd_sc_hd__or4_4 _05395_ (.A(_01930_),
    .B(_01931_),
    .C(_01932_),
    .D(_01933_),
    .X(_01934_));
 sky130_fd_sc_hd__mux2_1 _05396_ (.A0(\tms1x00.ins_pla_ands[25][3] ),
    .A1(\tms1x00.ins_pla_ands[25][2] ),
    .S(net696),
    .X(_01935_));
 sky130_fd_sc_hd__mux2_1 _05397_ (.A0(\tms1x00.ins_pla_ands[25][13] ),
    .A1(\tms1x00.ins_pla_ands[25][12] ),
    .S(net673),
    .X(_01936_));
 sky130_fd_sc_hd__mux2_1 _05398_ (.A0(\tms1x00.ins_pla_ands[25][11] ),
    .A1(\tms1x00.ins_pla_ands[25][10] ),
    .S(net678),
    .X(_01937_));
 sky130_fd_sc_hd__mux2_1 _05399_ (.A0(\tms1x00.ins_pla_ands[25][15] ),
    .A1(\tms1x00.ins_pla_ands[25][14] ),
    .S(net667),
    .X(_01938_));
 sky130_fd_sc_hd__or4_4 _05400_ (.A(_01935_),
    .B(_01936_),
    .C(_01937_),
    .D(_01938_),
    .X(_01939_));
 sky130_fd_sc_hd__nor2_8 _05401_ (.A(_01934_),
    .B(_01939_),
    .Y(_01940_));
 sky130_fd_sc_hd__mux2_1 _05402_ (.A0(\tms1x00.ins_pla_ands[5][11] ),
    .A1(\tms1x00.ins_pla_ands[5][10] ),
    .S(net680),
    .X(_01941_));
 sky130_fd_sc_hd__mux2_1 _05403_ (.A0(\tms1x00.ins_pla_ands[5][7] ),
    .A1(\tms1x00.ins_pla_ands[5][6] ),
    .S(net688),
    .X(_01942_));
 sky130_fd_sc_hd__mux2_1 _05404_ (.A0(\tms1x00.ins_pla_ands[5][3] ),
    .A1(\tms1x00.ins_pla_ands[5][2] ),
    .S(net698),
    .X(_01943_));
 sky130_fd_sc_hd__mux2_1 _05405_ (.A0(\tms1x00.ins_pla_ands[5][5] ),
    .A1(\tms1x00.ins_pla_ands[5][4] ),
    .S(net694),
    .X(_01944_));
 sky130_fd_sc_hd__or4_2 _05406_ (.A(_01941_),
    .B(_01942_),
    .C(_01943_),
    .D(_01944_),
    .X(_01945_));
 sky130_fd_sc_hd__mux2_1 _05407_ (.A0(\tms1x00.ins_pla_ands[5][1] ),
    .A1(\tms1x00.ins_pla_ands[5][0] ),
    .S(net703),
    .X(_01946_));
 sky130_fd_sc_hd__mux2_1 _05408_ (.A0(\tms1x00.ins_pla_ands[5][13] ),
    .A1(\tms1x00.ins_pla_ands[5][12] ),
    .S(net674),
    .X(_01947_));
 sky130_fd_sc_hd__mux2_1 _05409_ (.A0(\tms1x00.ins_pla_ands[5][15] ),
    .A1(\tms1x00.ins_pla_ands[5][14] ),
    .S(net671),
    .X(_01948_));
 sky130_fd_sc_hd__mux2_1 _05410_ (.A0(\tms1x00.ins_pla_ands[5][9] ),
    .A1(\tms1x00.ins_pla_ands[5][8] ),
    .S(net684),
    .X(_01949_));
 sky130_fd_sc_hd__or4_2 _05411_ (.A(_01946_),
    .B(_01947_),
    .C(_01948_),
    .D(_01949_),
    .X(_01950_));
 sky130_fd_sc_hd__nor2_4 _05412_ (.A(_01945_),
    .B(_01950_),
    .Y(_01951_));
 sky130_fd_sc_hd__mux2_1 _05413_ (.A0(\tms1x00.ins_pla_ands[6][11] ),
    .A1(\tms1x00.ins_pla_ands[6][10] ),
    .S(net680),
    .X(_01952_));
 sky130_fd_sc_hd__mux2_1 _05414_ (.A0(\tms1x00.ins_pla_ands[6][7] ),
    .A1(\tms1x00.ins_pla_ands[6][6] ),
    .S(net689),
    .X(_01953_));
 sky130_fd_sc_hd__mux2_1 _05415_ (.A0(\tms1x00.ins_pla_ands[6][3] ),
    .A1(\tms1x00.ins_pla_ands[6][2] ),
    .S(net698),
    .X(_01954_));
 sky130_fd_sc_hd__mux2_1 _05416_ (.A0(\tms1x00.ins_pla_ands[6][5] ),
    .A1(\tms1x00.ins_pla_ands[6][4] ),
    .S(net694),
    .X(_01955_));
 sky130_fd_sc_hd__or4_4 _05417_ (.A(_01952_),
    .B(_01953_),
    .C(_01954_),
    .D(_01955_),
    .X(_01956_));
 sky130_fd_sc_hd__mux2_1 _05418_ (.A0(\tms1x00.ins_pla_ands[6][1] ),
    .A1(\tms1x00.ins_pla_ands[6][0] ),
    .S(net703),
    .X(_01957_));
 sky130_fd_sc_hd__mux2_1 _05419_ (.A0(\tms1x00.ins_pla_ands[6][13] ),
    .A1(\tms1x00.ins_pla_ands[6][12] ),
    .S(net674),
    .X(_01958_));
 sky130_fd_sc_hd__mux2_1 _05420_ (.A0(\tms1x00.ins_pla_ands[6][15] ),
    .A1(\tms1x00.ins_pla_ands[6][14] ),
    .S(net670),
    .X(_01959_));
 sky130_fd_sc_hd__mux2_1 _05421_ (.A0(\tms1x00.ins_pla_ands[6][9] ),
    .A1(\tms1x00.ins_pla_ands[6][8] ),
    .S(net684),
    .X(_01960_));
 sky130_fd_sc_hd__or4_4 _05422_ (.A(_01957_),
    .B(_01958_),
    .C(_01959_),
    .D(_01960_),
    .X(_01961_));
 sky130_fd_sc_hd__nor2_8 _05423_ (.A(_01956_),
    .B(_01961_),
    .Y(_01962_));
 sky130_fd_sc_hd__mux2_1 _05424_ (.A0(\tms1x00.ins_pla_ands[8][5] ),
    .A1(\tms1x00.ins_pla_ands[8][4] ),
    .S(\tms1x00.ins_arg[5] ),
    .X(_01963_));
 sky130_fd_sc_hd__mux2_1 _05425_ (.A0(\tms1x00.ins_pla_ands[8][13] ),
    .A1(\tms1x00.ins_pla_ands[8][12] ),
    .S(net672),
    .X(_01964_));
 sky130_fd_sc_hd__mux2_1 _05426_ (.A0(\tms1x00.ins_pla_ands[8][7] ),
    .A1(\tms1x00.ins_pla_ands[8][6] ),
    .S(net686),
    .X(_01965_));
 sky130_fd_sc_hd__mux2_1 _05427_ (.A0(\tms1x00.ins_pla_ands[8][1] ),
    .A1(\tms1x00.ins_pla_ands[8][0] ),
    .S(net701),
    .X(_01966_));
 sky130_fd_sc_hd__or4_4 _05428_ (.A(_01963_),
    .B(_01964_),
    .C(_01965_),
    .D(_01966_),
    .X(_01967_));
 sky130_fd_sc_hd__mux2_1 _05429_ (.A0(\tms1x00.ins_pla_ands[8][3] ),
    .A1(\tms1x00.ins_pla_ands[8][2] ),
    .S(net697),
    .X(_01968_));
 sky130_fd_sc_hd__mux2_1 _05430_ (.A0(\tms1x00.ins_pla_ands[8][11] ),
    .A1(\tms1x00.ins_pla_ands[8][10] ),
    .S(net679),
    .X(_01969_));
 sky130_fd_sc_hd__mux2_1 _05431_ (.A0(\tms1x00.ins_pla_ands[8][15] ),
    .A1(\tms1x00.ins_pla_ands[8][14] ),
    .S(net669),
    .X(_01970_));
 sky130_fd_sc_hd__mux2_1 _05432_ (.A0(\tms1x00.ins_pla_ands[8][9] ),
    .A1(\tms1x00.ins_pla_ands[8][8] ),
    .S(net682),
    .X(_01971_));
 sky130_fd_sc_hd__or4_4 _05433_ (.A(_01968_),
    .B(_01969_),
    .C(_01970_),
    .D(_01971_),
    .X(_01972_));
 sky130_fd_sc_hd__nor2_8 _05434_ (.A(_01967_),
    .B(_01972_),
    .Y(_01973_));
 sky130_fd_sc_hd__a22o_1 _05435_ (.A1(\tms1x00.ins_pla_ors[1][10] ),
    .A2(net420),
    .B1(net416),
    .B2(\tms1x00.ins_pla_ors[1][22] ),
    .X(_01974_));
 sky130_fd_sc_hd__a22o_1 _05436_ (.A1(\tms1x00.ins_pla_ors[1][15] ),
    .A2(net410),
    .B1(net403),
    .B2(\tms1x00.ins_pla_ors[1][5] ),
    .X(_01975_));
 sky130_fd_sc_hd__a22o_1 _05437_ (.A1(\tms1x00.ins_pla_ors[1][18] ),
    .A2(net431),
    .B1(net414),
    .B2(\tms1x00.ins_pla_ors[1][9] ),
    .X(_01976_));
 sky130_fd_sc_hd__a22o_1 _05438_ (.A1(\tms1x00.ins_pla_ors[1][11] ),
    .A2(net448),
    .B1(net442),
    .B2(\tms1x00.ins_pla_ors[1][4] ),
    .X(_01977_));
 sky130_fd_sc_hd__a22o_1 _05439_ (.A1(\tms1x00.ins_pla_ors[1][16] ),
    .A2(net444),
    .B1(net412),
    .B2(\tms1x00.ins_pla_ors[1][17] ),
    .X(_01978_));
 sky130_fd_sc_hd__a22o_1 _05440_ (.A1(\tms1x00.ins_pla_ors[1][25] ),
    .A2(net404),
    .B1(net398),
    .B2(\tms1x00.ins_pla_ors[1][8] ),
    .X(_01979_));
 sky130_fd_sc_hd__a221o_1 _05441_ (.A1(\tms1x00.ins_pla_ors[1][2] ),
    .A2(net438),
    .B1(net434),
    .B2(\tms1x00.ins_pla_ors[1][1] ),
    .C1(_01979_),
    .X(_01980_));
 sky130_fd_sc_hd__a22o_1 _05442_ (.A1(\tms1x00.ins_pla_ors[1][27] ),
    .A2(net422),
    .B1(net406),
    .B2(\tms1x00.ins_pla_ors[1][19] ),
    .X(_01981_));
 sky130_fd_sc_hd__a221o_1 _05443_ (.A1(\tms1x00.ins_pla_ors[1][29] ),
    .A2(net428),
    .B1(net424),
    .B2(\tms1x00.ins_pla_ors[1][12] ),
    .C1(_01981_),
    .X(_01982_));
 sky130_fd_sc_hd__a22o_1 _05444_ (.A1(\tms1x00.ins_pla_ors[1][24] ),
    .A2(net456),
    .B1(net440),
    .B2(\tms1x00.ins_pla_ors[1][0] ),
    .X(_01983_));
 sky130_fd_sc_hd__a221o_2 _05445_ (.A1(\tms1x00.ins_pla_ors[1][20] ),
    .A2(net452),
    .B1(net408),
    .B2(\tms1x00.ins_pla_ors[1][14] ),
    .C1(_01978_),
    .X(_01984_));
 sky130_fd_sc_hd__a221o_1 _05446_ (.A1(\tms1x00.ins_pla_ors[1][7] ),
    .A2(net450),
    .B1(net432),
    .B2(\tms1x00.ins_pla_ors[1][3] ),
    .C1(_01977_),
    .X(_01985_));
 sky130_fd_sc_hd__a221o_1 _05447_ (.A1(\tms1x00.ins_pla_ors[1][13] ),
    .A2(net436),
    .B1(net400),
    .B2(\tms1x00.ins_pla_ors[1][6] ),
    .C1(_01983_),
    .X(_01986_));
 sky130_fd_sc_hd__a221o_2 _05448_ (.A1(\tms1x00.ins_pla_ors[1][26] ),
    .A2(net454),
    .B1(net446),
    .B2(\tms1x00.ins_pla_ors[1][28] ),
    .C1(_01974_),
    .X(_01987_));
 sky130_fd_sc_hd__or4_1 _05449_ (.A(_01984_),
    .B(_01985_),
    .C(_01986_),
    .D(_01987_),
    .X(_01988_));
 sky130_fd_sc_hd__a221o_1 _05450_ (.A1(\tms1x00.ins_pla_ors[1][23] ),
    .A2(net426),
    .B1(net418),
    .B2(\tms1x00.ins_pla_ors[1][21] ),
    .C1(_01976_),
    .X(_01989_));
 sky130_fd_sc_hd__or4_1 _05451_ (.A(_01975_),
    .B(_01980_),
    .C(_01982_),
    .D(_01989_),
    .X(_01990_));
 sky130_fd_sc_hd__or2_4 _05452_ (.A(_01988_),
    .B(_01990_),
    .X(_01991_));
 sky130_fd_sc_hd__a22o_1 _05453_ (.A1(\tms1x00.ins_pla_ors[0][25] ),
    .A2(net405),
    .B1(net399),
    .B2(\tms1x00.ins_pla_ors[0][8] ),
    .X(_01992_));
 sky130_fd_sc_hd__a22o_1 _05454_ (.A1(\tms1x00.ins_pla_ors[0][27] ),
    .A2(net423),
    .B1(net406),
    .B2(\tms1x00.ins_pla_ors[0][19] ),
    .X(_01993_));
 sky130_fd_sc_hd__a221o_1 _05455_ (.A1(\tms1x00.ins_pla_ors[0][29] ),
    .A2(net428),
    .B1(net425),
    .B2(\tms1x00.ins_pla_ors[0][12] ),
    .C1(_01993_),
    .X(_01994_));
 sky130_fd_sc_hd__a221o_1 _05456_ (.A1(\tms1x00.ins_pla_ors[0][2] ),
    .A2(net439),
    .B1(net435),
    .B2(\tms1x00.ins_pla_ors[0][1] ),
    .C1(_01992_),
    .X(_01995_));
 sky130_fd_sc_hd__a22o_1 _05457_ (.A1(\tms1x00.ins_pla_ors[0][16] ),
    .A2(net445),
    .B1(net413),
    .B2(\tms1x00.ins_pla_ors[0][17] ),
    .X(_01996_));
 sky130_fd_sc_hd__a22o_1 _05458_ (.A1(\tms1x00.ins_pla_ors[0][11] ),
    .A2(net448),
    .B1(net443),
    .B2(\tms1x00.ins_pla_ors[0][4] ),
    .X(_01997_));
 sky130_fd_sc_hd__a22o_1 _05459_ (.A1(\tms1x00.ins_pla_ors[0][18] ),
    .A2(net431),
    .B1(net414),
    .B2(\tms1x00.ins_pla_ors[0][9] ),
    .X(_01998_));
 sky130_fd_sc_hd__a22o_1 _05460_ (.A1(\tms1x00.ins_pla_ors[0][10] ),
    .A2(net421),
    .B1(net416),
    .B2(\tms1x00.ins_pla_ors[0][22] ),
    .X(_01999_));
 sky130_fd_sc_hd__a22o_1 _05461_ (.A1(\tms1x00.ins_pla_ors[0][24] ),
    .A2(net457),
    .B1(net441),
    .B2(\tms1x00.ins_pla_ors[0][0] ),
    .X(_02000_));
 sky130_fd_sc_hd__a221o_2 _05462_ (.A1(\tms1x00.ins_pla_ors[0][20] ),
    .A2(net453),
    .B1(net408),
    .B2(\tms1x00.ins_pla_ors[0][14] ),
    .C1(_01996_),
    .X(_02001_));
 sky130_fd_sc_hd__a221o_1 _05463_ (.A1(\tms1x00.ins_pla_ors[0][7] ),
    .A2(net451),
    .B1(net433),
    .B2(\tms1x00.ins_pla_ors[0][3] ),
    .C1(_01997_),
    .X(_02002_));
 sky130_fd_sc_hd__a221o_1 _05464_ (.A1(\tms1x00.ins_pla_ors[0][13] ),
    .A2(net437),
    .B1(net401),
    .B2(\tms1x00.ins_pla_ors[0][6] ),
    .C1(_02000_),
    .X(_02003_));
 sky130_fd_sc_hd__a221o_2 _05465_ (.A1(\tms1x00.ins_pla_ors[0][26] ),
    .A2(net455),
    .B1(net446),
    .B2(\tms1x00.ins_pla_ors[0][28] ),
    .C1(_01999_),
    .X(_02004_));
 sky130_fd_sc_hd__or4_1 _05466_ (.A(_02001_),
    .B(_02002_),
    .C(_02003_),
    .D(_02004_),
    .X(_02005_));
 sky130_fd_sc_hd__a221o_1 _05467_ (.A1(\tms1x00.ins_pla_ors[0][23] ),
    .A2(net426),
    .B1(net419),
    .B2(\tms1x00.ins_pla_ors[0][21] ),
    .C1(_01998_),
    .X(_02006_));
 sky130_fd_sc_hd__a22o_1 _05468_ (.A1(\tms1x00.ins_pla_ors[0][15] ),
    .A2(net410),
    .B1(net403),
    .B2(\tms1x00.ins_pla_ors[0][5] ),
    .X(_02007_));
 sky130_fd_sc_hd__or4_1 _05469_ (.A(_01994_),
    .B(_01995_),
    .C(_02006_),
    .D(_02007_),
    .X(_02008_));
 sky130_fd_sc_hd__or2_4 _05470_ (.A(_02005_),
    .B(_02008_),
    .X(_02009_));
 sky130_fd_sc_hd__or3_1 _05471_ (.A(net670),
    .B(net675),
    .C(_01625_),
    .X(_02010_));
 sky130_fd_sc_hd__or2_2 _05472_ (.A(_01626_),
    .B(_02010_),
    .X(_02011_));
 sky130_fd_sc_hd__nor2_2 _05473_ (.A(net688),
    .B(_02011_),
    .Y(_02012_));
 sky130_fd_sc_hd__or3_4 _05474_ (.A(_01991_),
    .B(_02009_),
    .C(_02012_),
    .X(_02013_));
 sky130_fd_sc_hd__and4b_4 _05475_ (.A_N(\tms1x00.cycle[2] ),
    .B(\tms1x00.cycle[1] ),
    .C(_01622_),
    .D(_02013_),
    .X(net157));
 sky130_fd_sc_hd__nor2_8 _05476_ (.A(net77),
    .B(net78),
    .Y(_02014_));
 sky130_fd_sc_hd__mux2_1 _05477_ (.A0(\wbs_o_buff[0] ),
    .A1(net42),
    .S(_02014_),
    .X(net180));
 sky130_fd_sc_hd__mux2_1 _05478_ (.A0(\wbs_o_buff[1] ),
    .A1(net53),
    .S(_02014_),
    .X(net191));
 sky130_fd_sc_hd__mux2_1 _05479_ (.A0(\wbs_o_buff[2] ),
    .A1(net64),
    .S(_02014_),
    .X(net202));
 sky130_fd_sc_hd__mux2_1 _05480_ (.A0(\wbs_o_buff[3] ),
    .A1(net67),
    .S(_02014_),
    .X(net205));
 sky130_fd_sc_hd__mux2_1 _05481_ (.A0(\wbs_o_buff[4] ),
    .A1(net68),
    .S(_02014_),
    .X(net206));
 sky130_fd_sc_hd__mux2_1 _05482_ (.A0(\wbs_o_buff[5] ),
    .A1(net69),
    .S(_02014_),
    .X(net207));
 sky130_fd_sc_hd__mux2_1 _05483_ (.A0(\wbs_o_buff[6] ),
    .A1(net70),
    .S(_02014_),
    .X(net208));
 sky130_fd_sc_hd__mux2_1 _05484_ (.A0(\wbs_o_buff[7] ),
    .A1(net71),
    .S(_02014_),
    .X(net209));
 sky130_fd_sc_hd__mux2_1 _05485_ (.A0(\wbs_o_buff[8] ),
    .A1(net72),
    .S(_02014_),
    .X(net210));
 sky130_fd_sc_hd__mux2_1 _05486_ (.A0(\wbs_o_buff[9] ),
    .A1(net73),
    .S(_02014_),
    .X(net211));
 sky130_fd_sc_hd__mux2_1 _05487_ (.A0(\wbs_o_buff[10] ),
    .A1(net43),
    .S(_02014_),
    .X(net181));
 sky130_fd_sc_hd__mux2_1 _05488_ (.A0(\wbs_o_buff[11] ),
    .A1(net44),
    .S(_02014_),
    .X(net182));
 sky130_fd_sc_hd__mux2_1 _05489_ (.A0(\wbs_o_buff[12] ),
    .A1(net45),
    .S(_02014_),
    .X(net183));
 sky130_fd_sc_hd__mux2_1 _05490_ (.A0(\wbs_o_buff[13] ),
    .A1(net46),
    .S(_02014_),
    .X(net184));
 sky130_fd_sc_hd__mux2_2 _05491_ (.A0(\wbs_o_buff[14] ),
    .A1(net47),
    .S(_02014_),
    .X(net185));
 sky130_fd_sc_hd__mux2_2 _05492_ (.A0(\wbs_o_buff[15] ),
    .A1(net48),
    .S(_02014_),
    .X(net186));
 sky130_fd_sc_hd__mux2_1 _05493_ (.A0(\wbs_o_buff[16] ),
    .A1(net49),
    .S(_02014_),
    .X(net187));
 sky130_fd_sc_hd__mux2_1 _05494_ (.A0(\wbs_o_buff[17] ),
    .A1(net50),
    .S(_02014_),
    .X(net188));
 sky130_fd_sc_hd__mux2_1 _05495_ (.A0(\wbs_o_buff[18] ),
    .A1(net51),
    .S(_02014_),
    .X(net189));
 sky130_fd_sc_hd__mux2_1 _05496_ (.A0(\wbs_o_buff[19] ),
    .A1(net52),
    .S(_02014_),
    .X(net190));
 sky130_fd_sc_hd__mux2_1 _05497_ (.A0(\wbs_o_buff[20] ),
    .A1(net54),
    .S(_02014_),
    .X(net192));
 sky130_fd_sc_hd__mux2_1 _05498_ (.A0(\wbs_o_buff[21] ),
    .A1(net55),
    .S(_02014_),
    .X(net193));
 sky130_fd_sc_hd__mux2_1 _05499_ (.A0(\wbs_o_buff[22] ),
    .A1(net56),
    .S(_02014_),
    .X(net194));
 sky130_fd_sc_hd__mux2_1 _05500_ (.A0(\wbs_o_buff[23] ),
    .A1(net57),
    .S(_02014_),
    .X(net195));
 sky130_fd_sc_hd__mux2_2 _05501_ (.A0(\wbs_o_buff[24] ),
    .A1(net58),
    .S(_02014_),
    .X(net196));
 sky130_fd_sc_hd__mux2_1 _05502_ (.A0(\wbs_o_buff[25] ),
    .A1(net59),
    .S(_02014_),
    .X(net197));
 sky130_fd_sc_hd__mux2_2 _05503_ (.A0(\wbs_o_buff[26] ),
    .A1(net60),
    .S(_02014_),
    .X(net198));
 sky130_fd_sc_hd__mux2_2 _05504_ (.A0(\wbs_o_buff[27] ),
    .A1(net61),
    .S(_02014_),
    .X(net199));
 sky130_fd_sc_hd__mux2_2 _05505_ (.A0(\wbs_o_buff[28] ),
    .A1(net62),
    .S(_02014_),
    .X(net200));
 sky130_fd_sc_hd__mux2_2 _05506_ (.A0(\wbs_o_buff[29] ),
    .A1(net63),
    .S(_02014_),
    .X(net201));
 sky130_fd_sc_hd__mux2_4 _05507_ (.A0(\wbs_o_buff[30] ),
    .A1(net65),
    .S(_02014_),
    .X(net203));
 sky130_fd_sc_hd__mux2_2 _05508_ (.A0(\wbs_o_buff[31] ),
    .A1(net66),
    .S(_02014_),
    .X(net204));
 sky130_fd_sc_hd__mux2_1 _05509_ (.A0(net2),
    .A1(\K_override[0] ),
    .S(net145),
    .X(\tms1x00.K_in[0] ));
 sky130_fd_sc_hd__mux2_1 _05510_ (.A0(net3),
    .A1(\K_override[1] ),
    .S(net145),
    .X(\tms1x00.K_in[1] ));
 sky130_fd_sc_hd__mux2_1 _05511_ (.A0(net4),
    .A1(\K_override[2] ),
    .S(net145),
    .X(\tms1x00.K_in[2] ));
 sky130_fd_sc_hd__mux2_1 _05512_ (.A0(net5),
    .A1(\K_override[3] ),
    .S(net145),
    .X(\tms1x00.K_in[3] ));
 sky130_fd_sc_hd__a22o_1 _05513_ (.A1(net644),
    .A2(\tms1x00.O_pla_ands[19][7] ),
    .B1(\tms1x00.O_pla_ands[19][4] ),
    .B2(net662),
    .X(_02015_));
 sky130_fd_sc_hd__a22o_1 _05514_ (.A1(net657),
    .A2(\tms1x00.O_pla_ands[19][8] ),
    .B1(\tms1x00.O_pla_ands[19][2] ),
    .B2(net663),
    .X(_02016_));
 sky130_fd_sc_hd__a221o_4 _05515_ (.A1(net640),
    .A2(\tms1x00.O_pla_ands[19][3] ),
    .B1(\tms1x00.O_pla_ands[19][0] ),
    .B2(net665),
    .C1(_02015_),
    .X(_02017_));
 sky130_fd_sc_hd__a221o_1 _05516_ (.A1(net646),
    .A2(\tms1x00.O_pla_ands[19][9] ),
    .B1(\tms1x00.O_pla_ands[19][5] ),
    .B2(net642),
    .C1(_02016_),
    .X(_02018_));
 sky130_fd_sc_hd__a221o_4 _05517_ (.A1(net659),
    .A2(\tms1x00.O_pla_ands[19][6] ),
    .B1(\tms1x00.O_pla_ands[19][1] ),
    .B2(net638),
    .C1(_02018_),
    .X(_02019_));
 sky130_fd_sc_hd__nor2_8 _05518_ (.A(_02017_),
    .B(_02019_),
    .Y(_02020_));
 sky130_fd_sc_hd__a22o_1 _05519_ (.A1(net645),
    .A2(\tms1x00.O_pla_ands[10][7] ),
    .B1(\tms1x00.O_pla_ands[10][4] ),
    .B2(net661),
    .X(_02021_));
 sky130_fd_sc_hd__a22o_1 _05520_ (.A1(net658),
    .A2(\tms1x00.O_pla_ands[10][8] ),
    .B1(\tms1x00.O_pla_ands[10][2] ),
    .B2(net664),
    .X(_02022_));
 sky130_fd_sc_hd__a221o_4 _05521_ (.A1(net641),
    .A2(\tms1x00.O_pla_ands[10][3] ),
    .B1(\tms1x00.O_pla_ands[10][0] ),
    .B2(net666),
    .C1(_02021_),
    .X(_02023_));
 sky130_fd_sc_hd__a221o_1 _05522_ (.A1(net647),
    .A2(\tms1x00.O_pla_ands[10][9] ),
    .B1(\tms1x00.O_pla_ands[10][5] ),
    .B2(net643),
    .C1(_02022_),
    .X(_02024_));
 sky130_fd_sc_hd__a221o_4 _05523_ (.A1(net660),
    .A2(\tms1x00.O_pla_ands[10][6] ),
    .B1(\tms1x00.O_pla_ands[10][1] ),
    .B2(net639),
    .C1(_02024_),
    .X(_02025_));
 sky130_fd_sc_hd__nor2_8 _05524_ (.A(_02023_),
    .B(_02025_),
    .Y(_02026_));
 sky130_fd_sc_hd__a22o_1 _05525_ (.A1(\tms1x00.O_pla_ors[0][19] ),
    .A2(_02020_),
    .B1(_02026_),
    .B2(\tms1x00.O_pla_ors[0][10] ),
    .X(_02027_));
 sky130_fd_sc_hd__a22o_1 _05526_ (.A1(net645),
    .A2(\tms1x00.O_pla_ands[2][7] ),
    .B1(\tms1x00.O_pla_ands[2][4] ),
    .B2(net661),
    .X(_02028_));
 sky130_fd_sc_hd__a22o_1 _05527_ (.A1(\tms1x00.O_latch[4] ),
    .A2(\tms1x00.O_pla_ands[2][8] ),
    .B1(\tms1x00.O_pla_ands[2][2] ),
    .B2(\tms1x00.O_latch[1] ),
    .X(_02029_));
 sky130_fd_sc_hd__a221o_4 _05528_ (.A1(net641),
    .A2(\tms1x00.O_pla_ands[2][3] ),
    .B1(\tms1x00.O_pla_ands[2][0] ),
    .B2(net666),
    .C1(_02028_),
    .X(_02030_));
 sky130_fd_sc_hd__a221o_1 _05529_ (.A1(net646),
    .A2(\tms1x00.O_pla_ands[2][9] ),
    .B1(\tms1x00.O_pla_ands[2][5] ),
    .B2(net642),
    .C1(_02029_),
    .X(_02031_));
 sky130_fd_sc_hd__a221o_4 _05530_ (.A1(net659),
    .A2(\tms1x00.O_pla_ands[2][6] ),
    .B1(\tms1x00.O_pla_ands[2][1] ),
    .B2(net638),
    .C1(_02031_),
    .X(_02032_));
 sky130_fd_sc_hd__nor2_8 _05531_ (.A(_02030_),
    .B(_02032_),
    .Y(_02033_));
 sky130_fd_sc_hd__a22o_1 _05532_ (.A1(net644),
    .A2(\tms1x00.O_pla_ands[6][7] ),
    .B1(\tms1x00.O_pla_ands[6][4] ),
    .B2(net662),
    .X(_02034_));
 sky130_fd_sc_hd__a22o_1 _05533_ (.A1(net657),
    .A2(\tms1x00.O_pla_ands[6][8] ),
    .B1(\tms1x00.O_pla_ands[6][2] ),
    .B2(net663),
    .X(_02035_));
 sky130_fd_sc_hd__a221o_4 _05534_ (.A1(net640),
    .A2(\tms1x00.O_pla_ands[6][3] ),
    .B1(\tms1x00.O_pla_ands[6][0] ),
    .B2(net665),
    .C1(_02034_),
    .X(_02036_));
 sky130_fd_sc_hd__a221o_1 _05535_ (.A1(net646),
    .A2(\tms1x00.O_pla_ands[6][9] ),
    .B1(\tms1x00.O_pla_ands[6][5] ),
    .B2(net642),
    .C1(_02035_),
    .X(_02037_));
 sky130_fd_sc_hd__a221o_4 _05536_ (.A1(net659),
    .A2(\tms1x00.O_pla_ands[6][6] ),
    .B1(\tms1x00.O_pla_ands[6][1] ),
    .B2(net638),
    .C1(_02037_),
    .X(_02038_));
 sky130_fd_sc_hd__nor2_8 _05537_ (.A(_02036_),
    .B(_02038_),
    .Y(_02039_));
 sky130_fd_sc_hd__a22o_1 _05538_ (.A1(net644),
    .A2(\tms1x00.O_pla_ands[17][7] ),
    .B1(\tms1x00.O_pla_ands[17][4] ),
    .B2(net662),
    .X(_02040_));
 sky130_fd_sc_hd__a22o_1 _05539_ (.A1(net657),
    .A2(\tms1x00.O_pla_ands[17][8] ),
    .B1(\tms1x00.O_pla_ands[17][2] ),
    .B2(net663),
    .X(_02041_));
 sky130_fd_sc_hd__a221o_4 _05540_ (.A1(net640),
    .A2(\tms1x00.O_pla_ands[17][3] ),
    .B1(\tms1x00.O_pla_ands[17][0] ),
    .B2(net665),
    .C1(_02040_),
    .X(_02042_));
 sky130_fd_sc_hd__a221o_1 _05541_ (.A1(net646),
    .A2(\tms1x00.O_pla_ands[17][9] ),
    .B1(\tms1x00.O_pla_ands[17][5] ),
    .B2(net642),
    .C1(_02041_),
    .X(_02043_));
 sky130_fd_sc_hd__a221o_4 _05542_ (.A1(net659),
    .A2(\tms1x00.O_pla_ands[17][6] ),
    .B1(\tms1x00.O_pla_ands[17][1] ),
    .B2(net638),
    .C1(_02043_),
    .X(_02044_));
 sky130_fd_sc_hd__nor2_8 _05543_ (.A(_02042_),
    .B(_02044_),
    .Y(_02045_));
 sky130_fd_sc_hd__a22o_1 _05544_ (.A1(net645),
    .A2(\tms1x00.O_pla_ands[8][7] ),
    .B1(\tms1x00.O_pla_ands[8][4] ),
    .B2(net661),
    .X(_02046_));
 sky130_fd_sc_hd__a22o_1 _05545_ (.A1(net658),
    .A2(\tms1x00.O_pla_ands[8][8] ),
    .B1(\tms1x00.O_pla_ands[8][2] ),
    .B2(net664),
    .X(_02047_));
 sky130_fd_sc_hd__a221o_4 _05546_ (.A1(net641),
    .A2(\tms1x00.O_pla_ands[8][3] ),
    .B1(\tms1x00.O_pla_ands[8][0] ),
    .B2(net666),
    .C1(_02046_),
    .X(_02048_));
 sky130_fd_sc_hd__a221o_1 _05547_ (.A1(net647),
    .A2(\tms1x00.O_pla_ands[8][9] ),
    .B1(\tms1x00.O_pla_ands[8][5] ),
    .B2(net643),
    .C1(_02047_),
    .X(_02049_));
 sky130_fd_sc_hd__a221o_4 _05548_ (.A1(net660),
    .A2(\tms1x00.O_pla_ands[8][6] ),
    .B1(\tms1x00.O_pla_ands[8][1] ),
    .B2(net639),
    .C1(_02049_),
    .X(_02050_));
 sky130_fd_sc_hd__nor2_8 _05549_ (.A(_02048_),
    .B(_02050_),
    .Y(_02051_));
 sky130_fd_sc_hd__a22o_1 _05550_ (.A1(net645),
    .A2(\tms1x00.O_pla_ands[11][7] ),
    .B1(\tms1x00.O_pla_ands[11][4] ),
    .B2(net661),
    .X(_02052_));
 sky130_fd_sc_hd__a22o_1 _05551_ (.A1(net658),
    .A2(\tms1x00.O_pla_ands[11][8] ),
    .B1(\tms1x00.O_pla_ands[11][2] ),
    .B2(\tms1x00.O_latch[1] ),
    .X(_02053_));
 sky130_fd_sc_hd__a221o_4 _05552_ (.A1(net641),
    .A2(\tms1x00.O_pla_ands[11][3] ),
    .B1(\tms1x00.O_pla_ands[11][0] ),
    .B2(net666),
    .C1(_02052_),
    .X(_02054_));
 sky130_fd_sc_hd__a221o_1 _05553_ (.A1(net647),
    .A2(\tms1x00.O_pla_ands[11][9] ),
    .B1(\tms1x00.O_pla_ands[11][5] ),
    .B2(net643),
    .C1(_02053_),
    .X(_02055_));
 sky130_fd_sc_hd__a221o_4 _05554_ (.A1(net660),
    .A2(\tms1x00.O_pla_ands[11][6] ),
    .B1(\tms1x00.O_pla_ands[11][1] ),
    .B2(net639),
    .C1(_02055_),
    .X(_02056_));
 sky130_fd_sc_hd__nor2_8 _05555_ (.A(_02054_),
    .B(_02056_),
    .Y(_02057_));
 sky130_fd_sc_hd__a22o_1 _05556_ (.A1(net645),
    .A2(\tms1x00.O_pla_ands[15][7] ),
    .B1(\tms1x00.O_pla_ands[15][4] ),
    .B2(net661),
    .X(_02058_));
 sky130_fd_sc_hd__a22o_1 _05557_ (.A1(net658),
    .A2(\tms1x00.O_pla_ands[15][8] ),
    .B1(\tms1x00.O_pla_ands[15][2] ),
    .B2(net664),
    .X(_02059_));
 sky130_fd_sc_hd__a221o_4 _05558_ (.A1(net641),
    .A2(\tms1x00.O_pla_ands[15][3] ),
    .B1(\tms1x00.O_pla_ands[15][0] ),
    .B2(net666),
    .C1(_02058_),
    .X(_02060_));
 sky130_fd_sc_hd__a221o_1 _05559_ (.A1(net647),
    .A2(\tms1x00.O_pla_ands[15][9] ),
    .B1(\tms1x00.O_pla_ands[15][5] ),
    .B2(net643),
    .C1(_02059_),
    .X(_02061_));
 sky130_fd_sc_hd__a221o_4 _05560_ (.A1(net660),
    .A2(\tms1x00.O_pla_ands[15][6] ),
    .B1(\tms1x00.O_pla_ands[15][1] ),
    .B2(net639),
    .C1(_02061_),
    .X(_02062_));
 sky130_fd_sc_hd__nor2_8 _05561_ (.A(_02060_),
    .B(_02062_),
    .Y(_02063_));
 sky130_fd_sc_hd__a22o_1 _05562_ (.A1(\tms1x00.O_pla_ands[3][7] ),
    .A2(net645),
    .B1(net661),
    .B2(\tms1x00.O_pla_ands[3][4] ),
    .X(_02064_));
 sky130_fd_sc_hd__a22o_1 _05563_ (.A1(\tms1x00.O_pla_ands[3][8] ),
    .A2(net658),
    .B1(net664),
    .B2(\tms1x00.O_pla_ands[3][2] ),
    .X(_02065_));
 sky130_fd_sc_hd__a221o_4 _05564_ (.A1(\tms1x00.O_pla_ands[3][3] ),
    .A2(net641),
    .B1(net639),
    .B2(\tms1x00.O_pla_ands[3][1] ),
    .C1(_02064_),
    .X(_02066_));
 sky130_fd_sc_hd__a221o_1 _05565_ (.A1(\tms1x00.O_pla_ands[3][9] ),
    .A2(net647),
    .B1(net643),
    .B2(\tms1x00.O_pla_ands[3][5] ),
    .C1(_02065_),
    .X(_02067_));
 sky130_fd_sc_hd__a221o_4 _05566_ (.A1(\tms1x00.O_pla_ands[3][6] ),
    .A2(net660),
    .B1(net665),
    .B2(\tms1x00.O_pla_ands[3][0] ),
    .C1(_02067_),
    .X(_02068_));
 sky130_fd_sc_hd__nor2_8 _05567_ (.A(_02066_),
    .B(_02068_),
    .Y(_02069_));
 sky130_fd_sc_hd__a22o_1 _05568_ (.A1(net658),
    .A2(\tms1x00.O_pla_ands[9][8] ),
    .B1(\tms1x00.O_pla_ands[9][2] ),
    .B2(net664),
    .X(_02070_));
 sky130_fd_sc_hd__a22o_1 _05569_ (.A1(net641),
    .A2(\tms1x00.O_pla_ands[9][3] ),
    .B1(\tms1x00.O_pla_ands[9][0] ),
    .B2(net666),
    .X(_02071_));
 sky130_fd_sc_hd__a221o_4 _05570_ (.A1(net645),
    .A2(\tms1x00.O_pla_ands[9][7] ),
    .B1(\tms1x00.O_pla_ands[9][4] ),
    .B2(net661),
    .C1(_02071_),
    .X(_02072_));
 sky130_fd_sc_hd__a221o_1 _05571_ (.A1(net647),
    .A2(\tms1x00.O_pla_ands[9][9] ),
    .B1(\tms1x00.O_pla_ands[9][5] ),
    .B2(net643),
    .C1(_02070_),
    .X(_02073_));
 sky130_fd_sc_hd__a221o_4 _05572_ (.A1(net660),
    .A2(\tms1x00.O_pla_ands[9][6] ),
    .B1(\tms1x00.O_pla_ands[9][1] ),
    .B2(net639),
    .C1(_02073_),
    .X(_02074_));
 sky130_fd_sc_hd__nor2_8 _05573_ (.A(_02072_),
    .B(_02074_),
    .Y(_02075_));
 sky130_fd_sc_hd__a22o_1 _05574_ (.A1(net644),
    .A2(\tms1x00.O_pla_ands[16][7] ),
    .B1(\tms1x00.O_pla_ands[16][4] ),
    .B2(net662),
    .X(_02076_));
 sky130_fd_sc_hd__a22o_1 _05575_ (.A1(net657),
    .A2(\tms1x00.O_pla_ands[16][8] ),
    .B1(\tms1x00.O_pla_ands[16][2] ),
    .B2(net663),
    .X(_02077_));
 sky130_fd_sc_hd__a221o_4 _05576_ (.A1(net640),
    .A2(\tms1x00.O_pla_ands[16][3] ),
    .B1(\tms1x00.O_pla_ands[16][0] ),
    .B2(net665),
    .C1(_02076_),
    .X(_02078_));
 sky130_fd_sc_hd__a221o_1 _05577_ (.A1(net646),
    .A2(\tms1x00.O_pla_ands[16][9] ),
    .B1(\tms1x00.O_pla_ands[16][5] ),
    .B2(net642),
    .C1(_02077_),
    .X(_02079_));
 sky130_fd_sc_hd__a221o_4 _05578_ (.A1(net659),
    .A2(\tms1x00.O_pla_ands[16][6] ),
    .B1(\tms1x00.O_pla_ands[16][1] ),
    .B2(net638),
    .C1(_02079_),
    .X(_02080_));
 sky130_fd_sc_hd__nor2_8 _05579_ (.A(_02078_),
    .B(_02080_),
    .Y(_02081_));
 sky130_fd_sc_hd__a22o_1 _05580_ (.A1(net645),
    .A2(\tms1x00.O_pla_ands[14][7] ),
    .B1(\tms1x00.O_pla_ands[14][4] ),
    .B2(net661),
    .X(_02082_));
 sky130_fd_sc_hd__a22o_1 _05581_ (.A1(net658),
    .A2(\tms1x00.O_pla_ands[14][8] ),
    .B1(\tms1x00.O_pla_ands[14][2] ),
    .B2(net664),
    .X(_02083_));
 sky130_fd_sc_hd__a221o_4 _05582_ (.A1(net641),
    .A2(\tms1x00.O_pla_ands[14][3] ),
    .B1(\tms1x00.O_pla_ands[14][0] ),
    .B2(net666),
    .C1(_02082_),
    .X(_02084_));
 sky130_fd_sc_hd__a221o_1 _05583_ (.A1(net647),
    .A2(\tms1x00.O_pla_ands[14][9] ),
    .B1(\tms1x00.O_pla_ands[14][5] ),
    .B2(net643),
    .C1(_02083_),
    .X(_02085_));
 sky130_fd_sc_hd__a221o_4 _05584_ (.A1(net660),
    .A2(\tms1x00.O_pla_ands[14][6] ),
    .B1(\tms1x00.O_pla_ands[14][1] ),
    .B2(net639),
    .C1(_02085_),
    .X(_02086_));
 sky130_fd_sc_hd__nor2_8 _05585_ (.A(_02084_),
    .B(_02086_),
    .Y(_02087_));
 sky130_fd_sc_hd__a22o_1 _05586_ (.A1(net644),
    .A2(\tms1x00.O_pla_ands[18][7] ),
    .B1(\tms1x00.O_pla_ands[18][4] ),
    .B2(net662),
    .X(_02088_));
 sky130_fd_sc_hd__a22o_1 _05587_ (.A1(net657),
    .A2(\tms1x00.O_pla_ands[18][8] ),
    .B1(\tms1x00.O_pla_ands[18][2] ),
    .B2(net663),
    .X(_02089_));
 sky130_fd_sc_hd__a221o_4 _05588_ (.A1(net640),
    .A2(\tms1x00.O_pla_ands[18][3] ),
    .B1(\tms1x00.O_pla_ands[18][0] ),
    .B2(net665),
    .C1(_02088_),
    .X(_02090_));
 sky130_fd_sc_hd__a221o_1 _05589_ (.A1(net646),
    .A2(\tms1x00.O_pla_ands[18][9] ),
    .B1(\tms1x00.O_pla_ands[18][5] ),
    .B2(net642),
    .C1(_02089_),
    .X(_02091_));
 sky130_fd_sc_hd__a221o_4 _05590_ (.A1(net659),
    .A2(\tms1x00.O_pla_ands[18][6] ),
    .B1(\tms1x00.O_pla_ands[18][1] ),
    .B2(net638),
    .C1(_02091_),
    .X(_02092_));
 sky130_fd_sc_hd__nor2_8 _05591_ (.A(_02090_),
    .B(_02092_),
    .Y(_02093_));
 sky130_fd_sc_hd__a22o_1 _05592_ (.A1(net644),
    .A2(\tms1x00.O_pla_ands[7][7] ),
    .B1(\tms1x00.O_pla_ands[7][4] ),
    .B2(net662),
    .X(_02094_));
 sky130_fd_sc_hd__a22o_1 _05593_ (.A1(net657),
    .A2(\tms1x00.O_pla_ands[7][8] ),
    .B1(\tms1x00.O_pla_ands[7][2] ),
    .B2(net663),
    .X(_02095_));
 sky130_fd_sc_hd__a221o_4 _05594_ (.A1(net640),
    .A2(\tms1x00.O_pla_ands[7][3] ),
    .B1(\tms1x00.O_pla_ands[7][0] ),
    .B2(net665),
    .C1(_02094_),
    .X(_02096_));
 sky130_fd_sc_hd__a221o_1 _05595_ (.A1(net647),
    .A2(\tms1x00.O_pla_ands[7][9] ),
    .B1(\tms1x00.O_pla_ands[7][5] ),
    .B2(net643),
    .C1(_02095_),
    .X(_02097_));
 sky130_fd_sc_hd__a221o_4 _05596_ (.A1(net659),
    .A2(\tms1x00.O_pla_ands[7][6] ),
    .B1(\tms1x00.O_pla_ands[7][1] ),
    .B2(net638),
    .C1(_02097_),
    .X(_02098_));
 sky130_fd_sc_hd__nor2_8 _05597_ (.A(_02096_),
    .B(_02098_),
    .Y(_02099_));
 sky130_fd_sc_hd__a22o_1 _05598_ (.A1(\tms1x00.O_pla_ands[4][7] ),
    .A2(net644),
    .B1(net662),
    .B2(\tms1x00.O_pla_ands[4][4] ),
    .X(_02100_));
 sky130_fd_sc_hd__a22o_1 _05599_ (.A1(\tms1x00.O_pla_ands[4][8] ),
    .A2(net657),
    .B1(net663),
    .B2(\tms1x00.O_pla_ands[4][2] ),
    .X(_02101_));
 sky130_fd_sc_hd__a221o_4 _05600_ (.A1(\tms1x00.O_pla_ands[4][3] ),
    .A2(net640),
    .B1(net639),
    .B2(\tms1x00.O_pla_ands[4][1] ),
    .C1(_02100_),
    .X(_02102_));
 sky130_fd_sc_hd__a221o_1 _05601_ (.A1(\tms1x00.O_pla_ands[4][9] ),
    .A2(net646),
    .B1(net642),
    .B2(\tms1x00.O_pla_ands[4][5] ),
    .C1(_02101_),
    .X(_02103_));
 sky130_fd_sc_hd__a221o_4 _05602_ (.A1(\tms1x00.O_pla_ands[4][6] ),
    .A2(net659),
    .B1(net666),
    .B2(\tms1x00.O_pla_ands[4][0] ),
    .C1(_02103_),
    .X(_02104_));
 sky130_fd_sc_hd__nor2_8 _05603_ (.A(_02102_),
    .B(_02104_),
    .Y(_02105_));
 sky130_fd_sc_hd__a22o_1 _05604_ (.A1(net644),
    .A2(\tms1x00.O_pla_ands[5][7] ),
    .B1(\tms1x00.O_pla_ands[5][4] ),
    .B2(net662),
    .X(_02106_));
 sky130_fd_sc_hd__a22o_1 _05605_ (.A1(net657),
    .A2(\tms1x00.O_pla_ands[5][8] ),
    .B1(\tms1x00.O_pla_ands[5][2] ),
    .B2(net663),
    .X(_02107_));
 sky130_fd_sc_hd__a221o_4 _05606_ (.A1(net640),
    .A2(\tms1x00.O_pla_ands[5][3] ),
    .B1(\tms1x00.O_pla_ands[5][0] ),
    .B2(net666),
    .C1(_02106_),
    .X(_02108_));
 sky130_fd_sc_hd__a221o_1 _05607_ (.A1(net646),
    .A2(\tms1x00.O_pla_ands[5][9] ),
    .B1(\tms1x00.O_pla_ands[5][5] ),
    .B2(net642),
    .C1(_02107_),
    .X(_02109_));
 sky130_fd_sc_hd__a221o_4 _05608_ (.A1(net659),
    .A2(\tms1x00.O_pla_ands[5][6] ),
    .B1(\tms1x00.O_pla_ands[5][1] ),
    .B2(net638),
    .C1(_02109_),
    .X(_02110_));
 sky130_fd_sc_hd__nor2_8 _05609_ (.A(_02108_),
    .B(_02110_),
    .Y(_02111_));
 sky130_fd_sc_hd__a22o_1 _05610_ (.A1(net658),
    .A2(\tms1x00.O_pla_ands[13][8] ),
    .B1(\tms1x00.O_pla_ands[13][2] ),
    .B2(net664),
    .X(_02112_));
 sky130_fd_sc_hd__a22o_1 _05611_ (.A1(net641),
    .A2(\tms1x00.O_pla_ands[13][3] ),
    .B1(\tms1x00.O_pla_ands[13][0] ),
    .B2(\tms1x00.O_latch[0] ),
    .X(_02113_));
 sky130_fd_sc_hd__a221o_4 _05612_ (.A1(net645),
    .A2(\tms1x00.O_pla_ands[13][7] ),
    .B1(\tms1x00.O_pla_ands[13][4] ),
    .B2(\tms1x00.O_latch[2] ),
    .C1(_02113_),
    .X(_02114_));
 sky130_fd_sc_hd__a221o_1 _05613_ (.A1(_01617_),
    .A2(\tms1x00.O_pla_ands[13][9] ),
    .B1(\tms1x00.O_pla_ands[13][5] ),
    .B2(_01619_),
    .C1(_02112_),
    .X(_02115_));
 sky130_fd_sc_hd__a221o_4 _05614_ (.A1(\tms1x00.O_latch[3] ),
    .A2(\tms1x00.O_pla_ands[13][6] ),
    .B1(\tms1x00.O_pla_ands[13][1] ),
    .B2(net639),
    .C1(_02115_),
    .X(_02116_));
 sky130_fd_sc_hd__nor2_8 _05615_ (.A(_02114_),
    .B(_02116_),
    .Y(_02117_));
 sky130_fd_sc_hd__a22o_1 _05616_ (.A1(net645),
    .A2(\tms1x00.O_pla_ands[12][7] ),
    .B1(\tms1x00.O_pla_ands[12][4] ),
    .B2(\tms1x00.O_latch[2] ),
    .X(_02118_));
 sky130_fd_sc_hd__a22o_1 _05617_ (.A1(net658),
    .A2(\tms1x00.O_pla_ands[12][8] ),
    .B1(\tms1x00.O_pla_ands[12][2] ),
    .B2(net664),
    .X(_02119_));
 sky130_fd_sc_hd__a221o_4 _05618_ (.A1(net641),
    .A2(\tms1x00.O_pla_ands[12][3] ),
    .B1(\tms1x00.O_pla_ands[12][0] ),
    .B2(\tms1x00.O_latch[0] ),
    .C1(_02118_),
    .X(_02120_));
 sky130_fd_sc_hd__a221o_1 _05619_ (.A1(net647),
    .A2(\tms1x00.O_pla_ands[12][9] ),
    .B1(\tms1x00.O_pla_ands[12][5] ),
    .B2(net643),
    .C1(_02119_),
    .X(_02121_));
 sky130_fd_sc_hd__a221o_4 _05620_ (.A1(net660),
    .A2(\tms1x00.O_pla_ands[12][6] ),
    .B1(\tms1x00.O_pla_ands[12][1] ),
    .B2(net639),
    .C1(_02121_),
    .X(_02122_));
 sky130_fd_sc_hd__nor2_8 _05621_ (.A(_02120_),
    .B(_02122_),
    .Y(_02123_));
 sky130_fd_sc_hd__a22o_1 _05622_ (.A1(\tms1x00.O_pla_ands[0][7] ),
    .A2(net644),
    .B1(net662),
    .B2(\tms1x00.O_pla_ands[0][4] ),
    .X(_02124_));
 sky130_fd_sc_hd__a22o_1 _05623_ (.A1(\tms1x00.O_pla_ands[0][8] ),
    .A2(net657),
    .B1(net663),
    .B2(\tms1x00.O_pla_ands[0][2] ),
    .X(_02125_));
 sky130_fd_sc_hd__a221o_4 _05624_ (.A1(\tms1x00.O_pla_ands[0][3] ),
    .A2(net640),
    .B1(net638),
    .B2(\tms1x00.O_pla_ands[0][1] ),
    .C1(_02124_),
    .X(_02126_));
 sky130_fd_sc_hd__a221o_1 _05625_ (.A1(\tms1x00.O_pla_ands[0][9] ),
    .A2(net646),
    .B1(net642),
    .B2(\tms1x00.O_pla_ands[0][5] ),
    .C1(_02125_),
    .X(_02127_));
 sky130_fd_sc_hd__a221o_4 _05626_ (.A1(\tms1x00.O_pla_ands[0][6] ),
    .A2(net659),
    .B1(net665),
    .B2(\tms1x00.O_pla_ands[0][0] ),
    .C1(_02127_),
    .X(_02128_));
 sky130_fd_sc_hd__nor2_8 _05627_ (.A(_02126_),
    .B(_02128_),
    .Y(_02129_));
 sky130_fd_sc_hd__a22o_1 _05628_ (.A1(\tms1x00.O_pla_ands[1][7] ),
    .A2(net644),
    .B1(net662),
    .B2(\tms1x00.O_pla_ands[1][4] ),
    .X(_02130_));
 sky130_fd_sc_hd__a22o_1 _05629_ (.A1(\tms1x00.O_pla_ands[1][8] ),
    .A2(net657),
    .B1(net663),
    .B2(\tms1x00.O_pla_ands[1][2] ),
    .X(_02131_));
 sky130_fd_sc_hd__a221o_4 _05630_ (.A1(\tms1x00.O_pla_ands[1][3] ),
    .A2(net640),
    .B1(net638),
    .B2(\tms1x00.O_pla_ands[1][1] ),
    .C1(_02130_),
    .X(_02132_));
 sky130_fd_sc_hd__a221o_1 _05631_ (.A1(\tms1x00.O_pla_ands[1][9] ),
    .A2(net646),
    .B1(net642),
    .B2(\tms1x00.O_pla_ands[1][5] ),
    .C1(_02131_),
    .X(_02133_));
 sky130_fd_sc_hd__a221o_4 _05632_ (.A1(\tms1x00.O_pla_ands[1][6] ),
    .A2(\tms1x00.O_latch[3] ),
    .B1(net665),
    .B2(\tms1x00.O_pla_ands[1][0] ),
    .C1(_02133_),
    .X(_02134_));
 sky130_fd_sc_hd__nor2_8 _05633_ (.A(_02132_),
    .B(_02134_),
    .Y(_02135_));
 sky130_fd_sc_hd__a22o_1 _05634_ (.A1(\tms1x00.O_pla_ors[0][5] ),
    .A2(_02111_),
    .B1(_02129_),
    .B2(\tms1x00.O_pla_ors[0][0] ),
    .X(_02136_));
 sky130_fd_sc_hd__a221o_1 _05635_ (.A1(\tms1x00.O_pla_ors[0][18] ),
    .A2(_02093_),
    .B1(_02135_),
    .B2(\tms1x00.O_pla_ors[0][1] ),
    .C1(_02136_),
    .X(_02137_));
 sky130_fd_sc_hd__a221o_1 _05636_ (.A1(\tms1x00.O_pla_ors[0][6] ),
    .A2(_02039_),
    .B1(_02075_),
    .B2(\tms1x00.O_pla_ors[0][9] ),
    .C1(_02027_),
    .X(_02138_));
 sky130_fd_sc_hd__a22o_1 _05637_ (.A1(\tms1x00.O_pla_ors[0][17] ),
    .A2(_02045_),
    .B1(_02105_),
    .B2(\tms1x00.O_pla_ors[0][4] ),
    .X(_02139_));
 sky130_fd_sc_hd__a221o_1 _05638_ (.A1(\tms1x00.O_pla_ors[0][13] ),
    .A2(_02117_),
    .B1(_02123_),
    .B2(\tms1x00.O_pla_ors[0][12] ),
    .C1(_02139_),
    .X(_02140_));
 sky130_fd_sc_hd__a22o_1 _05639_ (.A1(\tms1x00.O_pla_ors[0][2] ),
    .A2(_02033_),
    .B1(_02069_),
    .B2(\tms1x00.O_pla_ors[0][3] ),
    .X(_02141_));
 sky130_fd_sc_hd__a221o_1 _05640_ (.A1(\tms1x00.O_pla_ors[0][8] ),
    .A2(_02051_),
    .B1(_02057_),
    .B2(\tms1x00.O_pla_ors[0][11] ),
    .C1(_02141_),
    .X(_02142_));
 sky130_fd_sc_hd__a22o_1 _05641_ (.A1(\tms1x00.O_pla_ors[0][16] ),
    .A2(_02081_),
    .B1(_02099_),
    .B2(\tms1x00.O_pla_ors[0][7] ),
    .X(_02143_));
 sky130_fd_sc_hd__a221o_1 _05642_ (.A1(\tms1x00.O_pla_ors[0][15] ),
    .A2(_02063_),
    .B1(_02087_),
    .B2(\tms1x00.O_pla_ors[0][14] ),
    .C1(_02143_),
    .X(_02144_));
 sky130_fd_sc_hd__or3_1 _05643_ (.A(_02140_),
    .B(_02142_),
    .C(_02144_),
    .X(_02145_));
 sky130_fd_sc_hd__or3_4 _05644_ (.A(_02137_),
    .B(_02138_),
    .C(_02145_),
    .X(net120));
 sky130_fd_sc_hd__a22o_1 _05645_ (.A1(\tms1x00.O_pla_ors[1][15] ),
    .A2(_02063_),
    .B1(_02087_),
    .B2(\tms1x00.O_pla_ors[1][14] ),
    .X(_02146_));
 sky130_fd_sc_hd__a22o_1 _05646_ (.A1(\tms1x00.O_pla_ors[1][5] ),
    .A2(_02111_),
    .B1(_02129_),
    .B2(\tms1x00.O_pla_ors[1][0] ),
    .X(_02147_));
 sky130_fd_sc_hd__a22o_1 _05647_ (.A1(\tms1x00.O_pla_ors[1][18] ),
    .A2(_02093_),
    .B1(_02135_),
    .B2(\tms1x00.O_pla_ors[1][1] ),
    .X(_02148_));
 sky130_fd_sc_hd__a22o_1 _05648_ (.A1(\tms1x00.O_pla_ors[1][19] ),
    .A2(_02020_),
    .B1(_02026_),
    .B2(\tms1x00.O_pla_ors[1][10] ),
    .X(_02149_));
 sky130_fd_sc_hd__a221o_1 _05649_ (.A1(\tms1x00.O_pla_ors[1][6] ),
    .A2(_02039_),
    .B1(_02075_),
    .B2(\tms1x00.O_pla_ors[1][9] ),
    .C1(_02149_),
    .X(_02150_));
 sky130_fd_sc_hd__a22o_1 _05650_ (.A1(\tms1x00.O_pla_ors[1][17] ),
    .A2(_02045_),
    .B1(_02117_),
    .B2(\tms1x00.O_pla_ors[1][13] ),
    .X(_02151_));
 sky130_fd_sc_hd__a22o_1 _05651_ (.A1(\tms1x00.O_pla_ors[1][3] ),
    .A2(_02069_),
    .B1(_02123_),
    .B2(\tms1x00.O_pla_ors[1][12] ),
    .X(_02152_));
 sky130_fd_sc_hd__a221o_1 _05652_ (.A1(\tms1x00.O_pla_ors[1][2] ),
    .A2(_02033_),
    .B1(_02057_),
    .B2(\tms1x00.O_pla_ors[1][11] ),
    .C1(_02152_),
    .X(_02153_));
 sky130_fd_sc_hd__a211o_1 _05653_ (.A1(\tms1x00.O_pla_ors[1][8] ),
    .A2(_02051_),
    .B1(_02151_),
    .C1(_02153_),
    .X(_02154_));
 sky130_fd_sc_hd__a221o_1 _05654_ (.A1(\tms1x00.O_pla_ors[1][16] ),
    .A2(_02081_),
    .B1(_02099_),
    .B2(\tms1x00.O_pla_ors[1][7] ),
    .C1(_02146_),
    .X(_02155_));
 sky130_fd_sc_hd__or4_2 _05655_ (.A(_02147_),
    .B(_02148_),
    .C(_02150_),
    .D(_02155_),
    .X(_02156_));
 sky130_fd_sc_hd__a211o_4 _05656_ (.A1(\tms1x00.O_pla_ors[1][4] ),
    .A2(_02105_),
    .B1(_02154_),
    .C1(_02156_),
    .X(net121));
 sky130_fd_sc_hd__a22o_1 _05657_ (.A1(\tms1x00.O_pla_ors[2][17] ),
    .A2(_02045_),
    .B1(_02117_),
    .B2(\tms1x00.O_pla_ors[2][13] ),
    .X(_02157_));
 sky130_fd_sc_hd__a22o_1 _05658_ (.A1(\tms1x00.O_pla_ors[2][8] ),
    .A2(_02051_),
    .B1(_02105_),
    .B2(\tms1x00.O_pla_ors[2][4] ),
    .X(_02158_));
 sky130_fd_sc_hd__a22o_1 _05659_ (.A1(\tms1x00.O_pla_ors[2][3] ),
    .A2(_02069_),
    .B1(_02123_),
    .B2(\tms1x00.O_pla_ors[2][12] ),
    .X(_02159_));
 sky130_fd_sc_hd__a22o_1 _05660_ (.A1(\tms1x00.O_pla_ors[2][2] ),
    .A2(_02033_),
    .B1(_02057_),
    .B2(\tms1x00.O_pla_ors[2][11] ),
    .X(_02160_));
 sky130_fd_sc_hd__or4_2 _05661_ (.A(_02157_),
    .B(_02158_),
    .C(_02159_),
    .D(_02160_),
    .X(_02161_));
 sky130_fd_sc_hd__a22o_1 _05662_ (.A1(\tms1x00.O_pla_ors[2][5] ),
    .A2(_02111_),
    .B1(_02129_),
    .B2(\tms1x00.O_pla_ors[2][0] ),
    .X(_02162_));
 sky130_fd_sc_hd__a221o_2 _05663_ (.A1(\tms1x00.O_pla_ors[2][18] ),
    .A2(_02093_),
    .B1(_02135_),
    .B2(\tms1x00.O_pla_ors[2][1] ),
    .C1(_02162_),
    .X(_02163_));
 sky130_fd_sc_hd__a22o_1 _05664_ (.A1(\tms1x00.O_pla_ors[2][16] ),
    .A2(_02081_),
    .B1(_02099_),
    .B2(\tms1x00.O_pla_ors[2][7] ),
    .X(_02164_));
 sky130_fd_sc_hd__a221o_1 _05665_ (.A1(\tms1x00.O_pla_ors[2][15] ),
    .A2(_02063_),
    .B1(_02087_),
    .B2(\tms1x00.O_pla_ors[2][14] ),
    .C1(_02164_),
    .X(_02165_));
 sky130_fd_sc_hd__a22o_1 _05666_ (.A1(\tms1x00.O_pla_ors[2][19] ),
    .A2(_02020_),
    .B1(_02026_),
    .B2(\tms1x00.O_pla_ors[2][10] ),
    .X(_02166_));
 sky130_fd_sc_hd__a221o_2 _05667_ (.A1(\tms1x00.O_pla_ors[2][6] ),
    .A2(_02039_),
    .B1(_02075_),
    .B2(\tms1x00.O_pla_ors[2][9] ),
    .C1(_02166_),
    .X(_02167_));
 sky130_fd_sc_hd__or4_4 _05668_ (.A(_02161_),
    .B(_02163_),
    .C(_02165_),
    .D(_02167_),
    .X(net122));
 sky130_fd_sc_hd__a22o_1 _05669_ (.A1(\tms1x00.O_pla_ors[3][15] ),
    .A2(_02063_),
    .B1(_02087_),
    .B2(\tms1x00.O_pla_ors[3][14] ),
    .X(_02168_));
 sky130_fd_sc_hd__a22o_1 _05670_ (.A1(\tms1x00.O_pla_ors[3][2] ),
    .A2(_02033_),
    .B1(_02057_),
    .B2(\tms1x00.O_pla_ors[3][11] ),
    .X(_02169_));
 sky130_fd_sc_hd__a22o_1 _05671_ (.A1(\tms1x00.O_pla_ors[3][17] ),
    .A2(_02045_),
    .B1(_02117_),
    .B2(\tms1x00.O_pla_ors[3][13] ),
    .X(_02170_));
 sky130_fd_sc_hd__a22o_1 _05672_ (.A1(\tms1x00.O_pla_ors[3][8] ),
    .A2(_02051_),
    .B1(_02105_),
    .B2(\tms1x00.O_pla_ors[3][4] ),
    .X(_02171_));
 sky130_fd_sc_hd__a221o_1 _05673_ (.A1(\tms1x00.O_pla_ors[3][16] ),
    .A2(_02081_),
    .B1(_02099_),
    .B2(\tms1x00.O_pla_ors[3][7] ),
    .C1(_02168_),
    .X(_02172_));
 sky130_fd_sc_hd__a22o_1 _05674_ (.A1(\tms1x00.O_pla_ors[3][19] ),
    .A2(_02020_),
    .B1(_02026_),
    .B2(\tms1x00.O_pla_ors[3][10] ),
    .X(_02173_));
 sky130_fd_sc_hd__a221o_1 _05675_ (.A1(\tms1x00.O_pla_ors[3][6] ),
    .A2(_02039_),
    .B1(_02075_),
    .B2(\tms1x00.O_pla_ors[3][9] ),
    .C1(_02173_),
    .X(_02174_));
 sky130_fd_sc_hd__a22o_1 _05676_ (.A1(\tms1x00.O_pla_ors[3][3] ),
    .A2(_02069_),
    .B1(_02123_),
    .B2(\tms1x00.O_pla_ors[3][12] ),
    .X(_02175_));
 sky130_fd_sc_hd__a22o_1 _05677_ (.A1(\tms1x00.O_pla_ors[3][18] ),
    .A2(_02093_),
    .B1(_02135_),
    .B2(\tms1x00.O_pla_ors[3][1] ),
    .X(_02176_));
 sky130_fd_sc_hd__a221o_1 _05678_ (.A1(\tms1x00.O_pla_ors[3][5] ),
    .A2(_02111_),
    .B1(_02129_),
    .B2(\tms1x00.O_pla_ors[3][0] ),
    .C1(_02176_),
    .X(_02177_));
 sky130_fd_sc_hd__or4_2 _05679_ (.A(_02169_),
    .B(_02170_),
    .C(_02171_),
    .D(_02175_),
    .X(_02178_));
 sky130_fd_sc_hd__or4_4 _05680_ (.A(_02172_),
    .B(_02174_),
    .C(_02177_),
    .D(_02178_),
    .X(net123));
 sky130_fd_sc_hd__a22o_1 _05681_ (.A1(\tms1x00.O_pla_ors[4][17] ),
    .A2(_02045_),
    .B1(_02099_),
    .B2(\tms1x00.O_pla_ors[4][7] ),
    .X(_02179_));
 sky130_fd_sc_hd__a221o_1 _05682_ (.A1(\tms1x00.O_pla_ors[4][2] ),
    .A2(_02033_),
    .B1(_02093_),
    .B2(\tms1x00.O_pla_ors[4][18] ),
    .C1(_02179_),
    .X(_02180_));
 sky130_fd_sc_hd__a22o_1 _05683_ (.A1(\tms1x00.O_pla_ors[4][15] ),
    .A2(_02063_),
    .B1(_02069_),
    .B2(\tms1x00.O_pla_ors[4][3] ),
    .X(_02181_));
 sky130_fd_sc_hd__a221o_1 _05684_ (.A1(\tms1x00.O_pla_ors[4][8] ),
    .A2(_02051_),
    .B1(_02105_),
    .B2(\tms1x00.O_pla_ors[4][4] ),
    .C1(_02181_),
    .X(_02182_));
 sky130_fd_sc_hd__a22o_1 _05685_ (.A1(\tms1x00.O_pla_ors[4][6] ),
    .A2(_02039_),
    .B1(_02135_),
    .B2(\tms1x00.O_pla_ors[4][1] ),
    .X(_02183_));
 sky130_fd_sc_hd__a221o_1 _05686_ (.A1(\tms1x00.O_pla_ors[4][11] ),
    .A2(_02057_),
    .B1(_02129_),
    .B2(\tms1x00.O_pla_ors[4][0] ),
    .C1(_02183_),
    .X(_02184_));
 sky130_fd_sc_hd__a22o_1 _05687_ (.A1(\tms1x00.O_pla_ors[4][10] ),
    .A2(_02026_),
    .B1(_02087_),
    .B2(\tms1x00.O_pla_ors[4][14] ),
    .X(_02185_));
 sky130_fd_sc_hd__a221o_2 _05688_ (.A1(\tms1x00.O_pla_ors[4][9] ),
    .A2(_02075_),
    .B1(_02081_),
    .B2(\tms1x00.O_pla_ors[4][16] ),
    .C1(_02185_),
    .X(_02186_));
 sky130_fd_sc_hd__a22o_1 _05689_ (.A1(\tms1x00.O_pla_ors[4][19] ),
    .A2(_02020_),
    .B1(_02123_),
    .B2(\tms1x00.O_pla_ors[4][12] ),
    .X(_02187_));
 sky130_fd_sc_hd__a221o_1 _05690_ (.A1(\tms1x00.O_pla_ors[4][5] ),
    .A2(_02111_),
    .B1(_02117_),
    .B2(\tms1x00.O_pla_ors[4][13] ),
    .C1(_02187_),
    .X(_02188_));
 sky130_fd_sc_hd__or3_1 _05691_ (.A(_02184_),
    .B(_02186_),
    .C(_02188_),
    .X(_02189_));
 sky130_fd_sc_hd__or3_4 _05692_ (.A(_02180_),
    .B(_02182_),
    .C(_02189_),
    .X(net124));
 sky130_fd_sc_hd__a22o_1 _05693_ (.A1(\tms1x00.O_pla_ors[5][5] ),
    .A2(_02111_),
    .B1(_02129_),
    .B2(\tms1x00.O_pla_ors[5][0] ),
    .X(_02190_));
 sky130_fd_sc_hd__a221o_1 _05694_ (.A1(\tms1x00.O_pla_ors[5][18] ),
    .A2(_02093_),
    .B1(_02135_),
    .B2(\tms1x00.O_pla_ors[5][1] ),
    .C1(_02190_),
    .X(_02191_));
 sky130_fd_sc_hd__a22o_1 _05695_ (.A1(\tms1x00.O_pla_ors[5][19] ),
    .A2(_02020_),
    .B1(_02026_),
    .B2(\tms1x00.O_pla_ors[5][10] ),
    .X(_02192_));
 sky130_fd_sc_hd__a221o_1 _05696_ (.A1(\tms1x00.O_pla_ors[5][6] ),
    .A2(_02039_),
    .B1(_02075_),
    .B2(\tms1x00.O_pla_ors[5][9] ),
    .C1(_02192_),
    .X(_02193_));
 sky130_fd_sc_hd__a22o_1 _05697_ (.A1(\tms1x00.O_pla_ors[5][17] ),
    .A2(_02045_),
    .B1(_02105_),
    .B2(\tms1x00.O_pla_ors[5][4] ),
    .X(_02194_));
 sky130_fd_sc_hd__a221o_1 _05698_ (.A1(\tms1x00.O_pla_ors[5][13] ),
    .A2(_02117_),
    .B1(_02123_),
    .B2(\tms1x00.O_pla_ors[5][12] ),
    .C1(_02194_),
    .X(_02195_));
 sky130_fd_sc_hd__a22o_1 _05699_ (.A1(\tms1x00.O_pla_ors[5][2] ),
    .A2(_02033_),
    .B1(_02069_),
    .B2(\tms1x00.O_pla_ors[5][3] ),
    .X(_02196_));
 sky130_fd_sc_hd__a221o_1 _05700_ (.A1(\tms1x00.O_pla_ors[5][8] ),
    .A2(_02051_),
    .B1(_02057_),
    .B2(\tms1x00.O_pla_ors[5][11] ),
    .C1(_02196_),
    .X(_02197_));
 sky130_fd_sc_hd__a22o_1 _05701_ (.A1(\tms1x00.O_pla_ors[5][16] ),
    .A2(_02081_),
    .B1(_02099_),
    .B2(\tms1x00.O_pla_ors[5][7] ),
    .X(_02198_));
 sky130_fd_sc_hd__a221o_1 _05702_ (.A1(\tms1x00.O_pla_ors[5][15] ),
    .A2(_02063_),
    .B1(_02087_),
    .B2(\tms1x00.O_pla_ors[5][14] ),
    .C1(_02198_),
    .X(_02199_));
 sky130_fd_sc_hd__or3_1 _05703_ (.A(_02195_),
    .B(_02197_),
    .C(_02199_),
    .X(_02200_));
 sky130_fd_sc_hd__or3_4 _05704_ (.A(_02191_),
    .B(_02193_),
    .C(_02200_),
    .X(net125));
 sky130_fd_sc_hd__a22o_1 _05705_ (.A1(\tms1x00.O_pla_ors[6][17] ),
    .A2(_02045_),
    .B1(_02117_),
    .B2(\tms1x00.O_pla_ors[6][13] ),
    .X(_02201_));
 sky130_fd_sc_hd__a22o_1 _05706_ (.A1(\tms1x00.O_pla_ors[6][8] ),
    .A2(_02051_),
    .B1(_02105_),
    .B2(\tms1x00.O_pla_ors[6][4] ),
    .X(_02202_));
 sky130_fd_sc_hd__a22o_1 _05707_ (.A1(\tms1x00.O_pla_ors[6][3] ),
    .A2(_02069_),
    .B1(_02123_),
    .B2(\tms1x00.O_pla_ors[6][12] ),
    .X(_02203_));
 sky130_fd_sc_hd__a22o_1 _05708_ (.A1(\tms1x00.O_pla_ors[6][2] ),
    .A2(_02033_),
    .B1(_02057_),
    .B2(\tms1x00.O_pla_ors[6][11] ),
    .X(_02204_));
 sky130_fd_sc_hd__or4_2 _05709_ (.A(_02201_),
    .B(_02202_),
    .C(_02203_),
    .D(_02204_),
    .X(_02205_));
 sky130_fd_sc_hd__a22o_1 _05710_ (.A1(\tms1x00.O_pla_ors[6][5] ),
    .A2(_02111_),
    .B1(_02129_),
    .B2(\tms1x00.O_pla_ors[6][0] ),
    .X(_02206_));
 sky130_fd_sc_hd__a221o_2 _05711_ (.A1(\tms1x00.O_pla_ors[6][18] ),
    .A2(_02093_),
    .B1(_02135_),
    .B2(\tms1x00.O_pla_ors[6][1] ),
    .C1(_02206_),
    .X(_02207_));
 sky130_fd_sc_hd__a22o_1 _05712_ (.A1(\tms1x00.O_pla_ors[6][19] ),
    .A2(_02020_),
    .B1(_02026_),
    .B2(\tms1x00.O_pla_ors[6][10] ),
    .X(_02208_));
 sky130_fd_sc_hd__a22o_1 _05713_ (.A1(\tms1x00.O_pla_ors[6][16] ),
    .A2(_02081_),
    .B1(_02099_),
    .B2(\tms1x00.O_pla_ors[6][7] ),
    .X(_02209_));
 sky130_fd_sc_hd__a221o_1 _05714_ (.A1(\tms1x00.O_pla_ors[6][15] ),
    .A2(_02063_),
    .B1(_02087_),
    .B2(\tms1x00.O_pla_ors[6][14] ),
    .C1(_02209_),
    .X(_02210_));
 sky130_fd_sc_hd__a221o_2 _05715_ (.A1(\tms1x00.O_pla_ors[6][6] ),
    .A2(_02039_),
    .B1(_02075_),
    .B2(\tms1x00.O_pla_ors[6][9] ),
    .C1(_02208_),
    .X(_02211_));
 sky130_fd_sc_hd__or4_4 _05716_ (.A(_02205_),
    .B(_02207_),
    .C(_02210_),
    .D(_02211_),
    .X(net126));
 sky130_fd_sc_hd__a22o_1 _05717_ (.A1(\tms1x00.O_pla_ors[7][17] ),
    .A2(_02045_),
    .B1(_02117_),
    .B2(\tms1x00.O_pla_ors[7][13] ),
    .X(_02212_));
 sky130_fd_sc_hd__a22o_1 _05718_ (.A1(\tms1x00.O_pla_ors[7][8] ),
    .A2(_02051_),
    .B1(_02105_),
    .B2(\tms1x00.O_pla_ors[7][4] ),
    .X(_02213_));
 sky130_fd_sc_hd__a22o_1 _05719_ (.A1(\tms1x00.O_pla_ors[7][16] ),
    .A2(_02081_),
    .B1(_02099_),
    .B2(\tms1x00.O_pla_ors[7][7] ),
    .X(_02214_));
 sky130_fd_sc_hd__a221o_1 _05720_ (.A1(\tms1x00.O_pla_ors[7][15] ),
    .A2(_02063_),
    .B1(_02087_),
    .B2(\tms1x00.O_pla_ors[7][14] ),
    .C1(_02214_),
    .X(_02215_));
 sky130_fd_sc_hd__a22o_1 _05721_ (.A1(\tms1x00.O_pla_ors[7][19] ),
    .A2(_02020_),
    .B1(_02026_),
    .B2(\tms1x00.O_pla_ors[7][10] ),
    .X(_02216_));
 sky130_fd_sc_hd__a221o_1 _05722_ (.A1(\tms1x00.O_pla_ors[7][6] ),
    .A2(_02039_),
    .B1(_02075_),
    .B2(\tms1x00.O_pla_ors[7][9] ),
    .C1(_02216_),
    .X(_02217_));
 sky130_fd_sc_hd__a22o_1 _05723_ (.A1(\tms1x00.O_pla_ors[7][3] ),
    .A2(_02069_),
    .B1(_02123_),
    .B2(\tms1x00.O_pla_ors[7][12] ),
    .X(_02218_));
 sky130_fd_sc_hd__a22o_1 _05724_ (.A1(\tms1x00.O_pla_ors[7][18] ),
    .A2(_02093_),
    .B1(_02135_),
    .B2(\tms1x00.O_pla_ors[7][1] ),
    .X(_02219_));
 sky130_fd_sc_hd__a221o_2 _05725_ (.A1(\tms1x00.O_pla_ors[7][5] ),
    .A2(_02111_),
    .B1(_02129_),
    .B2(\tms1x00.O_pla_ors[7][0] ),
    .C1(_02219_),
    .X(_02220_));
 sky130_fd_sc_hd__a22o_1 _05726_ (.A1(\tms1x00.O_pla_ors[7][2] ),
    .A2(_02033_),
    .B1(_02057_),
    .B2(\tms1x00.O_pla_ors[7][11] ),
    .X(_02221_));
 sky130_fd_sc_hd__or4_2 _05727_ (.A(_02212_),
    .B(_02213_),
    .C(_02218_),
    .D(_02221_),
    .X(_02222_));
 sky130_fd_sc_hd__or4_4 _05728_ (.A(_02215_),
    .B(_02217_),
    .C(_02220_),
    .D(_02222_),
    .X(net127));
 sky130_fd_sc_hd__and3_4 _05729_ (.A(net118),
    .B(net87),
    .C(net78),
    .X(_02223_));
 sky130_fd_sc_hd__nand2_8 _05730_ (.A(net78),
    .B(valid),
    .Y(_02224_));
 sky130_fd_sc_hd__and2_1 _05731_ (.A(net906),
    .B(\wbs_o_buff[0] ),
    .X(_02225_));
 sky130_fd_sc_hd__nand2_8 _05732_ (.A(net77),
    .B(valid),
    .Y(_02226_));
 sky130_fd_sc_hd__nor2_8 _05733_ (.A(net119),
    .B(_02226_),
    .Y(_02227_));
 sky130_fd_sc_hd__or2_4 _05734_ (.A(net119),
    .B(_02226_),
    .X(_02228_));
 sky130_fd_sc_hd__nand2_4 _05735_ (.A(net1003),
    .B(net1001),
    .Y(_02229_));
 sky130_fd_sc_hd__nor2_8 _05736_ (.A(net1005),
    .B(_02229_),
    .Y(_02230_));
 sky130_fd_sc_hd__or2_4 _05737_ (.A(net1005),
    .B(_02229_),
    .X(_02231_));
 sky130_fd_sc_hd__and3b_2 _05738_ (.A_N(net1003),
    .B(net1001),
    .C(net1005),
    .X(_02232_));
 sky130_fd_sc_hd__nand3b_2 _05739_ (.A_N(net1003),
    .B(net1002),
    .C(net1005),
    .Y(_02233_));
 sky130_fd_sc_hd__and3b_2 _05740_ (.A_N(net1001),
    .B(net1003),
    .C(net1005),
    .X(_02234_));
 sky130_fd_sc_hd__nand3b_4 _05741_ (.A_N(net1001),
    .B(net1003),
    .C(net1005),
    .Y(_02235_));
 sky130_fd_sc_hd__nor3_4 _05742_ (.A(net1005),
    .B(net1003),
    .C(net1001),
    .Y(_02236_));
 sky130_fd_sc_hd__or3_4 _05743_ (.A(net1005),
    .B(net1003),
    .C(net1001),
    .X(_02237_));
 sky130_fd_sc_hd__nor3b_4 _05744_ (.A(net1006),
    .B(net1003),
    .C_N(net1001),
    .Y(_02238_));
 sky130_fd_sc_hd__or3b_4 _05745_ (.A(net1005),
    .B(net1003),
    .C_N(net1001),
    .X(_02239_));
 sky130_fd_sc_hd__and3_4 _05746_ (.A(net1006),
    .B(net1004),
    .C(net1002),
    .X(_02240_));
 sky130_fd_sc_hd__nand3_2 _05747_ (.A(net79),
    .B(net1004),
    .C(net1002),
    .Y(_02241_));
 sky130_fd_sc_hd__nor3b_4 _05748_ (.A(net1004),
    .B(net1002),
    .C_N(net1006),
    .Y(_02242_));
 sky130_fd_sc_hd__or3b_4 _05749_ (.A(net1003),
    .B(net1001),
    .C_N(net1005),
    .X(_02243_));
 sky130_fd_sc_hd__nor3b_4 _05750_ (.A(net1006),
    .B(net1002),
    .C_N(net1004),
    .Y(_02244_));
 sky130_fd_sc_hd__or3b_4 _05751_ (.A(net1006),
    .B(net1001),
    .C_N(net1004),
    .X(_02245_));
 sky130_fd_sc_hd__o22a_1 _05752_ (.A1(\tms1x00.O_pla_ands[6][0] ),
    .A2(net622),
    .B1(net788),
    .B2(\tms1x00.O_pla_ands[7][0] ),
    .X(_02246_));
 sky130_fd_sc_hd__o221a_1 _05753_ (.A1(\tms1x00.O_pla_ands[0][0] ),
    .A2(net834),
    .B1(net754),
    .B2(\tms1x00.O_pla_ands[1][0] ),
    .C1(net915),
    .X(_02247_));
 sky130_fd_sc_hd__o22a_1 _05754_ (.A1(\tms1x00.O_pla_ands[3][0] ),
    .A2(net868),
    .B1(net734),
    .B2(\tms1x00.O_pla_ands[2][0] ),
    .X(_02248_));
 sky130_fd_sc_hd__o211a_1 _05755_ (.A1(\tms1x00.O_pla_ands[5][0] ),
    .A2(net896),
    .B1(_02247_),
    .C1(_02248_),
    .X(_02249_));
 sky130_fd_sc_hd__o211a_1 _05756_ (.A1(\tms1x00.O_pla_ands[4][0] ),
    .A2(net814),
    .B1(_02246_),
    .C1(_02249_),
    .X(_02250_));
 sky130_fd_sc_hd__o22a_1 _05757_ (.A1(\tms1x00.O_pla_ands[13][0] ),
    .A2(net897),
    .B1(net765),
    .B2(\tms1x00.O_pla_ands[9][0] ),
    .X(_02251_));
 sky130_fd_sc_hd__o22a_1 _05758_ (.A1(\tms1x00.O_pla_ands[8][0] ),
    .A2(net843),
    .B1(net791),
    .B2(\tms1x00.O_pla_ands[15][0] ),
    .X(_02252_));
 sky130_fd_sc_hd__o221a_2 _05759_ (.A1(\tms1x00.O_pla_ands[12][0] ),
    .A2(net817),
    .B1(net735),
    .B2(\tms1x00.O_pla_ands[10][0] ),
    .C1(_02252_),
    .X(_02253_));
 sky130_fd_sc_hd__o211a_1 _05760_ (.A1(\tms1x00.O_pla_ands[11][0] ),
    .A2(net869),
    .B1(_02253_),
    .C1(net999),
    .X(_02254_));
 sky130_fd_sc_hd__o211a_1 _05761_ (.A1(\tms1x00.O_pla_ands[14][0] ),
    .A2(net623),
    .B1(_02251_),
    .C1(_02254_),
    .X(_02255_));
 sky130_fd_sc_hd__or3_2 _05762_ (.A(net988),
    .B(_02250_),
    .C(_02255_),
    .X(_02256_));
 sky130_fd_sc_hd__o22a_1 _05763_ (.A1(\tms1x00.O_pla_ands[30][0] ),
    .A2(net611),
    .B1(net777),
    .B2(\tms1x00.O_pla_ands[31][0] ),
    .X(_02257_));
 sky130_fd_sc_hd__o22a_1 _05764_ (.A1(\tms1x00.O_pla_ands[27][0] ),
    .A2(net855),
    .B1(net722),
    .B2(\tms1x00.O_pla_ands[26][0] ),
    .X(_02258_));
 sky130_fd_sc_hd__o221a_1 _05765_ (.A1(\tms1x00.O_pla_ands[29][0] ),
    .A2(net884),
    .B1(net803),
    .B2(\tms1x00.O_pla_ands[28][0] ),
    .C1(net992),
    .X(_02259_));
 sky130_fd_sc_hd__o211a_1 _05766_ (.A1(\tms1x00.O_pla_ands[25][0] ),
    .A2(net748),
    .B1(_02258_),
    .C1(_02259_),
    .X(_02260_));
 sky130_fd_sc_hd__o211a_4 _05767_ (.A1(\tms1x00.O_pla_ands[24][0] ),
    .A2(net830),
    .B1(_02257_),
    .C1(_02260_),
    .X(_02261_));
 sky130_fd_sc_hd__o22a_2 _05768_ (.A1(\tms1x00.O_pla_ands[22][0] ),
    .A2(net610),
    .B1(net776),
    .B2(\tms1x00.O_pla_ands[23][0] ),
    .X(_02262_));
 sky130_fd_sc_hd__o221a_1 _05769_ (.A1(\tms1x00.O_pla_ands[16][0] ),
    .A2(net834),
    .B1(net752),
    .B2(\tms1x00.O_pla_ands[17][0] ),
    .C1(net915),
    .X(_02263_));
 sky130_fd_sc_hd__o22a_1 _05770_ (.A1(\tms1x00.O_pla_ands[19][0] ),
    .A2(net860),
    .B1(net724),
    .B2(\tms1x00.O_pla_ands[18][0] ),
    .X(_02264_));
 sky130_fd_sc_hd__o211a_1 _05771_ (.A1(\tms1x00.O_pla_ands[21][0] ),
    .A2(net885),
    .B1(_02263_),
    .C1(_02264_),
    .X(_02265_));
 sky130_fd_sc_hd__o211a_1 _05772_ (.A1(\tms1x00.O_pla_ands[20][0] ),
    .A2(net805),
    .B1(_02262_),
    .C1(_02265_),
    .X(_02266_));
 sky130_fd_sc_hd__o311a_2 _05773_ (.A1(net925),
    .A2(_02261_),
    .A3(_02266_),
    .B1(net905),
    .C1(_02256_),
    .X(_02267_));
 sky130_fd_sc_hd__nor2_4 _05774_ (.A(net905),
    .B(net984),
    .Y(_02268_));
 sky130_fd_sc_hd__o22a_1 _05775_ (.A1(\tms1x00.ins_pla_ors[11][0] ),
    .A2(net852),
    .B1(net717),
    .B2(\tms1x00.ins_pla_ors[10][0] ),
    .X(_02269_));
 sky130_fd_sc_hd__o22a_1 _05776_ (.A1(\tms1x00.ins_pla_ors[12][0] ),
    .A2(net799),
    .B1(net772),
    .B2(\tms1x00.ins_pla_ors[15][0] ),
    .X(_02270_));
 sky130_fd_sc_hd__o221a_1 _05777_ (.A1(\tms1x00.ins_pla_ors[14][0] ),
    .A2(net605),
    .B1(net827),
    .B2(\tms1x00.ins_pla_ors[8][0] ),
    .C1(_02270_),
    .X(_02271_));
 sky130_fd_sc_hd__o211a_1 _05778_ (.A1(\tms1x00.ins_pla_ors[9][0] ),
    .A2(net745),
    .B1(_02271_),
    .C1(net996),
    .X(_02272_));
 sky130_fd_sc_hd__o211a_1 _05779_ (.A1(\tms1x00.ins_pla_ors[13][0] ),
    .A2(net880),
    .B1(_02269_),
    .C1(_02272_),
    .X(_02273_));
 sky130_fd_sc_hd__o22a_1 _05780_ (.A1(\tms1x00.ins_pla_ors[3][0] ),
    .A2(net866),
    .B1(net759),
    .B2(\tms1x00.ins_pla_ors[1][0] ),
    .X(_02274_));
 sky130_fd_sc_hd__o22a_1 _05781_ (.A1(\tms1x00.ins_pla_ors[7][0] ),
    .A2(net786),
    .B1(net730),
    .B2(\tms1x00.ins_pla_ors[2][0] ),
    .X(_02275_));
 sky130_fd_sc_hd__o221a_1 _05782_ (.A1(\tms1x00.ins_pla_ors[0][0] ),
    .A2(net840),
    .B1(net810),
    .B2(\tms1x00.ins_pla_ors[4][0] ),
    .C1(_02275_),
    .X(_02276_));
 sky130_fd_sc_hd__o211a_1 _05783_ (.A1(\tms1x00.ins_pla_ors[5][0] ),
    .A2(net893),
    .B1(_02276_),
    .C1(net919),
    .X(_02277_));
 sky130_fd_sc_hd__o211a_4 _05784_ (.A1(\tms1x00.ins_pla_ors[6][0] ),
    .A2(net620),
    .B1(_02274_),
    .C1(_02277_),
    .X(_02278_));
 sky130_fd_sc_hd__o21a_1 _05785_ (.A1(_02273_),
    .A2(_02278_),
    .B1(net600),
    .X(_02279_));
 sky130_fd_sc_hd__nor2_1 _05786_ (.A(net985),
    .B(net984),
    .Y(_02280_));
 sky130_fd_sc_hd__or2_2 _05787_ (.A(net985),
    .B(net984),
    .X(_02281_));
 sky130_fd_sc_hd__o22a_1 _05788_ (.A1(\tms1x00.O_pla_ors[3][0] ),
    .A2(net872),
    .B1(net816),
    .B2(\tms1x00.O_pla_ors[4][0] ),
    .X(_02282_));
 sky130_fd_sc_hd__nor2_8 _05789_ (.A(net905),
    .B(_01637_),
    .Y(_02283_));
 sky130_fd_sc_hd__o22a_1 _05790_ (.A1(\tms1x00.O_pla_ors[7][0] ),
    .A2(net790),
    .B1(net763),
    .B2(\tms1x00.O_pla_ors[1][0] ),
    .X(_02284_));
 sky130_fd_sc_hd__o221a_1 _05791_ (.A1(\tms1x00.O_pla_ors[0][0] ),
    .A2(net843),
    .B1(net736),
    .B2(\tms1x00.O_pla_ors[2][0] ),
    .C1(_02284_),
    .X(_02285_));
 sky130_fd_sc_hd__o211a_1 _05792_ (.A1(\tms1x00.O_pla_ors[5][0] ),
    .A2(net899),
    .B1(_02283_),
    .C1(_02285_),
    .X(_02286_));
 sky130_fd_sc_hd__o211a_4 _05793_ (.A1(\tms1x00.O_pla_ors[6][0] ),
    .A2(net624),
    .B1(_02282_),
    .C1(_02286_),
    .X(_02287_));
 sky130_fd_sc_hd__o22a_1 _05794_ (.A1(\tms1x00.ins_pla_ands[28][0] ),
    .A2(net798),
    .B1(net772),
    .B2(\tms1x00.ins_pla_ands[31][0] ),
    .X(_02288_));
 sky130_fd_sc_hd__o22a_1 _05795_ (.A1(\tms1x00.ins_pla_ands[29][0] ),
    .A2(net879),
    .B1(net827),
    .B2(\tms1x00.ins_pla_ands[24][0] ),
    .X(_02289_));
 sky130_fd_sc_hd__o221a_1 _05796_ (.A1(\tms1x00.ins_pla_ands[25][0] ),
    .A2(net745),
    .B1(net717),
    .B2(\tms1x00.ins_pla_ands[26][0] ),
    .C1(_02289_),
    .X(_02290_));
 sky130_fd_sc_hd__o211a_1 _05797_ (.A1(\tms1x00.ins_pla_ands[27][0] ),
    .A2(net852),
    .B1(_02290_),
    .C1(net990),
    .X(_02291_));
 sky130_fd_sc_hd__o211a_1 _05798_ (.A1(\tms1x00.ins_pla_ands[30][0] ),
    .A2(net605),
    .B1(_02288_),
    .C1(_02291_),
    .X(_02292_));
 sky130_fd_sc_hd__o22a_1 _05799_ (.A1(\tms1x00.ins_pla_ands[22][0] ),
    .A2(net604),
    .B1(net771),
    .B2(\tms1x00.ins_pla_ands[23][0] ),
    .X(_02293_));
 sky130_fd_sc_hd__o221a_2 _05800_ (.A1(\tms1x00.ins_pla_ands[21][0] ),
    .A2(net878),
    .B1(net797),
    .B2(\tms1x00.ins_pla_ands[20][0] ),
    .C1(net911),
    .X(_02294_));
 sky130_fd_sc_hd__o22a_1 _05801_ (.A1(\tms1x00.ins_pla_ands[19][0] ),
    .A2(net853),
    .B1(net718),
    .B2(\tms1x00.ins_pla_ands[18][0] ),
    .X(_02295_));
 sky130_fd_sc_hd__o211a_1 _05802_ (.A1(\tms1x00.ins_pla_ands[16][0] ),
    .A2(net827),
    .B1(_02294_),
    .C1(_02295_),
    .X(_02296_));
 sky130_fd_sc_hd__o211a_1 _05803_ (.A1(\tms1x00.ins_pla_ands[17][0] ),
    .A2(net746),
    .B1(_02293_),
    .C1(_02296_),
    .X(_02297_));
 sky130_fd_sc_hd__o22a_1 _05804_ (.A1(\tms1x00.ins_pla_ands[3][0] ),
    .A2(net859),
    .B1(net725),
    .B2(\tms1x00.ins_pla_ands[2][0] ),
    .X(_02298_));
 sky130_fd_sc_hd__o221a_1 _05805_ (.A1(\tms1x00.ins_pla_ands[6][0] ),
    .A2(net613),
    .B1(net751),
    .B2(\tms1x00.ins_pla_ands[1][0] ),
    .C1(_02298_),
    .X(_02299_));
 sky130_fd_sc_hd__o221a_2 _05806_ (.A1(\tms1x00.ins_pla_ands[5][0] ),
    .A2(net894),
    .B1(net812),
    .B2(\tms1x00.ins_pla_ands[4][0] ),
    .C1(net921),
    .X(_02300_));
 sky130_fd_sc_hd__o221a_1 _05807_ (.A1(\tms1x00.ins_pla_ands[0][0] ),
    .A2(net832),
    .B1(net780),
    .B2(\tms1x00.ins_pla_ands[7][0] ),
    .C1(_02300_),
    .X(_02301_));
 sky130_fd_sc_hd__o22a_1 _05808_ (.A1(\tms1x00.ins_pla_ands[14][0] ),
    .A2(net608),
    .B1(net779),
    .B2(\tms1x00.ins_pla_ands[15][0] ),
    .X(_02302_));
 sky130_fd_sc_hd__o221a_1 _05809_ (.A1(\tms1x00.ins_pla_ands[13][0] ),
    .A2(net882),
    .B1(net801),
    .B2(\tms1x00.ins_pla_ands[12][0] ),
    .C1(net993),
    .X(_02303_));
 sky130_fd_sc_hd__o22a_1 _05810_ (.A1(\tms1x00.ins_pla_ands[11][0] ),
    .A2(net854),
    .B1(net720),
    .B2(\tms1x00.ins_pla_ands[10][0] ),
    .X(_02304_));
 sky130_fd_sc_hd__o211a_1 _05811_ (.A1(\tms1x00.ins_pla_ands[8][0] ),
    .A2(net829),
    .B1(_02303_),
    .C1(_02304_),
    .X(_02305_));
 sky130_fd_sc_hd__o211a_1 _05812_ (.A1(\tms1x00.ins_pla_ands[9][0] ),
    .A2(net747),
    .B1(_02302_),
    .C1(_02305_),
    .X(_02306_));
 sky130_fd_sc_hd__a211o_1 _05813_ (.A1(_02299_),
    .A2(_02301_),
    .B1(_02306_),
    .C1(net986),
    .X(_02307_));
 sky130_fd_sc_hd__o31a_1 _05814_ (.A1(_02267_),
    .A2(_02279_),
    .A3(_02287_),
    .B1(net711),
    .X(_02308_));
 sky130_fd_sc_hd__o311a_1 _05815_ (.A1(net923),
    .A2(_02292_),
    .A3(_02297_),
    .B1(_02307_),
    .C1(net712),
    .X(_02309_));
 sky130_fd_sc_hd__or3_1 _05816_ (.A(net586),
    .B(_02308_),
    .C(_02309_),
    .X(_02310_));
 sky130_fd_sc_hd__o211a_1 _05817_ (.A1(_02225_),
    .A2(net589),
    .B1(_02310_),
    .C1(net629),
    .X(_02311_));
 sky130_fd_sc_hd__nor2_8 _05818_ (.A(net178),
    .B(net630),
    .Y(_02312_));
 sky130_fd_sc_hd__nor2_8 _05819_ (.A(net119),
    .B(net630),
    .Y(_02313_));
 sky130_fd_sc_hd__nand2_8 _05820_ (.A(net178),
    .B(_02223_),
    .Y(_02314_));
 sky130_fd_sc_hd__a221o_1 _05821_ (.A1(_02225_),
    .A2(net583),
    .B1(net579),
    .B2(net120),
    .C1(_02311_),
    .X(_00005_));
 sky130_fd_sc_hd__and2_1 _05822_ (.A(net906),
    .B(\wbs_o_buff[1] ),
    .X(_02315_));
 sky130_fd_sc_hd__o22a_1 _05823_ (.A1(\tms1x00.O_pla_ands[5][1] ),
    .A2(net896),
    .B1(net733),
    .B2(\tms1x00.O_pla_ands[2][1] ),
    .X(_02316_));
 sky130_fd_sc_hd__o221a_1 _05824_ (.A1(\tms1x00.O_pla_ands[6][1] ),
    .A2(net622),
    .B1(net788),
    .B2(\tms1x00.O_pla_ands[7][1] ),
    .C1(_02316_),
    .X(_02317_));
 sky130_fd_sc_hd__o221a_1 _05825_ (.A1(\tms1x00.O_pla_ands[0][1] ),
    .A2(net836),
    .B1(net754),
    .B2(\tms1x00.O_pla_ands[1][1] ),
    .C1(net914),
    .X(_02318_));
 sky130_fd_sc_hd__o221a_1 _05826_ (.A1(\tms1x00.O_pla_ands[3][1] ),
    .A2(net868),
    .B1(net813),
    .B2(\tms1x00.O_pla_ands[4][1] ),
    .C1(_02318_),
    .X(_02319_));
 sky130_fd_sc_hd__o22a_1 _05827_ (.A1(\tms1x00.O_pla_ands[11][1] ),
    .A2(net871),
    .B1(net816),
    .B2(\tms1x00.O_pla_ands[12][1] ),
    .X(_02320_));
 sky130_fd_sc_hd__o221a_1 _05828_ (.A1(\tms1x00.O_pla_ands[8][1] ),
    .A2(net842),
    .B1(net762),
    .B2(\tms1x00.O_pla_ands[9][1] ),
    .C1(net999),
    .X(_02321_));
 sky130_fd_sc_hd__o22a_1 _05829_ (.A1(\tms1x00.O_pla_ands[13][1] ),
    .A2(net898),
    .B1(net736),
    .B2(\tms1x00.O_pla_ands[10][1] ),
    .X(_02322_));
 sky130_fd_sc_hd__o221a_1 _05830_ (.A1(\tms1x00.O_pla_ands[14][1] ),
    .A2(net624),
    .B1(net790),
    .B2(\tms1x00.O_pla_ands[15][1] ),
    .C1(_02322_),
    .X(_02323_));
 sky130_fd_sc_hd__a31o_1 _05831_ (.A1(_02320_),
    .A2(_02321_),
    .A3(_02323_),
    .B1(net988),
    .X(_02324_));
 sky130_fd_sc_hd__a21o_1 _05832_ (.A1(_02317_),
    .A2(_02319_),
    .B1(_02324_),
    .X(_02325_));
 sky130_fd_sc_hd__o22a_1 _05833_ (.A1(\tms1x00.O_pla_ands[24][1] ),
    .A2(net831),
    .B1(net775),
    .B2(\tms1x00.O_pla_ands[31][1] ),
    .X(_02326_));
 sky130_fd_sc_hd__o221a_1 _05834_ (.A1(\tms1x00.O_pla_ands[29][1] ),
    .A2(net884),
    .B1(net803),
    .B2(\tms1x00.O_pla_ands[28][1] ),
    .C1(net992),
    .X(_02327_));
 sky130_fd_sc_hd__o22a_1 _05835_ (.A1(\tms1x00.O_pla_ands[27][1] ),
    .A2(net856),
    .B1(net723),
    .B2(\tms1x00.O_pla_ands[26][1] ),
    .X(_02328_));
 sky130_fd_sc_hd__o221a_1 _05836_ (.A1(\tms1x00.O_pla_ands[30][1] ),
    .A2(net611),
    .B1(net748),
    .B2(\tms1x00.O_pla_ands[25][1] ),
    .C1(_02328_),
    .X(_02329_));
 sky130_fd_sc_hd__o22a_1 _05837_ (.A1(\tms1x00.O_pla_ands[22][1] ),
    .A2(net610),
    .B1(net775),
    .B2(\tms1x00.O_pla_ands[23][1] ),
    .X(_02330_));
 sky130_fd_sc_hd__o221a_1 _05838_ (.A1(\tms1x00.O_pla_ands[16][1] ),
    .A2(net835),
    .B1(net753),
    .B2(\tms1x00.O_pla_ands[17][1] ),
    .C1(net914),
    .X(_02331_));
 sky130_fd_sc_hd__o22a_1 _05839_ (.A1(\tms1x00.O_pla_ands[19][1] ),
    .A2(net858),
    .B1(net724),
    .B2(\tms1x00.O_pla_ands[18][1] ),
    .X(_02332_));
 sky130_fd_sc_hd__o211a_1 _05840_ (.A1(\tms1x00.O_pla_ands[21][1] ),
    .A2(net885),
    .B1(_02331_),
    .C1(_02332_),
    .X(_02333_));
 sky130_fd_sc_hd__o211a_1 _05841_ (.A1(\tms1x00.O_pla_ands[20][1] ),
    .A2(net804),
    .B1(_02330_),
    .C1(_02333_),
    .X(_02334_));
 sky130_fd_sc_hd__a31o_4 _05842_ (.A1(_02326_),
    .A2(_02327_),
    .A3(_02329_),
    .B1(_02334_),
    .X(_02335_));
 sky130_fd_sc_hd__o211a_1 _05843_ (.A1(net925),
    .A2(_02335_),
    .B1(_02325_),
    .C1(_01636_),
    .X(_02336_));
 sky130_fd_sc_hd__o22a_1 _05844_ (.A1(\tms1x00.ins_pla_ors[11][1] ),
    .A2(net853),
    .B1(net719),
    .B2(\tms1x00.ins_pla_ors[10][1] ),
    .X(_02337_));
 sky130_fd_sc_hd__o22a_1 _05845_ (.A1(\tms1x00.ins_pla_ors[12][1] ),
    .A2(net799),
    .B1(net773),
    .B2(\tms1x00.ins_pla_ors[15][1] ),
    .X(_02338_));
 sky130_fd_sc_hd__o221a_1 _05846_ (.A1(\tms1x00.ins_pla_ors[14][1] ),
    .A2(net605),
    .B1(net828),
    .B2(\tms1x00.ins_pla_ors[8][1] ),
    .C1(_02338_),
    .X(_02339_));
 sky130_fd_sc_hd__o211a_1 _05847_ (.A1(\tms1x00.ins_pla_ors[9][1] ),
    .A2(net757),
    .B1(_02339_),
    .C1(net996),
    .X(_02340_));
 sky130_fd_sc_hd__o211a_2 _05848_ (.A1(\tms1x00.ins_pla_ors[13][1] ),
    .A2(net890),
    .B1(_02337_),
    .C1(_02340_),
    .X(_02341_));
 sky130_fd_sc_hd__or2_1 _05849_ (.A(\tms1x00.ins_pla_ors[1][1] ),
    .B(net759),
    .X(_02342_));
 sky130_fd_sc_hd__or2_1 _05850_ (.A(\tms1x00.ins_pla_ors[0][1] ),
    .B(net840),
    .X(_02343_));
 sky130_fd_sc_hd__o221a_1 _05851_ (.A1(\tms1x00.ins_pla_ors[5][1] ),
    .A2(net890),
    .B1(net807),
    .B2(\tms1x00.ins_pla_ors[4][1] ),
    .C1(net920),
    .X(_02344_));
 sky130_fd_sc_hd__o221a_2 _05852_ (.A1(\tms1x00.ins_pla_ors[6][1] ),
    .A2(net620),
    .B1(net786),
    .B2(\tms1x00.ins_pla_ors[7][1] ),
    .C1(_02342_),
    .X(_02345_));
 sky130_fd_sc_hd__o221a_1 _05853_ (.A1(\tms1x00.ins_pla_ors[3][1] ),
    .A2(net866),
    .B1(net730),
    .B2(\tms1x00.ins_pla_ors[2][1] ),
    .C1(_02343_),
    .X(_02346_));
 sky130_fd_sc_hd__a31o_2 _05854_ (.A1(_02344_),
    .A2(_02345_),
    .A3(_02346_),
    .B1(_02341_),
    .X(_02347_));
 sky130_fd_sc_hd__o22a_1 _05855_ (.A1(\tms1x00.O_pla_ors[3][1] ),
    .A2(net873),
    .B1(net736),
    .B2(\tms1x00.O_pla_ors[2][1] ),
    .X(_02348_));
 sky130_fd_sc_hd__o221a_1 _05856_ (.A1(\tms1x00.O_pla_ors[0][1] ),
    .A2(net843),
    .B1(net763),
    .B2(\tms1x00.O_pla_ors[1][1] ),
    .C1(net599),
    .X(_02349_));
 sky130_fd_sc_hd__o22a_1 _05857_ (.A1(\tms1x00.O_pla_ors[6][1] ),
    .A2(net625),
    .B1(net791),
    .B2(\tms1x00.O_pla_ors[7][1] ),
    .X(_02350_));
 sky130_fd_sc_hd__o211a_1 _05858_ (.A1(\tms1x00.O_pla_ors[4][1] ),
    .A2(net817),
    .B1(_02349_),
    .C1(_02350_),
    .X(_02351_));
 sky130_fd_sc_hd__o211a_4 _05859_ (.A1(\tms1x00.O_pla_ors[5][1] ),
    .A2(net899),
    .B1(_02348_),
    .C1(_02351_),
    .X(_02352_));
 sky130_fd_sc_hd__o22a_1 _05860_ (.A1(\tms1x00.ins_pla_ands[19][1] ),
    .A2(net853),
    .B1(net718),
    .B2(\tms1x00.ins_pla_ands[18][1] ),
    .X(_02353_));
 sky130_fd_sc_hd__o22a_1 _05861_ (.A1(\tms1x00.ins_pla_ands[16][1] ),
    .A2(net825),
    .B1(net771),
    .B2(\tms1x00.ins_pla_ands[23][1] ),
    .X(_02354_));
 sky130_fd_sc_hd__o221a_1 _05862_ (.A1(\tms1x00.ins_pla_ands[21][1] ),
    .A2(net878),
    .B1(net797),
    .B2(\tms1x00.ins_pla_ands[20][1] ),
    .C1(net912),
    .X(_02355_));
 sky130_fd_sc_hd__o221a_1 _05863_ (.A1(\tms1x00.ins_pla_ands[22][1] ),
    .A2(net604),
    .B1(net744),
    .B2(\tms1x00.ins_pla_ands[17][1] ),
    .C1(_02353_),
    .X(_02356_));
 sky130_fd_sc_hd__and3_1 _05864_ (.A(_02354_),
    .B(_02355_),
    .C(_02356_),
    .X(_02357_));
 sky130_fd_sc_hd__or2_1 _05865_ (.A(\tms1x00.ins_pla_ands[31][1] ),
    .B(net769),
    .X(_02358_));
 sky130_fd_sc_hd__o221a_1 _05866_ (.A1(\tms1x00.ins_pla_ands[30][1] ),
    .A2(net603),
    .B1(net877),
    .B2(\tms1x00.ins_pla_ands[29][1] ),
    .C1(_02358_),
    .X(_02359_));
 sky130_fd_sc_hd__o22a_1 _05867_ (.A1(\tms1x00.ins_pla_ands[28][1] ),
    .A2(net798),
    .B1(net743),
    .B2(\tms1x00.ins_pla_ands[25][1] ),
    .X(_02360_));
 sky130_fd_sc_hd__o221a_1 _05868_ (.A1(\tms1x00.ins_pla_ands[24][1] ),
    .A2(net823),
    .B1(net716),
    .B2(\tms1x00.ins_pla_ands[26][1] ),
    .C1(_02360_),
    .X(_02361_));
 sky130_fd_sc_hd__o211a_1 _05869_ (.A1(\tms1x00.ins_pla_ands[27][1] ),
    .A2(net850),
    .B1(_02361_),
    .C1(net990),
    .X(_02362_));
 sky130_fd_sc_hd__a211o_2 _05870_ (.A1(_02359_),
    .A2(_02362_),
    .B1(net923),
    .C1(_02357_),
    .X(_02363_));
 sky130_fd_sc_hd__o22a_1 _05871_ (.A1(\tms1x00.ins_pla_ands[6][1] ),
    .A2(net614),
    .B1(net750),
    .B2(\tms1x00.ins_pla_ands[1][1] ),
    .X(_02364_));
 sky130_fd_sc_hd__o22a_1 _05872_ (.A1(\tms1x00.ins_pla_ands[3][1] ),
    .A2(net870),
    .B1(net815),
    .B2(\tms1x00.ins_pla_ands[4][1] ),
    .X(_02365_));
 sky130_fd_sc_hd__o221a_2 _05873_ (.A1(\tms1x00.ins_pla_ands[5][1] ),
    .A2(net894),
    .B1(net732),
    .B2(\tms1x00.ins_pla_ands[2][1] ),
    .C1(_02365_),
    .X(_02366_));
 sky130_fd_sc_hd__o211a_1 _05874_ (.A1(\tms1x00.ins_pla_ands[7][1] ),
    .A2(net779),
    .B1(_02366_),
    .C1(net916),
    .X(_02367_));
 sky130_fd_sc_hd__o211a_1 _05875_ (.A1(\tms1x00.ins_pla_ands[0][1] ),
    .A2(net832),
    .B1(_02364_),
    .C1(_02367_),
    .X(_02368_));
 sky130_fd_sc_hd__o22a_1 _05876_ (.A1(\tms1x00.ins_pla_ands[14][1] ),
    .A2(net609),
    .B1(net779),
    .B2(\tms1x00.ins_pla_ands[15][1] ),
    .X(_02369_));
 sky130_fd_sc_hd__o221a_1 _05877_ (.A1(\tms1x00.ins_pla_ands[13][1] ),
    .A2(net882),
    .B1(net801),
    .B2(\tms1x00.ins_pla_ands[12][1] ),
    .C1(net993),
    .X(_02370_));
 sky130_fd_sc_hd__o22a_1 _05878_ (.A1(\tms1x00.ins_pla_ands[11][1] ),
    .A2(net854),
    .B1(net720),
    .B2(\tms1x00.ins_pla_ands[10][1] ),
    .X(_02371_));
 sky130_fd_sc_hd__o211a_1 _05879_ (.A1(\tms1x00.ins_pla_ands[9][1] ),
    .A2(net747),
    .B1(_02370_),
    .C1(_02371_),
    .X(_02372_));
 sky130_fd_sc_hd__o211a_1 _05880_ (.A1(\tms1x00.ins_pla_ands[8][1] ),
    .A2(net832),
    .B1(_02369_),
    .C1(_02372_),
    .X(_02373_));
 sky130_fd_sc_hd__a211o_2 _05881_ (.A1(net600),
    .A2(_02347_),
    .B1(_02352_),
    .C1(_02336_),
    .X(_02374_));
 sky130_fd_sc_hd__o311a_1 _05882_ (.A1(net986),
    .A2(_02368_),
    .A3(_02373_),
    .B1(net712),
    .C1(_02363_),
    .X(_02375_));
 sky130_fd_sc_hd__a211o_1 _05883_ (.A1(net711),
    .A2(_02374_),
    .B1(_02375_),
    .C1(net586),
    .X(_02376_));
 sky130_fd_sc_hd__o211a_1 _05884_ (.A1(net589),
    .A2(_02315_),
    .B1(_02376_),
    .C1(net629),
    .X(_02377_));
 sky130_fd_sc_hd__a221o_1 _05885_ (.A1(net121),
    .A2(net579),
    .B1(_02315_),
    .B2(net583),
    .C1(_02377_),
    .X(_00016_));
 sky130_fd_sc_hd__and2_1 _05886_ (.A(net906),
    .B(\wbs_o_buff[2] ),
    .X(_02378_));
 sky130_fd_sc_hd__o22a_1 _05887_ (.A1(\tms1x00.O_pla_ands[6][2] ),
    .A2(net622),
    .B1(net788),
    .B2(\tms1x00.O_pla_ands[7][2] ),
    .X(_02379_));
 sky130_fd_sc_hd__o221a_1 _05888_ (.A1(\tms1x00.O_pla_ands[0][2] ),
    .A2(net834),
    .B1(net752),
    .B2(\tms1x00.O_pla_ands[1][2] ),
    .C1(net914),
    .X(_02380_));
 sky130_fd_sc_hd__o22a_1 _05889_ (.A1(\tms1x00.O_pla_ands[3][2] ),
    .A2(net868),
    .B1(net733),
    .B2(\tms1x00.O_pla_ands[2][2] ),
    .X(_02381_));
 sky130_fd_sc_hd__o211a_1 _05890_ (.A1(\tms1x00.O_pla_ands[5][2] ),
    .A2(net896),
    .B1(_02380_),
    .C1(_02381_),
    .X(_02382_));
 sky130_fd_sc_hd__o211a_1 _05891_ (.A1(\tms1x00.O_pla_ands[4][2] ),
    .A2(net813),
    .B1(_02379_),
    .C1(_02382_),
    .X(_02383_));
 sky130_fd_sc_hd__o22a_1 _05892_ (.A1(\tms1x00.O_pla_ands[11][2] ),
    .A2(net871),
    .B1(net816),
    .B2(\tms1x00.O_pla_ands[12][2] ),
    .X(_02384_));
 sky130_fd_sc_hd__o221a_1 _05893_ (.A1(\tms1x00.O_pla_ands[8][2] ),
    .A2(net842),
    .B1(net762),
    .B2(\tms1x00.O_pla_ands[9][2] ),
    .C1(net999),
    .X(_02385_));
 sky130_fd_sc_hd__o22a_1 _05894_ (.A1(\tms1x00.O_pla_ands[13][2] ),
    .A2(net898),
    .B1(net735),
    .B2(\tms1x00.O_pla_ands[10][2] ),
    .X(_02386_));
 sky130_fd_sc_hd__o221a_1 _05895_ (.A1(\tms1x00.O_pla_ands[14][2] ),
    .A2(net624),
    .B1(net790),
    .B2(\tms1x00.O_pla_ands[15][2] ),
    .C1(_02386_),
    .X(_02387_));
 sky130_fd_sc_hd__a31o_2 _05896_ (.A1(_02384_),
    .A2(_02385_),
    .A3(_02387_),
    .B1(net988),
    .X(_02388_));
 sky130_fd_sc_hd__o22a_1 _05897_ (.A1(\tms1x00.O_pla_ands[30][2] ),
    .A2(net611),
    .B1(net775),
    .B2(\tms1x00.O_pla_ands[31][2] ),
    .X(_02389_));
 sky130_fd_sc_hd__o22a_1 _05898_ (.A1(\tms1x00.O_pla_ands[27][2] ),
    .A2(net856),
    .B1(net722),
    .B2(\tms1x00.O_pla_ands[26][2] ),
    .X(_02390_));
 sky130_fd_sc_hd__o221a_1 _05899_ (.A1(\tms1x00.O_pla_ands[29][2] ),
    .A2(net884),
    .B1(net803),
    .B2(\tms1x00.O_pla_ands[28][2] ),
    .C1(net992),
    .X(_02391_));
 sky130_fd_sc_hd__o211a_1 _05900_ (.A1(\tms1x00.O_pla_ands[25][2] ),
    .A2(net748),
    .B1(_02390_),
    .C1(_02391_),
    .X(_02392_));
 sky130_fd_sc_hd__o211a_1 _05901_ (.A1(\tms1x00.O_pla_ands[24][2] ),
    .A2(net830),
    .B1(_02389_),
    .C1(_02392_),
    .X(_02393_));
 sky130_fd_sc_hd__o22a_1 _05902_ (.A1(\tms1x00.O_pla_ands[21][2] ),
    .A2(net885),
    .B1(net723),
    .B2(\tms1x00.O_pla_ands[18][2] ),
    .X(_02394_));
 sky130_fd_sc_hd__o221a_1 _05903_ (.A1(\tms1x00.O_pla_ands[22][2] ),
    .A2(net612),
    .B1(net776),
    .B2(\tms1x00.O_pla_ands[23][2] ),
    .C1(_02394_),
    .X(_02395_));
 sky130_fd_sc_hd__o221a_1 _05904_ (.A1(\tms1x00.O_pla_ands[16][2] ),
    .A2(net835),
    .B1(net749),
    .B2(\tms1x00.O_pla_ands[17][2] ),
    .C1(net917),
    .X(_02396_));
 sky130_fd_sc_hd__o221a_1 _05905_ (.A1(\tms1x00.O_pla_ands[19][2] ),
    .A2(net858),
    .B1(net805),
    .B2(\tms1x00.O_pla_ands[20][2] ),
    .C1(_02396_),
    .X(_02397_));
 sky130_fd_sc_hd__a21o_2 _05906_ (.A1(_02395_),
    .A2(_02397_),
    .B1(_02393_),
    .X(_02398_));
 sky130_fd_sc_hd__o22a_1 _05907_ (.A1(_02383_),
    .A2(_02388_),
    .B1(_02398_),
    .B2(net926),
    .X(_02399_));
 sky130_fd_sc_hd__o22a_2 _05908_ (.A1(\tms1x00.ins_pla_ors[11][2] ),
    .A2(net852),
    .B1(net719),
    .B2(\tms1x00.ins_pla_ors[10][2] ),
    .X(_02400_));
 sky130_fd_sc_hd__o22a_1 _05909_ (.A1(\tms1x00.ins_pla_ors[12][2] ),
    .A2(net807),
    .B1(net757),
    .B2(\tms1x00.ins_pla_ors[9][2] ),
    .X(_02401_));
 sky130_fd_sc_hd__o221a_1 _05910_ (.A1(\tms1x00.ins_pla_ors[13][2] ),
    .A2(net889),
    .B1(net784),
    .B2(\tms1x00.ins_pla_ors[15][2] ),
    .C1(_02401_),
    .X(_02402_));
 sky130_fd_sc_hd__o211a_1 _05911_ (.A1(\tms1x00.ins_pla_ors[8][2] ),
    .A2(net838),
    .B1(_02402_),
    .C1(net996),
    .X(_02403_));
 sky130_fd_sc_hd__o211a_1 _05912_ (.A1(\tms1x00.ins_pla_ors[14][2] ),
    .A2(net617),
    .B1(_02400_),
    .C1(_02403_),
    .X(_02404_));
 sky130_fd_sc_hd__o22a_1 _05913_ (.A1(\tms1x00.ins_pla_ors[0][2] ),
    .A2(net841),
    .B1(net787),
    .B2(\tms1x00.ins_pla_ors[7][2] ),
    .X(_02405_));
 sky130_fd_sc_hd__o22a_1 _05914_ (.A1(\tms1x00.ins_pla_ors[3][2] ),
    .A2(net867),
    .B1(net760),
    .B2(\tms1x00.ins_pla_ors[1][2] ),
    .X(_02406_));
 sky130_fd_sc_hd__o221a_1 _05915_ (.A1(\tms1x00.ins_pla_ors[6][2] ),
    .A2(net619),
    .B1(net730),
    .B2(\tms1x00.ins_pla_ors[2][2] ),
    .C1(_02406_),
    .X(_02407_));
 sky130_fd_sc_hd__o211a_1 _05916_ (.A1(\tms1x00.ins_pla_ors[4][2] ),
    .A2(net811),
    .B1(_02407_),
    .C1(net919),
    .X(_02408_));
 sky130_fd_sc_hd__o211a_2 _05917_ (.A1(\tms1x00.ins_pla_ors[5][2] ),
    .A2(net892),
    .B1(_02405_),
    .C1(_02408_),
    .X(_02409_));
 sky130_fd_sc_hd__o21a_2 _05918_ (.A1(_02404_),
    .A2(_02409_),
    .B1(net600),
    .X(_02410_));
 sky130_fd_sc_hd__o221a_1 _05919_ (.A1(\tms1x00.O_pla_ors[0][2] ),
    .A2(net842),
    .B1(net762),
    .B2(\tms1x00.O_pla_ors[1][2] ),
    .C1(net599),
    .X(_02411_));
 sky130_fd_sc_hd__o22a_1 _05920_ (.A1(\tms1x00.O_pla_ors[6][2] ),
    .A2(net623),
    .B1(net789),
    .B2(\tms1x00.O_pla_ors[7][2] ),
    .X(_02412_));
 sky130_fd_sc_hd__o22a_1 _05921_ (.A1(\tms1x00.O_pla_ors[5][2] ),
    .A2(net898),
    .B1(net734),
    .B2(\tms1x00.O_pla_ors[2][2] ),
    .X(_02413_));
 sky130_fd_sc_hd__and3_1 _05922_ (.A(_02411_),
    .B(_02412_),
    .C(_02413_),
    .X(_02414_));
 sky130_fd_sc_hd__o221a_2 _05923_ (.A1(\tms1x00.O_pla_ors[3][2] ),
    .A2(net869),
    .B1(net814),
    .B2(\tms1x00.O_pla_ors[4][2] ),
    .C1(_02414_),
    .X(_02415_));
 sky130_fd_sc_hd__o22a_1 _05924_ (.A1(\tms1x00.ins_pla_ands[22][2] ),
    .A2(net606),
    .B1(net772),
    .B2(\tms1x00.ins_pla_ands[23][2] ),
    .X(_02416_));
 sky130_fd_sc_hd__o221a_1 _05925_ (.A1(\tms1x00.ins_pla_ands[21][2] ),
    .A2(net877),
    .B1(net797),
    .B2(\tms1x00.ins_pla_ands[20][2] ),
    .C1(net911),
    .X(_02417_));
 sky130_fd_sc_hd__o22a_1 _05926_ (.A1(\tms1x00.ins_pla_ands[19][2] ),
    .A2(net851),
    .B1(net715),
    .B2(\tms1x00.ins_pla_ands[18][2] ),
    .X(_02418_));
 sky130_fd_sc_hd__o211a_1 _05927_ (.A1(\tms1x00.ins_pla_ands[16][2] ),
    .A2(net826),
    .B1(_02417_),
    .C1(_02418_),
    .X(_02419_));
 sky130_fd_sc_hd__o211a_1 _05928_ (.A1(\tms1x00.ins_pla_ands[17][2] ),
    .A2(net746),
    .B1(_02416_),
    .C1(_02419_),
    .X(_02420_));
 sky130_fd_sc_hd__o22a_1 _05929_ (.A1(\tms1x00.ins_pla_ands[29][2] ),
    .A2(net879),
    .B1(net772),
    .B2(\tms1x00.ins_pla_ands[31][2] ),
    .X(_02421_));
 sky130_fd_sc_hd__o22a_1 _05930_ (.A1(\tms1x00.ins_pla_ands[24][2] ),
    .A2(net823),
    .B1(net796),
    .B2(\tms1x00.ins_pla_ands[28][2] ),
    .X(_02422_));
 sky130_fd_sc_hd__o221a_1 _05931_ (.A1(\tms1x00.ins_pla_ands[25][2] ),
    .A2(net743),
    .B1(net714),
    .B2(\tms1x00.ins_pla_ands[26][2] ),
    .C1(_02422_),
    .X(_02423_));
 sky130_fd_sc_hd__o211a_1 _05932_ (.A1(\tms1x00.ins_pla_ands[27][2] ),
    .A2(net850),
    .B1(_02423_),
    .C1(net990),
    .X(_02424_));
 sky130_fd_sc_hd__o211a_1 _05933_ (.A1(\tms1x00.ins_pla_ands[30][2] ),
    .A2(net605),
    .B1(_02421_),
    .C1(_02424_),
    .X(_02425_));
 sky130_fd_sc_hd__or3_2 _05934_ (.A(net924),
    .B(_02420_),
    .C(_02425_),
    .X(_02426_));
 sky130_fd_sc_hd__o22a_1 _05935_ (.A1(\tms1x00.ins_pla_ands[6][2] ),
    .A2(net613),
    .B1(net750),
    .B2(\tms1x00.ins_pla_ands[1][2] ),
    .X(_02427_));
 sky130_fd_sc_hd__o22a_1 _05936_ (.A1(\tms1x00.ins_pla_ands[5][2] ),
    .A2(net894),
    .B1(net870),
    .B2(\tms1x00.ins_pla_ands[3][2] ),
    .X(_02428_));
 sky130_fd_sc_hd__o221a_2 _05937_ (.A1(\tms1x00.ins_pla_ands[4][2] ),
    .A2(net812),
    .B1(net732),
    .B2(\tms1x00.ins_pla_ands[2][2] ),
    .C1(_02428_),
    .X(_02429_));
 sky130_fd_sc_hd__o211a_1 _05938_ (.A1(\tms1x00.ins_pla_ands[7][2] ),
    .A2(net779),
    .B1(_02429_),
    .C1(net916),
    .X(_02430_));
 sky130_fd_sc_hd__o211a_1 _05939_ (.A1(\tms1x00.ins_pla_ands[0][2] ),
    .A2(net832),
    .B1(_02427_),
    .C1(_02430_),
    .X(_02431_));
 sky130_fd_sc_hd__o22a_1 _05940_ (.A1(\tms1x00.ins_pla_ands[14][2] ),
    .A2(net609),
    .B1(net774),
    .B2(\tms1x00.ins_pla_ands[15][2] ),
    .X(_02432_));
 sky130_fd_sc_hd__o221a_1 _05941_ (.A1(\tms1x00.ins_pla_ands[13][2] ),
    .A2(net883),
    .B1(net801),
    .B2(\tms1x00.ins_pla_ands[12][2] ),
    .C1(net993),
    .X(_02433_));
 sky130_fd_sc_hd__o22a_1 _05942_ (.A1(\tms1x00.ins_pla_ands[11][2] ),
    .A2(net855),
    .B1(net721),
    .B2(\tms1x00.ins_pla_ands[10][2] ),
    .X(_02434_));
 sky130_fd_sc_hd__o211a_1 _05943_ (.A1(\tms1x00.ins_pla_ands[8][2] ),
    .A2(net829),
    .B1(_02433_),
    .C1(_02434_),
    .X(_02435_));
 sky130_fd_sc_hd__o211a_1 _05944_ (.A1(\tms1x00.ins_pla_ands[9][2] ),
    .A2(net751),
    .B1(_02432_),
    .C1(_02435_),
    .X(_02436_));
 sky130_fd_sc_hd__a211o_4 _05945_ (.A1(_01636_),
    .A2(_02399_),
    .B1(_02410_),
    .C1(_02415_),
    .X(_02437_));
 sky130_fd_sc_hd__o311a_1 _05946_ (.A1(net986),
    .A2(_02431_),
    .A3(_02436_),
    .B1(net712),
    .C1(_02426_),
    .X(_02438_));
 sky130_fd_sc_hd__a211o_1 _05947_ (.A1(net711),
    .A2(_02437_),
    .B1(_02438_),
    .C1(net586),
    .X(_02439_));
 sky130_fd_sc_hd__o211a_1 _05948_ (.A1(net589),
    .A2(_02378_),
    .B1(_02439_),
    .C1(net629),
    .X(_02440_));
 sky130_fd_sc_hd__a22o_1 _05949_ (.A1(net122),
    .A2(net579),
    .B1(_02378_),
    .B2(net583),
    .X(_02441_));
 sky130_fd_sc_hd__or2_1 _05950_ (.A(_02440_),
    .B(_02441_),
    .X(_00027_));
 sky130_fd_sc_hd__nand2_1 _05951_ (.A(net906),
    .B(\wbs_o_buff[3] ),
    .Y(_02442_));
 sky130_fd_sc_hd__o22a_1 _05952_ (.A1(\tms1x00.O_pla_ands[6][3] ),
    .A2(net622),
    .B1(net789),
    .B2(\tms1x00.O_pla_ands[7][3] ),
    .X(_02443_));
 sky130_fd_sc_hd__o221a_1 _05953_ (.A1(\tms1x00.O_pla_ands[0][3] ),
    .A2(net836),
    .B1(net753),
    .B2(\tms1x00.O_pla_ands[1][3] ),
    .C1(net914),
    .X(_02444_));
 sky130_fd_sc_hd__o22a_1 _05954_ (.A1(\tms1x00.O_pla_ands[3][3] ),
    .A2(net868),
    .B1(net733),
    .B2(\tms1x00.O_pla_ands[2][3] ),
    .X(_02445_));
 sky130_fd_sc_hd__o211a_1 _05955_ (.A1(\tms1x00.O_pla_ands[4][3] ),
    .A2(net814),
    .B1(_02444_),
    .C1(_02445_),
    .X(_02446_));
 sky130_fd_sc_hd__o211a_1 _05956_ (.A1(\tms1x00.O_pla_ands[5][3] ),
    .A2(net897),
    .B1(_02443_),
    .C1(_02446_),
    .X(_02447_));
 sky130_fd_sc_hd__o22a_1 _05957_ (.A1(\tms1x00.O_pla_ands[13][3] ),
    .A2(net899),
    .B1(net791),
    .B2(\tms1x00.O_pla_ands[15][3] ),
    .X(_02448_));
 sky130_fd_sc_hd__o22a_1 _05958_ (.A1(\tms1x00.O_pla_ands[8][3] ),
    .A2(net842),
    .B1(net762),
    .B2(\tms1x00.O_pla_ands[9][3] ),
    .X(_02449_));
 sky130_fd_sc_hd__o221a_1 _05959_ (.A1(\tms1x00.O_pla_ands[14][3] ),
    .A2(net624),
    .B1(net735),
    .B2(\tms1x00.O_pla_ands[10][3] ),
    .C1(_02449_),
    .X(_02450_));
 sky130_fd_sc_hd__o211a_1 _05960_ (.A1(\tms1x00.O_pla_ands[11][3] ),
    .A2(net871),
    .B1(_02450_),
    .C1(net999),
    .X(_02451_));
 sky130_fd_sc_hd__o211a_2 _05961_ (.A1(\tms1x00.O_pla_ands[12][3] ),
    .A2(net817),
    .B1(_02448_),
    .C1(_02451_),
    .X(_02452_));
 sky130_fd_sc_hd__or3_4 _05962_ (.A(net988),
    .B(_02447_),
    .C(_02452_),
    .X(_02453_));
 sky130_fd_sc_hd__o22a_1 _05963_ (.A1(\tms1x00.O_pla_ands[30][3] ),
    .A2(net611),
    .B1(net777),
    .B2(\tms1x00.O_pla_ands[31][3] ),
    .X(_02454_));
 sky130_fd_sc_hd__o221a_1 _05964_ (.A1(\tms1x00.O_pla_ands[29][3] ),
    .A2(net884),
    .B1(net803),
    .B2(\tms1x00.O_pla_ands[28][3] ),
    .C1(net992),
    .X(_02455_));
 sky130_fd_sc_hd__o22a_1 _05965_ (.A1(\tms1x00.O_pla_ands[27][3] ),
    .A2(net855),
    .B1(net722),
    .B2(\tms1x00.O_pla_ands[26][3] ),
    .X(_02456_));
 sky130_fd_sc_hd__o211a_1 _05966_ (.A1(\tms1x00.O_pla_ands[24][3] ),
    .A2(net830),
    .B1(_02455_),
    .C1(_02456_),
    .X(_02457_));
 sky130_fd_sc_hd__o211a_4 _05967_ (.A1(\tms1x00.O_pla_ands[25][3] ),
    .A2(net748),
    .B1(_02454_),
    .C1(_02457_),
    .X(_02458_));
 sky130_fd_sc_hd__o22a_2 _05968_ (.A1(\tms1x00.O_pla_ands[22][3] ),
    .A2(net610),
    .B1(net775),
    .B2(\tms1x00.O_pla_ands[23][3] ),
    .X(_02459_));
 sky130_fd_sc_hd__o221a_1 _05969_ (.A1(\tms1x00.O_pla_ands[16][3] ),
    .A2(net834),
    .B1(net752),
    .B2(\tms1x00.O_pla_ands[17][3] ),
    .C1(net915),
    .X(_02460_));
 sky130_fd_sc_hd__o22a_1 _05970_ (.A1(\tms1x00.O_pla_ands[19][3] ),
    .A2(net860),
    .B1(net724),
    .B2(\tms1x00.O_pla_ands[18][3] ),
    .X(_02461_));
 sky130_fd_sc_hd__o211a_1 _05971_ (.A1(\tms1x00.O_pla_ands[21][3] ),
    .A2(net885),
    .B1(_02460_),
    .C1(_02461_),
    .X(_02462_));
 sky130_fd_sc_hd__o211a_1 _05972_ (.A1(\tms1x00.O_pla_ands[20][3] ),
    .A2(net805),
    .B1(_02459_),
    .C1(_02462_),
    .X(_02463_));
 sky130_fd_sc_hd__o311a_4 _05973_ (.A1(net926),
    .A2(_02458_),
    .A3(_02463_),
    .B1(net905),
    .C1(_02453_),
    .X(_02464_));
 sky130_fd_sc_hd__or2_1 _05974_ (.A(\tms1x00.ins_pla_ors[1][3] ),
    .B(net759),
    .X(_02465_));
 sky130_fd_sc_hd__or2_1 _05975_ (.A(\tms1x00.ins_pla_ors[0][3] ),
    .B(net840),
    .X(_02466_));
 sky130_fd_sc_hd__o221a_1 _05976_ (.A1(\tms1x00.ins_pla_ors[5][3] ),
    .A2(net890),
    .B1(net807),
    .B2(\tms1x00.ins_pla_ors[4][3] ),
    .C1(net920),
    .X(_02467_));
 sky130_fd_sc_hd__o221a_1 _05977_ (.A1(\tms1x00.ins_pla_ors[6][3] ),
    .A2(net619),
    .B1(net786),
    .B2(\tms1x00.ins_pla_ors[7][3] ),
    .C1(_02465_),
    .X(_02468_));
 sky130_fd_sc_hd__o221a_1 _05978_ (.A1(\tms1x00.ins_pla_ors[3][3] ),
    .A2(net866),
    .B1(net730),
    .B2(\tms1x00.ins_pla_ors[2][3] ),
    .C1(_02466_),
    .X(_02469_));
 sky130_fd_sc_hd__o22a_1 _05979_ (.A1(\tms1x00.ins_pla_ors[11][3] ),
    .A2(net862),
    .B1(net727),
    .B2(\tms1x00.ins_pla_ors[10][3] ),
    .X(_02470_));
 sky130_fd_sc_hd__o22a_1 _05980_ (.A1(\tms1x00.ins_pla_ors[14][3] ),
    .A2(net605),
    .B1(net783),
    .B2(\tms1x00.ins_pla_ors[15][3] ),
    .X(_02471_));
 sky130_fd_sc_hd__o221a_1 _05981_ (.A1(\tms1x00.ins_pla_ors[8][3] ),
    .A2(net837),
    .B1(net745),
    .B2(\tms1x00.ins_pla_ors[9][3] ),
    .C1(net997),
    .X(_02472_));
 sky130_fd_sc_hd__o211a_1 _05982_ (.A1(\tms1x00.ins_pla_ors[12][3] ),
    .A2(net806),
    .B1(_02471_),
    .C1(_02472_),
    .X(_02473_));
 sky130_fd_sc_hd__o211a_2 _05983_ (.A1(\tms1x00.ins_pla_ors[13][3] ),
    .A2(net888),
    .B1(_02470_),
    .C1(_02473_),
    .X(_02474_));
 sky130_fd_sc_hd__a31o_2 _05984_ (.A1(_02467_),
    .A2(_02468_),
    .A3(_02469_),
    .B1(_02474_),
    .X(_02475_));
 sky130_fd_sc_hd__o221a_1 _05985_ (.A1(\tms1x00.O_pla_ors[0][3] ),
    .A2(net842),
    .B1(net762),
    .B2(\tms1x00.O_pla_ors[1][3] ),
    .C1(net599),
    .X(_02476_));
 sky130_fd_sc_hd__o22a_1 _05986_ (.A1(\tms1x00.O_pla_ors[6][3] ),
    .A2(net626),
    .B1(net789),
    .B2(\tms1x00.O_pla_ors[7][3] ),
    .X(_02477_));
 sky130_fd_sc_hd__o22a_1 _05987_ (.A1(\tms1x00.O_pla_ors[5][3] ),
    .A2(net900),
    .B1(net737),
    .B2(\tms1x00.O_pla_ors[2][3] ),
    .X(_02478_));
 sky130_fd_sc_hd__and3_1 _05988_ (.A(_02476_),
    .B(_02477_),
    .C(_02478_),
    .X(_02479_));
 sky130_fd_sc_hd__o221a_2 _05989_ (.A1(\tms1x00.O_pla_ors[3][3] ),
    .A2(net872),
    .B1(net818),
    .B2(\tms1x00.O_pla_ors[4][3] ),
    .C1(_02479_),
    .X(_02480_));
 sky130_fd_sc_hd__o22a_1 _05990_ (.A1(\tms1x00.ins_pla_ands[22][3] ),
    .A2(net606),
    .B1(net772),
    .B2(\tms1x00.ins_pla_ands[23][3] ),
    .X(_02481_));
 sky130_fd_sc_hd__o221a_1 _05991_ (.A1(\tms1x00.ins_pla_ands[21][3] ),
    .A2(net878),
    .B1(net797),
    .B2(\tms1x00.ins_pla_ands[20][3] ),
    .C1(net911),
    .X(_02482_));
 sky130_fd_sc_hd__o22a_1 _05992_ (.A1(\tms1x00.ins_pla_ands[19][3] ),
    .A2(net851),
    .B1(net715),
    .B2(\tms1x00.ins_pla_ands[18][3] ),
    .X(_02483_));
 sky130_fd_sc_hd__o211a_1 _05993_ (.A1(\tms1x00.ins_pla_ands[16][3] ),
    .A2(net826),
    .B1(_02482_),
    .C1(_02483_),
    .X(_02484_));
 sky130_fd_sc_hd__o211a_1 _05994_ (.A1(\tms1x00.ins_pla_ands[17][3] ),
    .A2(net746),
    .B1(_02481_),
    .C1(_02484_),
    .X(_02485_));
 sky130_fd_sc_hd__o22a_1 _05995_ (.A1(\tms1x00.ins_pla_ands[27][3] ),
    .A2(net850),
    .B1(net714),
    .B2(\tms1x00.ins_pla_ands[26][3] ),
    .X(_02486_));
 sky130_fd_sc_hd__o221a_1 _05996_ (.A1(\tms1x00.ins_pla_ands[29][3] ),
    .A2(net877),
    .B1(net796),
    .B2(\tms1x00.ins_pla_ands[28][3] ),
    .C1(net991),
    .X(_02487_));
 sky130_fd_sc_hd__o22a_1 _05997_ (.A1(\tms1x00.ins_pla_ands[30][3] ),
    .A2(net602),
    .B1(net769),
    .B2(\tms1x00.ins_pla_ands[31][3] ),
    .X(_02488_));
 sky130_fd_sc_hd__o211a_1 _05998_ (.A1(\tms1x00.ins_pla_ands[25][3] ),
    .A2(net742),
    .B1(_02487_),
    .C1(_02488_),
    .X(_02489_));
 sky130_fd_sc_hd__o211a_2 _05999_ (.A1(\tms1x00.ins_pla_ands[24][3] ),
    .A2(net823),
    .B1(_02486_),
    .C1(_02489_),
    .X(_02490_));
 sky130_fd_sc_hd__or3_2 _06000_ (.A(net924),
    .B(_02485_),
    .C(_02490_),
    .X(_02491_));
 sky130_fd_sc_hd__o22a_1 _06001_ (.A1(\tms1x00.ins_pla_ands[14][3] ),
    .A2(net609),
    .B1(net779),
    .B2(\tms1x00.ins_pla_ands[15][3] ),
    .X(_02492_));
 sky130_fd_sc_hd__o221a_1 _06002_ (.A1(\tms1x00.ins_pla_ands[13][3] ),
    .A2(net882),
    .B1(net801),
    .B2(\tms1x00.ins_pla_ands[12][3] ),
    .C1(net993),
    .X(_02493_));
 sky130_fd_sc_hd__o22a_1 _06003_ (.A1(\tms1x00.ins_pla_ands[11][3] ),
    .A2(net855),
    .B1(net720),
    .B2(\tms1x00.ins_pla_ands[10][3] ),
    .X(_02494_));
 sky130_fd_sc_hd__o211a_1 _06004_ (.A1(\tms1x00.ins_pla_ands[8][3] ),
    .A2(net829),
    .B1(_02493_),
    .C1(_02494_),
    .X(_02495_));
 sky130_fd_sc_hd__o211a_1 _06005_ (.A1(\tms1x00.ins_pla_ands[9][3] ),
    .A2(net751),
    .B1(_02492_),
    .C1(_02495_),
    .X(_02496_));
 sky130_fd_sc_hd__o22a_1 _06006_ (.A1(\tms1x00.ins_pla_ands[5][3] ),
    .A2(net894),
    .B1(net732),
    .B2(\tms1x00.ins_pla_ands[2][3] ),
    .X(_02497_));
 sky130_fd_sc_hd__o22a_1 _06007_ (.A1(\tms1x00.ins_pla_ands[0][3] ),
    .A2(net832),
    .B1(net779),
    .B2(\tms1x00.ins_pla_ands[7][3] ),
    .X(_02498_));
 sky130_fd_sc_hd__o221a_1 _06008_ (.A1(\tms1x00.ins_pla_ands[6][3] ),
    .A2(net613),
    .B1(net859),
    .B2(\tms1x00.ins_pla_ands[3][3] ),
    .C1(_02498_),
    .X(_02499_));
 sky130_fd_sc_hd__o211a_1 _06009_ (.A1(\tms1x00.ins_pla_ands[4][3] ),
    .A2(net812),
    .B1(_02499_),
    .C1(net916),
    .X(_02500_));
 sky130_fd_sc_hd__o211a_1 _06010_ (.A1(\tms1x00.ins_pla_ands[1][3] ),
    .A2(net750),
    .B1(_02497_),
    .C1(_02500_),
    .X(_02501_));
 sky130_fd_sc_hd__a211o_2 _06011_ (.A1(net600),
    .A2(_02475_),
    .B1(_02480_),
    .C1(_02464_),
    .X(_02502_));
 sky130_fd_sc_hd__o311a_1 _06012_ (.A1(net986),
    .A2(_02496_),
    .A3(_02501_),
    .B1(net712),
    .C1(_02491_),
    .X(_02503_));
 sky130_fd_sc_hd__a211o_1 _06013_ (.A1(_02281_),
    .A2(_02502_),
    .B1(_02503_),
    .C1(net586),
    .X(_02504_));
 sky130_fd_sc_hd__a21oi_1 _06014_ (.A1(net586),
    .A2(_02442_),
    .B1(_02223_),
    .Y(_02505_));
 sky130_fd_sc_hd__a22o_1 _06015_ (.A1(net123),
    .A2(net579),
    .B1(_02504_),
    .B2(_02505_),
    .X(_02506_));
 sky130_fd_sc_hd__a31o_1 _06016_ (.A1(net906),
    .A2(\wbs_o_buff[3] ),
    .A3(net583),
    .B1(_02506_),
    .X(_00030_));
 sky130_fd_sc_hd__nand2_1 _06017_ (.A(net906),
    .B(\wbs_o_buff[4] ),
    .Y(_02507_));
 sky130_fd_sc_hd__o22a_1 _06018_ (.A1(\tms1x00.O_pla_ands[6][4] ),
    .A2(net622),
    .B1(net788),
    .B2(\tms1x00.O_pla_ands[7][4] ),
    .X(_02508_));
 sky130_fd_sc_hd__o221a_2 _06019_ (.A1(\tms1x00.O_pla_ands[0][4] ),
    .A2(net834),
    .B1(net752),
    .B2(\tms1x00.O_pla_ands[1][4] ),
    .C1(net915),
    .X(_02509_));
 sky130_fd_sc_hd__o22a_1 _06020_ (.A1(\tms1x00.O_pla_ands[3][4] ),
    .A2(net869),
    .B1(net733),
    .B2(\tms1x00.O_pla_ands[2][4] ),
    .X(_02510_));
 sky130_fd_sc_hd__o211a_1 _06021_ (.A1(\tms1x00.O_pla_ands[5][4] ),
    .A2(net897),
    .B1(_02509_),
    .C1(_02510_),
    .X(_02511_));
 sky130_fd_sc_hd__o211a_1 _06022_ (.A1(\tms1x00.O_pla_ands[4][4] ),
    .A2(net814),
    .B1(_02508_),
    .C1(_02511_),
    .X(_02512_));
 sky130_fd_sc_hd__or2_1 _06023_ (.A(\tms1x00.O_pla_ands[9][4] ),
    .B(net765),
    .X(_02513_));
 sky130_fd_sc_hd__o221a_1 _06024_ (.A1(\tms1x00.O_pla_ands[14][4] ),
    .A2(net623),
    .B1(net897),
    .B2(\tms1x00.O_pla_ands[13][4] ),
    .C1(_02513_),
    .X(_02514_));
 sky130_fd_sc_hd__o22a_1 _06025_ (.A1(\tms1x00.O_pla_ands[8][4] ),
    .A2(net843),
    .B1(net790),
    .B2(\tms1x00.O_pla_ands[15][4] ),
    .X(_02515_));
 sky130_fd_sc_hd__o221a_2 _06026_ (.A1(\tms1x00.O_pla_ands[12][4] ),
    .A2(net817),
    .B1(net735),
    .B2(\tms1x00.O_pla_ands[10][4] ),
    .C1(_02515_),
    .X(_02516_));
 sky130_fd_sc_hd__o211a_1 _06027_ (.A1(\tms1x00.O_pla_ands[11][4] ),
    .A2(net869),
    .B1(_02516_),
    .C1(net999),
    .X(_02517_));
 sky130_fd_sc_hd__a211o_2 _06028_ (.A1(_02514_),
    .A2(_02517_),
    .B1(net988),
    .C1(_02512_),
    .X(_02518_));
 sky130_fd_sc_hd__o22a_1 _06029_ (.A1(\tms1x00.O_pla_ands[30][4] ),
    .A2(net611),
    .B1(net777),
    .B2(\tms1x00.O_pla_ands[31][4] ),
    .X(_02519_));
 sky130_fd_sc_hd__o22a_1 _06030_ (.A1(\tms1x00.O_pla_ands[27][4] ),
    .A2(net855),
    .B1(net722),
    .B2(\tms1x00.O_pla_ands[26][4] ),
    .X(_02520_));
 sky130_fd_sc_hd__o221a_1 _06031_ (.A1(\tms1x00.O_pla_ands[29][4] ),
    .A2(net884),
    .B1(net803),
    .B2(\tms1x00.O_pla_ands[28][4] ),
    .C1(net992),
    .X(_02521_));
 sky130_fd_sc_hd__o211a_1 _06032_ (.A1(\tms1x00.O_pla_ands[24][4] ),
    .A2(net830),
    .B1(_02520_),
    .C1(_02521_),
    .X(_02522_));
 sky130_fd_sc_hd__o211a_4 _06033_ (.A1(\tms1x00.O_pla_ands[25][4] ),
    .A2(net748),
    .B1(_02519_),
    .C1(_02522_),
    .X(_02523_));
 sky130_fd_sc_hd__o22a_1 _06034_ (.A1(\tms1x00.O_pla_ands[22][4] ),
    .A2(net610),
    .B1(net775),
    .B2(\tms1x00.O_pla_ands[23][4] ),
    .X(_02524_));
 sky130_fd_sc_hd__o221a_1 _06035_ (.A1(\tms1x00.O_pla_ands[16][4] ),
    .A2(net835),
    .B1(net753),
    .B2(\tms1x00.O_pla_ands[17][4] ),
    .C1(net914),
    .X(_02525_));
 sky130_fd_sc_hd__o22a_1 _06036_ (.A1(\tms1x00.O_pla_ands[19][4] ),
    .A2(net858),
    .B1(net724),
    .B2(\tms1x00.O_pla_ands[18][4] ),
    .X(_02526_));
 sky130_fd_sc_hd__o211a_1 _06037_ (.A1(\tms1x00.O_pla_ands[21][4] ),
    .A2(net886),
    .B1(_02525_),
    .C1(_02526_),
    .X(_02527_));
 sky130_fd_sc_hd__o211a_1 _06038_ (.A1(\tms1x00.O_pla_ands[20][4] ),
    .A2(net805),
    .B1(_02524_),
    .C1(_02527_),
    .X(_02528_));
 sky130_fd_sc_hd__o311a_2 _06039_ (.A1(net925),
    .A2(_02523_),
    .A3(_02528_),
    .B1(net905),
    .C1(_02518_),
    .X(_02529_));
 sky130_fd_sc_hd__o22a_1 _06040_ (.A1(\tms1x00.ins_pla_ors[11][4] ),
    .A2(net863),
    .B1(net807),
    .B2(\tms1x00.ins_pla_ors[12][4] ),
    .X(_02530_));
 sky130_fd_sc_hd__o22a_1 _06041_ (.A1(\tms1x00.ins_pla_ors[13][4] ),
    .A2(net881),
    .B1(net717),
    .B2(\tms1x00.ins_pla_ors[10][4] ),
    .X(_02531_));
 sky130_fd_sc_hd__o221a_2 _06042_ (.A1(\tms1x00.ins_pla_ors[14][4] ),
    .A2(net606),
    .B1(net773),
    .B2(\tms1x00.ins_pla_ors[15][4] ),
    .C1(_02531_),
    .X(_02532_));
 sky130_fd_sc_hd__o221a_1 _06043_ (.A1(\tms1x00.ins_pla_ors[8][4] ),
    .A2(net838),
    .B1(net757),
    .B2(\tms1x00.ins_pla_ors[9][4] ),
    .C1(net996),
    .X(_02533_));
 sky130_fd_sc_hd__o22a_1 _06044_ (.A1(\tms1x00.ins_pla_ors[0][4] ),
    .A2(net840),
    .B1(net759),
    .B2(\tms1x00.ins_pla_ors[1][4] ),
    .X(_02534_));
 sky130_fd_sc_hd__o22a_1 _06045_ (.A1(\tms1x00.ins_pla_ors[3][4] ),
    .A2(net866),
    .B1(net786),
    .B2(\tms1x00.ins_pla_ors[7][4] ),
    .X(_02535_));
 sky130_fd_sc_hd__o221a_2 _06046_ (.A1(\tms1x00.ins_pla_ors[6][4] ),
    .A2(net620),
    .B1(net730),
    .B2(\tms1x00.ins_pla_ors[2][4] ),
    .C1(_02535_),
    .X(_02536_));
 sky130_fd_sc_hd__o211a_1 _06047_ (.A1(\tms1x00.ins_pla_ors[4][4] ),
    .A2(net810),
    .B1(_02536_),
    .C1(net920),
    .X(_02537_));
 sky130_fd_sc_hd__o211a_2 _06048_ (.A1(\tms1x00.ins_pla_ors[5][4] ),
    .A2(net892),
    .B1(_02534_),
    .C1(_02537_),
    .X(_02538_));
 sky130_fd_sc_hd__a31o_2 _06049_ (.A1(_02530_),
    .A2(_02532_),
    .A3(_02533_),
    .B1(_02538_),
    .X(_02539_));
 sky130_fd_sc_hd__o22a_1 _06050_ (.A1(\tms1x00.O_pla_ors[0][4] ),
    .A2(net845),
    .B1(net732),
    .B2(\tms1x00.O_pla_ors[2][4] ),
    .X(_02540_));
 sky130_fd_sc_hd__o22a_1 _06051_ (.A1(\tms1x00.O_pla_ors[7][4] ),
    .A2(net788),
    .B1(net765),
    .B2(\tms1x00.O_pla_ors[1][4] ),
    .X(_02541_));
 sky130_fd_sc_hd__o221a_1 _06052_ (.A1(\tms1x00.O_pla_ors[6][4] ),
    .A2(net623),
    .B1(net869),
    .B2(\tms1x00.O_pla_ors[3][4] ),
    .C1(_02541_),
    .X(_02542_));
 sky130_fd_sc_hd__o211a_1 _06053_ (.A1(\tms1x00.O_pla_ors[4][4] ),
    .A2(net814),
    .B1(net599),
    .C1(_02542_),
    .X(_02543_));
 sky130_fd_sc_hd__o211a_2 _06054_ (.A1(\tms1x00.O_pla_ors[5][4] ),
    .A2(net895),
    .B1(_02540_),
    .C1(_02543_),
    .X(_02544_));
 sky130_fd_sc_hd__o22a_1 _06055_ (.A1(\tms1x00.ins_pla_ands[27][4] ),
    .A2(net850),
    .B1(net716),
    .B2(\tms1x00.ins_pla_ands[26][4] ),
    .X(_02545_));
 sky130_fd_sc_hd__o221a_1 _06056_ (.A1(\tms1x00.ins_pla_ands[30][4] ),
    .A2(net602),
    .B1(net743),
    .B2(\tms1x00.ins_pla_ands[25][4] ),
    .C1(_02545_),
    .X(_02546_));
 sky130_fd_sc_hd__o221a_2 _06057_ (.A1(\tms1x00.ins_pla_ands[29][4] ),
    .A2(net879),
    .B1(net798),
    .B2(\tms1x00.ins_pla_ands[28][4] ),
    .C1(net990),
    .X(_02547_));
 sky130_fd_sc_hd__o221a_1 _06058_ (.A1(\tms1x00.ins_pla_ands[24][4] ),
    .A2(net824),
    .B1(net769),
    .B2(\tms1x00.ins_pla_ands[31][4] ),
    .C1(_02547_),
    .X(_02548_));
 sky130_fd_sc_hd__and2_2 _06059_ (.A(_02546_),
    .B(_02548_),
    .X(_02549_));
 sky130_fd_sc_hd__o22a_1 _06060_ (.A1(\tms1x00.ins_pla_ands[22][4] ),
    .A2(net606),
    .B1(net773),
    .B2(\tms1x00.ins_pla_ands[23][4] ),
    .X(_02550_));
 sky130_fd_sc_hd__o221a_4 _06061_ (.A1(\tms1x00.ins_pla_ands[21][4] ),
    .A2(net877),
    .B1(net796),
    .B2(\tms1x00.ins_pla_ands[20][4] ),
    .C1(net911),
    .X(_02551_));
 sky130_fd_sc_hd__o22a_1 _06062_ (.A1(\tms1x00.ins_pla_ands[19][4] ),
    .A2(net853),
    .B1(net718),
    .B2(\tms1x00.ins_pla_ands[18][4] ),
    .X(_02552_));
 sky130_fd_sc_hd__o211a_1 _06063_ (.A1(\tms1x00.ins_pla_ands[16][4] ),
    .A2(net828),
    .B1(_02551_),
    .C1(_02552_),
    .X(_02553_));
 sky130_fd_sc_hd__o211a_1 _06064_ (.A1(\tms1x00.ins_pla_ands[17][4] ),
    .A2(net745),
    .B1(_02550_),
    .C1(_02553_),
    .X(_02554_));
 sky130_fd_sc_hd__o22a_1 _06065_ (.A1(\tms1x00.ins_pla_ands[6][4] ),
    .A2(net614),
    .B1(net751),
    .B2(\tms1x00.ins_pla_ands[1][4] ),
    .X(_02555_));
 sky130_fd_sc_hd__o22a_1 _06066_ (.A1(\tms1x00.ins_pla_ands[3][4] ),
    .A2(net870),
    .B1(net815),
    .B2(\tms1x00.ins_pla_ands[4][4] ),
    .X(_02556_));
 sky130_fd_sc_hd__o221a_2 _06067_ (.A1(\tms1x00.ins_pla_ands[5][4] ),
    .A2(net894),
    .B1(net732),
    .B2(\tms1x00.ins_pla_ands[2][4] ),
    .C1(_02556_),
    .X(_02557_));
 sky130_fd_sc_hd__o211a_1 _06068_ (.A1(\tms1x00.ins_pla_ands[7][4] ),
    .A2(net780),
    .B1(_02557_),
    .C1(net916),
    .X(_02558_));
 sky130_fd_sc_hd__o211a_1 _06069_ (.A1(\tms1x00.ins_pla_ands[0][4] ),
    .A2(net833),
    .B1(_02555_),
    .C1(_02558_),
    .X(_02559_));
 sky130_fd_sc_hd__o22a_1 _06070_ (.A1(\tms1x00.ins_pla_ands[14][4] ),
    .A2(net608),
    .B1(net778),
    .B2(\tms1x00.ins_pla_ands[15][4] ),
    .X(_02560_));
 sky130_fd_sc_hd__o221a_1 _06071_ (.A1(\tms1x00.ins_pla_ands[13][4] ),
    .A2(net882),
    .B1(net801),
    .B2(\tms1x00.ins_pla_ands[12][4] ),
    .C1(net993),
    .X(_02561_));
 sky130_fd_sc_hd__o22a_1 _06072_ (.A1(\tms1x00.ins_pla_ands[11][4] ),
    .A2(net854),
    .B1(net720),
    .B2(\tms1x00.ins_pla_ands[10][4] ),
    .X(_02562_));
 sky130_fd_sc_hd__o211a_1 _06073_ (.A1(\tms1x00.ins_pla_ands[8][4] ),
    .A2(net831),
    .B1(_02561_),
    .C1(_02562_),
    .X(_02563_));
 sky130_fd_sc_hd__o211a_1 _06074_ (.A1(\tms1x00.ins_pla_ands[9][4] ),
    .A2(net747),
    .B1(_02560_),
    .C1(_02563_),
    .X(_02564_));
 sky130_fd_sc_hd__or3_1 _06075_ (.A(net986),
    .B(_02559_),
    .C(_02564_),
    .X(_02565_));
 sky130_fd_sc_hd__a211o_2 _06076_ (.A1(net600),
    .A2(_02539_),
    .B1(_02544_),
    .C1(_02529_),
    .X(_02566_));
 sky130_fd_sc_hd__o31a_1 _06077_ (.A1(net924),
    .A2(_02549_),
    .A3(_02554_),
    .B1(net712),
    .X(_02567_));
 sky130_fd_sc_hd__a221o_1 _06078_ (.A1(net711),
    .A2(_02566_),
    .B1(_02567_),
    .B2(_02565_),
    .C1(net586),
    .X(_02568_));
 sky130_fd_sc_hd__a21oi_1 _06079_ (.A1(net586),
    .A2(_02507_),
    .B1(_02223_),
    .Y(_02569_));
 sky130_fd_sc_hd__a22o_1 _06080_ (.A1(net124),
    .A2(net579),
    .B1(_02568_),
    .B2(_02569_),
    .X(_02570_));
 sky130_fd_sc_hd__a31o_1 _06081_ (.A1(net906),
    .A2(\wbs_o_buff[4] ),
    .A3(net583),
    .B1(_02570_),
    .X(_00031_));
 sky130_fd_sc_hd__and2_1 _06082_ (.A(net907),
    .B(\wbs_o_buff[5] ),
    .X(_02571_));
 sky130_fd_sc_hd__o22a_1 _06083_ (.A1(\tms1x00.O_pla_ands[6][5] ),
    .A2(net622),
    .B1(net788),
    .B2(\tms1x00.O_pla_ands[7][5] ),
    .X(_02572_));
 sky130_fd_sc_hd__o221a_1 _06084_ (.A1(\tms1x00.O_pla_ands[0][5] ),
    .A2(net834),
    .B1(net752),
    .B2(\tms1x00.O_pla_ands[1][5] ),
    .C1(net914),
    .X(_02573_));
 sky130_fd_sc_hd__o22a_1 _06085_ (.A1(\tms1x00.O_pla_ands[3][5] ),
    .A2(net868),
    .B1(net733),
    .B2(\tms1x00.O_pla_ands[2][5] ),
    .X(_02574_));
 sky130_fd_sc_hd__o211a_1 _06086_ (.A1(\tms1x00.O_pla_ands[5][5] ),
    .A2(net897),
    .B1(_02573_),
    .C1(_02574_),
    .X(_02575_));
 sky130_fd_sc_hd__o211a_1 _06087_ (.A1(\tms1x00.O_pla_ands[4][5] ),
    .A2(net813),
    .B1(_02572_),
    .C1(_02575_),
    .X(_02576_));
 sky130_fd_sc_hd__o22a_1 _06088_ (.A1(\tms1x00.O_pla_ands[13][5] ),
    .A2(net898),
    .B1(net790),
    .B2(\tms1x00.O_pla_ands[15][5] ),
    .X(_02577_));
 sky130_fd_sc_hd__o22a_1 _06089_ (.A1(\tms1x00.O_pla_ands[8][5] ),
    .A2(net842),
    .B1(net762),
    .B2(\tms1x00.O_pla_ands[9][5] ),
    .X(_02578_));
 sky130_fd_sc_hd__o221a_1 _06090_ (.A1(\tms1x00.O_pla_ands[12][5] ),
    .A2(net816),
    .B1(net735),
    .B2(\tms1x00.O_pla_ands[10][5] ),
    .C1(_02578_),
    .X(_02579_));
 sky130_fd_sc_hd__o211a_1 _06091_ (.A1(\tms1x00.O_pla_ands[11][5] ),
    .A2(net871),
    .B1(_02579_),
    .C1(net999),
    .X(_02580_));
 sky130_fd_sc_hd__o211a_2 _06092_ (.A1(\tms1x00.O_pla_ands[14][5] ),
    .A2(net624),
    .B1(_02577_),
    .C1(_02580_),
    .X(_02581_));
 sky130_fd_sc_hd__or3_2 _06093_ (.A(net988),
    .B(_02576_),
    .C(_02581_),
    .X(_02582_));
 sky130_fd_sc_hd__o22a_1 _06094_ (.A1(\tms1x00.O_pla_ands[30][5] ),
    .A2(net611),
    .B1(net777),
    .B2(\tms1x00.O_pla_ands[31][5] ),
    .X(_02583_));
 sky130_fd_sc_hd__o22a_1 _06095_ (.A1(\tms1x00.O_pla_ands[27][5] ),
    .A2(net856),
    .B1(net722),
    .B2(\tms1x00.O_pla_ands[26][5] ),
    .X(_02584_));
 sky130_fd_sc_hd__o221a_1 _06096_ (.A1(\tms1x00.O_pla_ands[29][5] ),
    .A2(net884),
    .B1(net803),
    .B2(\tms1x00.O_pla_ands[28][5] ),
    .C1(net992),
    .X(_02585_));
 sky130_fd_sc_hd__o211a_1 _06097_ (.A1(\tms1x00.O_pla_ands[24][5] ),
    .A2(net830),
    .B1(_02584_),
    .C1(_02585_),
    .X(_02586_));
 sky130_fd_sc_hd__o211a_2 _06098_ (.A1(\tms1x00.O_pla_ands[25][5] ),
    .A2(net748),
    .B1(_02583_),
    .C1(_02586_),
    .X(_02587_));
 sky130_fd_sc_hd__o22a_1 _06099_ (.A1(\tms1x00.O_pla_ands[22][5] ),
    .A2(net610),
    .B1(net775),
    .B2(\tms1x00.O_pla_ands[23][5] ),
    .X(_02588_));
 sky130_fd_sc_hd__o221a_1 _06100_ (.A1(\tms1x00.O_pla_ands[16][5] ),
    .A2(net835),
    .B1(net753),
    .B2(\tms1x00.O_pla_ands[17][5] ),
    .C1(net914),
    .X(_02589_));
 sky130_fd_sc_hd__o22a_1 _06101_ (.A1(\tms1x00.O_pla_ands[19][5] ),
    .A2(net858),
    .B1(net724),
    .B2(\tms1x00.O_pla_ands[18][5] ),
    .X(_02590_));
 sky130_fd_sc_hd__o211a_1 _06102_ (.A1(\tms1x00.O_pla_ands[21][5] ),
    .A2(net885),
    .B1(_02589_),
    .C1(_02590_),
    .X(_02591_));
 sky130_fd_sc_hd__o211a_2 _06103_ (.A1(\tms1x00.O_pla_ands[20][5] ),
    .A2(net805),
    .B1(_02588_),
    .C1(_02591_),
    .X(_02592_));
 sky130_fd_sc_hd__o311a_2 _06104_ (.A1(net926),
    .A2(_02587_),
    .A3(_02592_),
    .B1(net905),
    .C1(_02582_),
    .X(_02593_));
 sky130_fd_sc_hd__o22a_1 _06105_ (.A1(\tms1x00.ins_pla_ors[11][5] ),
    .A2(net853),
    .B1(net719),
    .B2(\tms1x00.ins_pla_ors[10][5] ),
    .X(_02594_));
 sky130_fd_sc_hd__or2_1 _06106_ (.A(\tms1x00.ins_pla_ors[14][5] ),
    .B(net617),
    .X(_02595_));
 sky130_fd_sc_hd__o22a_1 _06107_ (.A1(\tms1x00.ins_pla_ors[13][5] ),
    .A2(net889),
    .B1(net757),
    .B2(\tms1x00.ins_pla_ors[9][5] ),
    .X(_02596_));
 sky130_fd_sc_hd__o221a_1 _06108_ (.A1(\tms1x00.ins_pla_ors[12][5] ),
    .A2(net807),
    .B1(net784),
    .B2(\tms1x00.ins_pla_ors[15][5] ),
    .C1(_02596_),
    .X(_02597_));
 sky130_fd_sc_hd__o211a_1 _06109_ (.A1(\tms1x00.ins_pla_ors[8][5] ),
    .A2(net838),
    .B1(_02597_),
    .C1(net996),
    .X(_02598_));
 sky130_fd_sc_hd__o22a_1 _06110_ (.A1(\tms1x00.ins_pla_ors[7][5] ),
    .A2(net786),
    .B1(net730),
    .B2(\tms1x00.ins_pla_ors[2][5] ),
    .X(_02599_));
 sky130_fd_sc_hd__o22a_1 _06111_ (.A1(\tms1x00.ins_pla_ors[3][5] ),
    .A2(net866),
    .B1(net759),
    .B2(\tms1x00.ins_pla_ors[1][5] ),
    .X(_02600_));
 sky130_fd_sc_hd__o221a_2 _06112_ (.A1(\tms1x00.ins_pla_ors[6][5] ),
    .A2(net619),
    .B1(net840),
    .B2(\tms1x00.ins_pla_ors[0][5] ),
    .C1(_02600_),
    .X(_02601_));
 sky130_fd_sc_hd__o211a_1 _06113_ (.A1(\tms1x00.ins_pla_ors[4][5] ),
    .A2(net810),
    .B1(_02601_),
    .C1(net919),
    .X(_02602_));
 sky130_fd_sc_hd__o211a_2 _06114_ (.A1(\tms1x00.ins_pla_ors[5][5] ),
    .A2(net892),
    .B1(_02599_),
    .C1(_02602_),
    .X(_02603_));
 sky130_fd_sc_hd__a31o_1 _06115_ (.A1(_02594_),
    .A2(_02595_),
    .A3(_02598_),
    .B1(_02603_),
    .X(_02604_));
 sky130_fd_sc_hd__o221a_1 _06116_ (.A1(\tms1x00.O_pla_ors[0][5] ),
    .A2(net843),
    .B1(net763),
    .B2(\tms1x00.O_pla_ors[1][5] ),
    .C1(net599),
    .X(_02605_));
 sky130_fd_sc_hd__o22a_1 _06117_ (.A1(\tms1x00.O_pla_ors[6][5] ),
    .A2(net625),
    .B1(net791),
    .B2(\tms1x00.O_pla_ors[7][5] ),
    .X(_02606_));
 sky130_fd_sc_hd__o22a_1 _06118_ (.A1(\tms1x00.O_pla_ors[5][5] ),
    .A2(net899),
    .B1(net736),
    .B2(\tms1x00.O_pla_ors[2][5] ),
    .X(_02607_));
 sky130_fd_sc_hd__and3_2 _06119_ (.A(_02605_),
    .B(_02606_),
    .C(_02607_),
    .X(_02608_));
 sky130_fd_sc_hd__o221a_4 _06120_ (.A1(\tms1x00.O_pla_ors[3][5] ),
    .A2(net872),
    .B1(net817),
    .B2(\tms1x00.O_pla_ors[4][5] ),
    .C1(_02608_),
    .X(_02609_));
 sky130_fd_sc_hd__o22a_1 _06121_ (.A1(\tms1x00.ins_pla_ands[16][5] ),
    .A2(net827),
    .B1(net773),
    .B2(\tms1x00.ins_pla_ands[23][5] ),
    .X(_02610_));
 sky130_fd_sc_hd__o221a_2 _06122_ (.A1(\tms1x00.ins_pla_ands[21][5] ),
    .A2(net877),
    .B1(net796),
    .B2(\tms1x00.ins_pla_ands[20][5] ),
    .C1(net911),
    .X(_02611_));
 sky130_fd_sc_hd__o22a_1 _06123_ (.A1(\tms1x00.ins_pla_ands[19][5] ),
    .A2(net853),
    .B1(net718),
    .B2(\tms1x00.ins_pla_ands[18][5] ),
    .X(_02612_));
 sky130_fd_sc_hd__o221a_1 _06124_ (.A1(\tms1x00.ins_pla_ands[22][5] ),
    .A2(net606),
    .B1(net745),
    .B2(\tms1x00.ins_pla_ands[17][5] ),
    .C1(_02612_),
    .X(_02613_));
 sky130_fd_sc_hd__and3_1 _06125_ (.A(_02610_),
    .B(_02611_),
    .C(_02613_),
    .X(_02614_));
 sky130_fd_sc_hd__or2_1 _06126_ (.A(\tms1x00.ins_pla_ands[25][5] ),
    .B(net742),
    .X(_02615_));
 sky130_fd_sc_hd__o221a_1 _06127_ (.A1(\tms1x00.ins_pla_ands[27][5] ),
    .A2(net850),
    .B1(net714),
    .B2(\tms1x00.ins_pla_ands[26][5] ),
    .C1(_02615_),
    .X(_02616_));
 sky130_fd_sc_hd__o221a_1 _06128_ (.A1(\tms1x00.ins_pla_ands[29][5] ),
    .A2(net879),
    .B1(net798),
    .B2(\tms1x00.ins_pla_ands[28][5] ),
    .C1(net990),
    .X(_02617_));
 sky130_fd_sc_hd__o22a_1 _06129_ (.A1(\tms1x00.ins_pla_ands[30][5] ),
    .A2(net603),
    .B1(net769),
    .B2(\tms1x00.ins_pla_ands[31][5] ),
    .X(_02618_));
 sky130_fd_sc_hd__o211a_1 _06130_ (.A1(\tms1x00.ins_pla_ands[24][5] ),
    .A2(net827),
    .B1(_02617_),
    .C1(_02618_),
    .X(_02619_));
 sky130_fd_sc_hd__a211o_2 _06131_ (.A1(_02616_),
    .A2(_02619_),
    .B1(net923),
    .C1(_02614_),
    .X(_02620_));
 sky130_fd_sc_hd__o22a_1 _06132_ (.A1(\tms1x00.ins_pla_ands[14][5] ),
    .A2(net609),
    .B1(net778),
    .B2(\tms1x00.ins_pla_ands[15][5] ),
    .X(_02621_));
 sky130_fd_sc_hd__o22a_1 _06133_ (.A1(\tms1x00.ins_pla_ands[11][5] ),
    .A2(net854),
    .B1(net721),
    .B2(\tms1x00.ins_pla_ands[10][5] ),
    .X(_02622_));
 sky130_fd_sc_hd__o221a_1 _06134_ (.A1(\tms1x00.ins_pla_ands[13][5] ),
    .A2(net882),
    .B1(net802),
    .B2(\tms1x00.ins_pla_ands[12][5] ),
    .C1(net993),
    .X(_02623_));
 sky130_fd_sc_hd__o211a_1 _06135_ (.A1(\tms1x00.ins_pla_ands[9][5] ),
    .A2(net747),
    .B1(_02622_),
    .C1(_02623_),
    .X(_02624_));
 sky130_fd_sc_hd__o211a_1 _06136_ (.A1(\tms1x00.ins_pla_ands[8][5] ),
    .A2(net829),
    .B1(_02621_),
    .C1(_02624_),
    .X(_02625_));
 sky130_fd_sc_hd__o22a_1 _06137_ (.A1(\tms1x00.ins_pla_ands[4][5] ),
    .A2(net812),
    .B1(net732),
    .B2(\tms1x00.ins_pla_ands[2][5] ),
    .X(_02626_));
 sky130_fd_sc_hd__o22a_1 _06138_ (.A1(\tms1x00.ins_pla_ands[3][5] ),
    .A2(net859),
    .B1(net780),
    .B2(\tms1x00.ins_pla_ands[7][5] ),
    .X(_02627_));
 sky130_fd_sc_hd__o221a_1 _06139_ (.A1(\tms1x00.ins_pla_ands[6][5] ),
    .A2(net614),
    .B1(net833),
    .B2(\tms1x00.ins_pla_ands[0][5] ),
    .C1(_02627_),
    .X(_02628_));
 sky130_fd_sc_hd__o211a_1 _06140_ (.A1(\tms1x00.ins_pla_ands[5][5] ),
    .A2(net886),
    .B1(_02628_),
    .C1(net916),
    .X(_02629_));
 sky130_fd_sc_hd__o211a_1 _06141_ (.A1(\tms1x00.ins_pla_ands[1][5] ),
    .A2(net751),
    .B1(_02626_),
    .C1(_02629_),
    .X(_02630_));
 sky130_fd_sc_hd__a211o_1 _06142_ (.A1(net600),
    .A2(_02604_),
    .B1(_02609_),
    .C1(_02593_),
    .X(_02631_));
 sky130_fd_sc_hd__o311a_2 _06143_ (.A1(net986),
    .A2(_02625_),
    .A3(_02630_),
    .B1(net713),
    .C1(_02620_),
    .X(_02632_));
 sky130_fd_sc_hd__a211o_1 _06144_ (.A1(net711),
    .A2(_02631_),
    .B1(_02632_),
    .C1(net586),
    .X(_02633_));
 sky130_fd_sc_hd__o211a_1 _06145_ (.A1(net590),
    .A2(_02571_),
    .B1(_02633_),
    .C1(net630),
    .X(_02634_));
 sky130_fd_sc_hd__a221o_1 _06146_ (.A1(net125),
    .A2(net580),
    .B1(_02571_),
    .B2(net585),
    .C1(_02634_),
    .X(_00032_));
 sky130_fd_sc_hd__o22a_1 _06147_ (.A1(\tms1x00.ins_pla_ands[16][6] ),
    .A2(net825),
    .B1(net770),
    .B2(\tms1x00.ins_pla_ands[23][6] ),
    .X(_02635_));
 sky130_fd_sc_hd__o221a_1 _06148_ (.A1(\tms1x00.ins_pla_ands[21][6] ),
    .A2(net877),
    .B1(net796),
    .B2(\tms1x00.ins_pla_ands[20][6] ),
    .C1(net911),
    .X(_02636_));
 sky130_fd_sc_hd__o22a_1 _06149_ (.A1(\tms1x00.ins_pla_ands[19][6] ),
    .A2(net853),
    .B1(net718),
    .B2(\tms1x00.ins_pla_ands[18][6] ),
    .X(_02637_));
 sky130_fd_sc_hd__o221a_1 _06150_ (.A1(\tms1x00.ins_pla_ands[22][6] ),
    .A2(net604),
    .B1(net746),
    .B2(\tms1x00.ins_pla_ands[17][6] ),
    .C1(_02637_),
    .X(_02638_));
 sky130_fd_sc_hd__and3_1 _06151_ (.A(_02635_),
    .B(_02636_),
    .C(_02638_),
    .X(_02639_));
 sky130_fd_sc_hd__or2_1 _06152_ (.A(\tms1x00.ins_pla_ands[28][6] ),
    .B(net797),
    .X(_02640_));
 sky130_fd_sc_hd__o221a_1 _06153_ (.A1(\tms1x00.ins_pla_ands[31][6] ),
    .A2(net769),
    .B1(net714),
    .B2(\tms1x00.ins_pla_ands[26][6] ),
    .C1(_02640_),
    .X(_02641_));
 sky130_fd_sc_hd__o22a_1 _06154_ (.A1(\tms1x00.ins_pla_ands[29][6] ),
    .A2(net877),
    .B1(net742),
    .B2(\tms1x00.ins_pla_ands[25][6] ),
    .X(_02642_));
 sky130_fd_sc_hd__o221a_1 _06155_ (.A1(\tms1x00.ins_pla_ands[27][6] ),
    .A2(net850),
    .B1(net824),
    .B2(\tms1x00.ins_pla_ands[24][6] ),
    .C1(_02642_),
    .X(_02643_));
 sky130_fd_sc_hd__o211a_1 _06156_ (.A1(\tms1x00.ins_pla_ands[30][6] ),
    .A2(net602),
    .B1(_02643_),
    .C1(net991),
    .X(_02644_));
 sky130_fd_sc_hd__a211o_2 _06157_ (.A1(_02641_),
    .A2(_02644_),
    .B1(net923),
    .C1(_02639_),
    .X(_02645_));
 sky130_fd_sc_hd__o22a_1 _06158_ (.A1(\tms1x00.ins_pla_ands[14][6] ),
    .A2(net609),
    .B1(net774),
    .B2(\tms1x00.ins_pla_ands[15][6] ),
    .X(_02646_));
 sky130_fd_sc_hd__o221a_1 _06159_ (.A1(\tms1x00.ins_pla_ands[13][6] ),
    .A2(net882),
    .B1(net801),
    .B2(\tms1x00.ins_pla_ands[12][6] ),
    .C1(net993),
    .X(_02647_));
 sky130_fd_sc_hd__o22a_1 _06160_ (.A1(\tms1x00.ins_pla_ands[11][6] ),
    .A2(net857),
    .B1(net721),
    .B2(\tms1x00.ins_pla_ands[10][6] ),
    .X(_02648_));
 sky130_fd_sc_hd__o211a_1 _06161_ (.A1(\tms1x00.ins_pla_ands[8][6] ),
    .A2(net831),
    .B1(_02647_),
    .C1(_02648_),
    .X(_02649_));
 sky130_fd_sc_hd__o211a_1 _06162_ (.A1(\tms1x00.ins_pla_ands[9][6] ),
    .A2(net749),
    .B1(_02646_),
    .C1(_02649_),
    .X(_02650_));
 sky130_fd_sc_hd__o22a_1 _06163_ (.A1(\tms1x00.ins_pla_ands[5][6] ),
    .A2(net894),
    .B1(net732),
    .B2(\tms1x00.ins_pla_ands[2][6] ),
    .X(_02651_));
 sky130_fd_sc_hd__o22a_1 _06164_ (.A1(\tms1x00.ins_pla_ands[7][6] ),
    .A2(net780),
    .B1(net750),
    .B2(\tms1x00.ins_pla_ands[1][6] ),
    .X(_02652_));
 sky130_fd_sc_hd__o221a_1 _06165_ (.A1(\tms1x00.ins_pla_ands[6][6] ),
    .A2(net613),
    .B1(net859),
    .B2(\tms1x00.ins_pla_ands[3][6] ),
    .C1(_02652_),
    .X(_02653_));
 sky130_fd_sc_hd__o211a_1 _06166_ (.A1(\tms1x00.ins_pla_ands[4][6] ),
    .A2(net819),
    .B1(_02653_),
    .C1(net916),
    .X(_02654_));
 sky130_fd_sc_hd__o211a_1 _06167_ (.A1(\tms1x00.ins_pla_ands[0][6] ),
    .A2(net833),
    .B1(_02651_),
    .C1(_02654_),
    .X(_02655_));
 sky130_fd_sc_hd__o22a_1 _06168_ (.A1(\tms1x00.O_pla_ands[6][6] ),
    .A2(net622),
    .B1(net788),
    .B2(\tms1x00.O_pla_ands[7][6] ),
    .X(_02656_));
 sky130_fd_sc_hd__o221a_1 _06169_ (.A1(\tms1x00.O_pla_ands[0][6] ),
    .A2(net845),
    .B1(net752),
    .B2(\tms1x00.O_pla_ands[1][6] ),
    .C1(net915),
    .X(_02657_));
 sky130_fd_sc_hd__o22a_1 _06170_ (.A1(\tms1x00.O_pla_ands[3][6] ),
    .A2(net868),
    .B1(net733),
    .B2(\tms1x00.O_pla_ands[2][6] ),
    .X(_02658_));
 sky130_fd_sc_hd__o211a_1 _06171_ (.A1(\tms1x00.O_pla_ands[4][6] ),
    .A2(net813),
    .B1(_02657_),
    .C1(_02658_),
    .X(_02659_));
 sky130_fd_sc_hd__o211a_1 _06172_ (.A1(\tms1x00.O_pla_ands[5][6] ),
    .A2(net896),
    .B1(_02656_),
    .C1(_02659_),
    .X(_02660_));
 sky130_fd_sc_hd__o22a_1 _06173_ (.A1(\tms1x00.O_pla_ands[15][6] ),
    .A2(net790),
    .B1(net736),
    .B2(\tms1x00.O_pla_ands[10][6] ),
    .X(_02661_));
 sky130_fd_sc_hd__o22a_1 _06174_ (.A1(\tms1x00.O_pla_ands[8][6] ),
    .A2(net842),
    .B1(net762),
    .B2(\tms1x00.O_pla_ands[9][6] ),
    .X(_02662_));
 sky130_fd_sc_hd__o221a_1 _06175_ (.A1(\tms1x00.O_pla_ands[13][6] ),
    .A2(net898),
    .B1(net816),
    .B2(\tms1x00.O_pla_ands[12][6] ),
    .C1(_02662_),
    .X(_02663_));
 sky130_fd_sc_hd__o211a_1 _06176_ (.A1(\tms1x00.O_pla_ands[11][6] ),
    .A2(net871),
    .B1(_02663_),
    .C1(net999),
    .X(_02664_));
 sky130_fd_sc_hd__o211a_2 _06177_ (.A1(\tms1x00.O_pla_ands[14][6] ),
    .A2(net624),
    .B1(_02661_),
    .C1(_02664_),
    .X(_02665_));
 sky130_fd_sc_hd__or3_2 _06178_ (.A(net989),
    .B(_02660_),
    .C(_02665_),
    .X(_02666_));
 sky130_fd_sc_hd__o22a_1 _06179_ (.A1(\tms1x00.O_pla_ands[30][6] ),
    .A2(net610),
    .B1(net775),
    .B2(\tms1x00.O_pla_ands[31][6] ),
    .X(_02667_));
 sky130_fd_sc_hd__o221a_1 _06180_ (.A1(\tms1x00.O_pla_ands[29][6] ),
    .A2(net884),
    .B1(net803),
    .B2(\tms1x00.O_pla_ands[28][6] ),
    .C1(net992),
    .X(_02668_));
 sky130_fd_sc_hd__o22a_1 _06181_ (.A1(\tms1x00.O_pla_ands[27][6] ),
    .A2(net855),
    .B1(net722),
    .B2(\tms1x00.O_pla_ands[26][6] ),
    .X(_02669_));
 sky130_fd_sc_hd__o211a_1 _06182_ (.A1(\tms1x00.O_pla_ands[24][6] ),
    .A2(net830),
    .B1(_02668_),
    .C1(_02669_),
    .X(_02670_));
 sky130_fd_sc_hd__o211a_2 _06183_ (.A1(\tms1x00.O_pla_ands[25][6] ),
    .A2(net749),
    .B1(_02667_),
    .C1(_02670_),
    .X(_02671_));
 sky130_fd_sc_hd__o22a_1 _06184_ (.A1(\tms1x00.O_pla_ands[22][6] ),
    .A2(net610),
    .B1(net775),
    .B2(\tms1x00.O_pla_ands[23][6] ),
    .X(_02672_));
 sky130_fd_sc_hd__o221a_1 _06185_ (.A1(\tms1x00.O_pla_ands[16][6] ),
    .A2(net835),
    .B1(net753),
    .B2(\tms1x00.O_pla_ands[17][6] ),
    .C1(net914),
    .X(_02673_));
 sky130_fd_sc_hd__o22a_1 _06186_ (.A1(\tms1x00.O_pla_ands[19][6] ),
    .A2(net858),
    .B1(net724),
    .B2(\tms1x00.O_pla_ands[18][6] ),
    .X(_02674_));
 sky130_fd_sc_hd__o211a_1 _06187_ (.A1(\tms1x00.O_pla_ands[21][6] ),
    .A2(net885),
    .B1(_02673_),
    .C1(_02674_),
    .X(_02675_));
 sky130_fd_sc_hd__o211a_1 _06188_ (.A1(\tms1x00.O_pla_ands[20][6] ),
    .A2(net805),
    .B1(_02672_),
    .C1(_02675_),
    .X(_02676_));
 sky130_fd_sc_hd__o311a_2 _06189_ (.A1(net926),
    .A2(_02671_),
    .A3(_02676_),
    .B1(net905),
    .C1(_02666_),
    .X(_02677_));
 sky130_fd_sc_hd__or2_1 _06190_ (.A(\tms1x00.ins_pla_ors[4][6] ),
    .B(net810),
    .X(_02678_));
 sky130_fd_sc_hd__o22a_2 _06191_ (.A1(\tms1x00.ins_pla_ors[1][6] ),
    .A2(net760),
    .B1(net731),
    .B2(\tms1x00.ins_pla_ors[2][6] ),
    .X(_02679_));
 sky130_fd_sc_hd__o22a_1 _06192_ (.A1(\tms1x00.ins_pla_ors[3][6] ),
    .A2(net864),
    .B1(net786),
    .B2(\tms1x00.ins_pla_ors[7][6] ),
    .X(_02680_));
 sky130_fd_sc_hd__o221a_2 _06193_ (.A1(\tms1x00.ins_pla_ors[6][6] ),
    .A2(net619),
    .B1(net840),
    .B2(\tms1x00.ins_pla_ors[0][6] ),
    .C1(_02680_),
    .X(_02681_));
 sky130_fd_sc_hd__o211a_1 _06194_ (.A1(\tms1x00.ins_pla_ors[5][6] ),
    .A2(net893),
    .B1(_02681_),
    .C1(net920),
    .X(_02682_));
 sky130_fd_sc_hd__o22a_1 _06195_ (.A1(\tms1x00.ins_pla_ors[13][6] ),
    .A2(net889),
    .B1(net863),
    .B2(\tms1x00.ins_pla_ors[11][6] ),
    .X(_02683_));
 sky130_fd_sc_hd__o22a_1 _06196_ (.A1(\tms1x00.ins_pla_ors[8][6] ),
    .A2(net838),
    .B1(net756),
    .B2(\tms1x00.ins_pla_ors[9][6] ),
    .X(_02684_));
 sky130_fd_sc_hd__o221a_1 _06197_ (.A1(\tms1x00.ins_pla_ors[15][6] ),
    .A2(net783),
    .B1(net727),
    .B2(\tms1x00.ins_pla_ors[10][6] ),
    .C1(_02684_),
    .X(_02685_));
 sky130_fd_sc_hd__o211a_1 _06198_ (.A1(\tms1x00.ins_pla_ors[14][6] ),
    .A2(net617),
    .B1(_02685_),
    .C1(net996),
    .X(_02686_));
 sky130_fd_sc_hd__o211a_1 _06199_ (.A1(\tms1x00.ins_pla_ors[12][6] ),
    .A2(net807),
    .B1(_02683_),
    .C1(_02686_),
    .X(_02687_));
 sky130_fd_sc_hd__a31o_4 _06200_ (.A1(_02678_),
    .A2(_02679_),
    .A3(_02682_),
    .B1(_02687_),
    .X(_02688_));
 sky130_fd_sc_hd__o22a_1 _06201_ (.A1(\tms1x00.O_pla_ors[3][6] ),
    .A2(net872),
    .B1(net792),
    .B2(\tms1x00.O_pla_ors[7][6] ),
    .X(_02689_));
 sky130_fd_sc_hd__o22a_1 _06202_ (.A1(\tms1x00.O_pla_ors[5][6] ),
    .A2(net899),
    .B1(net817),
    .B2(\tms1x00.O_pla_ors[4][6] ),
    .X(_02690_));
 sky130_fd_sc_hd__o221a_1 _06203_ (.A1(\tms1x00.O_pla_ors[6][6] ),
    .A2(net625),
    .B1(net764),
    .B2(\tms1x00.O_pla_ors[1][6] ),
    .C1(_02690_),
    .X(_02691_));
 sky130_fd_sc_hd__o211a_1 _06204_ (.A1(\tms1x00.O_pla_ors[0][6] ),
    .A2(net844),
    .B1(net599),
    .C1(_02691_),
    .X(_02692_));
 sky130_fd_sc_hd__o211a_4 _06205_ (.A1(\tms1x00.O_pla_ors[2][6] ),
    .A2(net737),
    .B1(_02689_),
    .C1(_02692_),
    .X(_02693_));
 sky130_fd_sc_hd__a211o_1 _06206_ (.A1(net600),
    .A2(_02688_),
    .B1(_02693_),
    .C1(_02677_),
    .X(_02694_));
 sky130_fd_sc_hd__o311a_2 _06207_ (.A1(net986),
    .A2(_02650_),
    .A3(_02655_),
    .B1(net712),
    .C1(_02645_),
    .X(_02695_));
 sky130_fd_sc_hd__a211o_1 _06208_ (.A1(net711),
    .A2(_02694_),
    .B1(_02695_),
    .C1(net587),
    .X(_02696_));
 sky130_fd_sc_hd__a21o_1 _06209_ (.A1(net907),
    .A2(\wbs_o_buff[6] ),
    .B1(net589),
    .X(_02697_));
 sky130_fd_sc_hd__a32o_1 _06210_ (.A1(net629),
    .A2(_02696_),
    .A3(_02697_),
    .B1(net579),
    .B2(net126),
    .X(_02698_));
 sky130_fd_sc_hd__a31o_1 _06211_ (.A1(net907),
    .A2(\wbs_o_buff[6] ),
    .A3(net585),
    .B1(_02698_),
    .X(_00033_));
 sky130_fd_sc_hd__nand2_1 _06212_ (.A(net906),
    .B(\wbs_o_buff[7] ),
    .Y(_02699_));
 sky130_fd_sc_hd__o22a_1 _06213_ (.A1(\tms1x00.O_pla_ands[6][7] ),
    .A2(net623),
    .B1(net789),
    .B2(\tms1x00.O_pla_ands[7][7] ),
    .X(_02700_));
 sky130_fd_sc_hd__o221a_2 _06214_ (.A1(\tms1x00.O_pla_ands[0][7] ),
    .A2(net834),
    .B1(net754),
    .B2(\tms1x00.O_pla_ands[1][7] ),
    .C1(net915),
    .X(_02701_));
 sky130_fd_sc_hd__o22a_1 _06215_ (.A1(\tms1x00.O_pla_ands[3][7] ),
    .A2(net869),
    .B1(net734),
    .B2(\tms1x00.O_pla_ands[2][7] ),
    .X(_02702_));
 sky130_fd_sc_hd__o211a_1 _06216_ (.A1(\tms1x00.O_pla_ands[5][7] ),
    .A2(net897),
    .B1(_02701_),
    .C1(_02702_),
    .X(_02703_));
 sky130_fd_sc_hd__o211a_1 _06217_ (.A1(\tms1x00.O_pla_ands[4][7] ),
    .A2(net814),
    .B1(_02700_),
    .C1(_02703_),
    .X(_02704_));
 sky130_fd_sc_hd__or2_1 _06218_ (.A(\tms1x00.O_pla_ands[14][7] ),
    .B(net623),
    .X(_02705_));
 sky130_fd_sc_hd__o22a_1 _06219_ (.A1(\tms1x00.O_pla_ands[13][7] ),
    .A2(net897),
    .B1(net765),
    .B2(\tms1x00.O_pla_ands[9][7] ),
    .X(_02706_));
 sky130_fd_sc_hd__o22a_1 _06220_ (.A1(\tms1x00.O_pla_ands[8][7] ),
    .A2(net844),
    .B1(net791),
    .B2(\tms1x00.O_pla_ands[15][7] ),
    .X(_02707_));
 sky130_fd_sc_hd__o221a_2 _06221_ (.A1(\tms1x00.O_pla_ands[12][7] ),
    .A2(net817),
    .B1(net735),
    .B2(\tms1x00.O_pla_ands[10][7] ),
    .C1(_02707_),
    .X(_02708_));
 sky130_fd_sc_hd__o211a_1 _06222_ (.A1(\tms1x00.O_pla_ands[11][7] ),
    .A2(net869),
    .B1(_02708_),
    .C1(net1000),
    .X(_02709_));
 sky130_fd_sc_hd__a31o_1 _06223_ (.A1(_02705_),
    .A2(_02706_),
    .A3(_02709_),
    .B1(_02704_),
    .X(_02710_));
 sky130_fd_sc_hd__o22a_1 _06224_ (.A1(\tms1x00.O_pla_ands[24][7] ),
    .A2(net830),
    .B1(net777),
    .B2(\tms1x00.O_pla_ands[31][7] ),
    .X(_02711_));
 sky130_fd_sc_hd__o22a_1 _06225_ (.A1(\tms1x00.O_pla_ands[27][7] ),
    .A2(net855),
    .B1(net722),
    .B2(\tms1x00.O_pla_ands[26][7] ),
    .X(_02712_));
 sky130_fd_sc_hd__o221a_1 _06226_ (.A1(\tms1x00.O_pla_ands[30][7] ),
    .A2(net611),
    .B1(net748),
    .B2(\tms1x00.O_pla_ands[25][7] ),
    .C1(_02712_),
    .X(_02713_));
 sky130_fd_sc_hd__o221a_1 _06227_ (.A1(\tms1x00.O_pla_ands[29][7] ),
    .A2(net886),
    .B1(net804),
    .B2(\tms1x00.O_pla_ands[28][7] ),
    .C1(net992),
    .X(_02714_));
 sky130_fd_sc_hd__o22a_2 _06228_ (.A1(\tms1x00.O_pla_ands[22][7] ),
    .A2(net612),
    .B1(net776),
    .B2(\tms1x00.O_pla_ands[23][7] ),
    .X(_02715_));
 sky130_fd_sc_hd__o221a_1 _06229_ (.A1(\tms1x00.O_pla_ands[16][7] ),
    .A2(net834),
    .B1(net753),
    .B2(\tms1x00.O_pla_ands[17][7] ),
    .C1(net914),
    .X(_02716_));
 sky130_fd_sc_hd__o22a_1 _06230_ (.A1(\tms1x00.O_pla_ands[19][7] ),
    .A2(net860),
    .B1(net725),
    .B2(\tms1x00.O_pla_ands[18][7] ),
    .X(_02717_));
 sky130_fd_sc_hd__o211a_1 _06231_ (.A1(\tms1x00.O_pla_ands[21][7] ),
    .A2(net885),
    .B1(_02716_),
    .C1(_02717_),
    .X(_02718_));
 sky130_fd_sc_hd__o211a_2 _06232_ (.A1(\tms1x00.O_pla_ands[20][7] ),
    .A2(net805),
    .B1(_02715_),
    .C1(_02718_),
    .X(_02719_));
 sky130_fd_sc_hd__a31o_4 _06233_ (.A1(_02711_),
    .A2(_02713_),
    .A3(_02714_),
    .B1(net925),
    .X(_02720_));
 sky130_fd_sc_hd__o221a_2 _06234_ (.A1(net989),
    .A2(_02710_),
    .B1(_02719_),
    .B2(_02720_),
    .C1(net905),
    .X(_02721_));
 sky130_fd_sc_hd__o22a_1 _06235_ (.A1(\tms1x00.ins_pla_ors[13][7] ),
    .A2(net881),
    .B1(net853),
    .B2(\tms1x00.ins_pla_ors[11][7] ),
    .X(_02722_));
 sky130_fd_sc_hd__o22a_1 _06236_ (.A1(\tms1x00.ins_pla_ors[12][7] ),
    .A2(net807),
    .B1(net757),
    .B2(\tms1x00.ins_pla_ors[9][7] ),
    .X(_02723_));
 sky130_fd_sc_hd__o221a_1 _06237_ (.A1(\tms1x00.ins_pla_ors[15][7] ),
    .A2(net773),
    .B1(net718),
    .B2(\tms1x00.ins_pla_ors[10][7] ),
    .C1(_02723_),
    .X(_02724_));
 sky130_fd_sc_hd__o211a_1 _06238_ (.A1(\tms1x00.ins_pla_ors[8][7] ),
    .A2(net828),
    .B1(_02724_),
    .C1(net991),
    .X(_02725_));
 sky130_fd_sc_hd__o211a_2 _06239_ (.A1(\tms1x00.ins_pla_ors[14][7] ),
    .A2(net606),
    .B1(_02722_),
    .C1(_02725_),
    .X(_02726_));
 sky130_fd_sc_hd__or2_1 _06240_ (.A(\tms1x00.ins_pla_ors[5][7] ),
    .B(net889),
    .X(_02727_));
 sky130_fd_sc_hd__o22a_1 _06241_ (.A1(\tms1x00.ins_pla_ors[0][7] ),
    .A2(net840),
    .B1(net786),
    .B2(\tms1x00.ins_pla_ors[7][7] ),
    .X(_02728_));
 sky130_fd_sc_hd__o22a_1 _06242_ (.A1(\tms1x00.ins_pla_ors[3][7] ),
    .A2(net866),
    .B1(net759),
    .B2(\tms1x00.ins_pla_ors[1][7] ),
    .X(_02729_));
 sky130_fd_sc_hd__o221a_1 _06243_ (.A1(\tms1x00.ins_pla_ors[6][7] ),
    .A2(net619),
    .B1(net730),
    .B2(\tms1x00.ins_pla_ors[2][7] ),
    .C1(_02729_),
    .X(_02730_));
 sky130_fd_sc_hd__o211a_1 _06244_ (.A1(\tms1x00.ins_pla_ors[4][7] ),
    .A2(net810),
    .B1(_02730_),
    .C1(net920),
    .X(_02731_));
 sky130_fd_sc_hd__a31o_1 _06245_ (.A1(_02727_),
    .A2(_02728_),
    .A3(_02731_),
    .B1(_02726_),
    .X(_02732_));
 sky130_fd_sc_hd__o22a_1 _06246_ (.A1(\tms1x00.O_pla_ors[0][7] ),
    .A2(net844),
    .B1(net818),
    .B2(\tms1x00.O_pla_ors[4][7] ),
    .X(_02733_));
 sky130_fd_sc_hd__o22a_1 _06247_ (.A1(\tms1x00.O_pla_ors[7][7] ),
    .A2(net792),
    .B1(net737),
    .B2(\tms1x00.O_pla_ors[2][7] ),
    .X(_02734_));
 sky130_fd_sc_hd__o221a_1 _06248_ (.A1(\tms1x00.O_pla_ors[5][7] ),
    .A2(net900),
    .B1(net872),
    .B2(\tms1x00.O_pla_ors[3][7] ),
    .C1(_02734_),
    .X(_02735_));
 sky130_fd_sc_hd__o211a_1 _06249_ (.A1(\tms1x00.O_pla_ors[1][7] ),
    .A2(net764),
    .B1(net599),
    .C1(_02735_),
    .X(_02736_));
 sky130_fd_sc_hd__o211a_1 _06250_ (.A1(\tms1x00.O_pla_ors[6][7] ),
    .A2(net625),
    .B1(_02733_),
    .C1(_02736_),
    .X(_02737_));
 sky130_fd_sc_hd__o22a_1 _06251_ (.A1(\tms1x00.ins_pla_ands[16][7] ),
    .A2(net826),
    .B1(net770),
    .B2(\tms1x00.ins_pla_ands[23][7] ),
    .X(_02738_));
 sky130_fd_sc_hd__o221a_1 _06252_ (.A1(\tms1x00.ins_pla_ands[21][7] ),
    .A2(net877),
    .B1(net796),
    .B2(\tms1x00.ins_pla_ands[20][7] ),
    .C1(net911),
    .X(_02739_));
 sky130_fd_sc_hd__o22a_1 _06253_ (.A1(\tms1x00.ins_pla_ands[19][7] ),
    .A2(net853),
    .B1(net718),
    .B2(\tms1x00.ins_pla_ands[18][7] ),
    .X(_02740_));
 sky130_fd_sc_hd__o221a_1 _06254_ (.A1(\tms1x00.ins_pla_ands[22][7] ),
    .A2(net606),
    .B1(net746),
    .B2(\tms1x00.ins_pla_ands[17][7] ),
    .C1(_02740_),
    .X(_02741_));
 sky130_fd_sc_hd__and3_1 _06255_ (.A(_02738_),
    .B(_02739_),
    .C(_02741_),
    .X(_02742_));
 sky130_fd_sc_hd__or2_1 _06256_ (.A(\tms1x00.ins_pla_ands[31][7] ),
    .B(net771),
    .X(_02743_));
 sky130_fd_sc_hd__o221a_1 _06257_ (.A1(\tms1x00.ins_pla_ands[30][7] ),
    .A2(net603),
    .B1(net796),
    .B2(\tms1x00.ins_pla_ands[28][7] ),
    .C1(_02743_),
    .X(_02744_));
 sky130_fd_sc_hd__o22a_1 _06258_ (.A1(\tms1x00.ins_pla_ands[29][7] ),
    .A2(net877),
    .B1(net714),
    .B2(\tms1x00.ins_pla_ands[26][7] ),
    .X(_02745_));
 sky130_fd_sc_hd__o221a_1 _06259_ (.A1(\tms1x00.ins_pla_ands[24][7] ),
    .A2(net823),
    .B1(net742),
    .B2(\tms1x00.ins_pla_ands[25][7] ),
    .C1(_02745_),
    .X(_02746_));
 sky130_fd_sc_hd__o211a_1 _06260_ (.A1(\tms1x00.ins_pla_ands[27][7] ),
    .A2(net850),
    .B1(_02746_),
    .C1(net991),
    .X(_02747_));
 sky130_fd_sc_hd__a211o_2 _06261_ (.A1(_02744_),
    .A2(_02747_),
    .B1(net923),
    .C1(_02742_),
    .X(_02748_));
 sky130_fd_sc_hd__o22a_1 _06262_ (.A1(\tms1x00.ins_pla_ands[6][7] ),
    .A2(net613),
    .B1(net750),
    .B2(\tms1x00.ins_pla_ands[1][7] ),
    .X(_02749_));
 sky130_fd_sc_hd__o22a_1 _06263_ (.A1(\tms1x00.ins_pla_ands[0][7] ),
    .A2(net845),
    .B1(net812),
    .B2(\tms1x00.ins_pla_ands[4][7] ),
    .X(_02750_));
 sky130_fd_sc_hd__o221a_1 _06264_ (.A1(\tms1x00.ins_pla_ands[5][7] ),
    .A2(net894),
    .B1(net732),
    .B2(\tms1x00.ins_pla_ands[2][7] ),
    .C1(_02750_),
    .X(_02751_));
 sky130_fd_sc_hd__o211a_1 _06265_ (.A1(\tms1x00.ins_pla_ands[7][7] ),
    .A2(net780),
    .B1(_02751_),
    .C1(net916),
    .X(_02752_));
 sky130_fd_sc_hd__o211a_1 _06266_ (.A1(\tms1x00.ins_pla_ands[3][7] ),
    .A2(net859),
    .B1(_02749_),
    .C1(_02752_),
    .X(_02753_));
 sky130_fd_sc_hd__o22a_1 _06267_ (.A1(\tms1x00.ins_pla_ands[14][7] ),
    .A2(net614),
    .B1(net779),
    .B2(\tms1x00.ins_pla_ands[15][7] ),
    .X(_02754_));
 sky130_fd_sc_hd__o221a_1 _06268_ (.A1(\tms1x00.ins_pla_ands[13][7] ),
    .A2(net883),
    .B1(net802),
    .B2(\tms1x00.ins_pla_ands[12][7] ),
    .C1(net993),
    .X(_02755_));
 sky130_fd_sc_hd__o22a_1 _06269_ (.A1(\tms1x00.ins_pla_ands[11][7] ),
    .A2(net857),
    .B1(net721),
    .B2(\tms1x00.ins_pla_ands[10][7] ),
    .X(_02756_));
 sky130_fd_sc_hd__o211a_1 _06270_ (.A1(\tms1x00.ins_pla_ands[9][7] ),
    .A2(net747),
    .B1(_02755_),
    .C1(_02756_),
    .X(_02757_));
 sky130_fd_sc_hd__o211a_1 _06271_ (.A1(\tms1x00.ins_pla_ands[8][7] ),
    .A2(net832),
    .B1(_02754_),
    .C1(_02757_),
    .X(_02758_));
 sky130_fd_sc_hd__a211o_4 _06272_ (.A1(net600),
    .A2(_02732_),
    .B1(_02737_),
    .C1(_02721_),
    .X(_02759_));
 sky130_fd_sc_hd__o311a_1 _06273_ (.A1(net986),
    .A2(_02753_),
    .A3(_02758_),
    .B1(net712),
    .C1(_02748_),
    .X(_02760_));
 sky130_fd_sc_hd__a211o_1 _06274_ (.A1(net711),
    .A2(_02759_),
    .B1(_02760_),
    .C1(net586),
    .X(_02761_));
 sky130_fd_sc_hd__a21oi_1 _06275_ (.A1(net586),
    .A2(_02699_),
    .B1(_02223_),
    .Y(_02762_));
 sky130_fd_sc_hd__a22o_1 _06276_ (.A1(net127),
    .A2(net579),
    .B1(_02761_),
    .B2(_02762_),
    .X(_02763_));
 sky130_fd_sc_hd__a31o_1 _06277_ (.A1(net906),
    .A2(\wbs_o_buff[7] ),
    .A3(net582),
    .B1(_02763_),
    .X(_00034_));
 sky130_fd_sc_hd__o22a_1 _06278_ (.A1(\tms1x00.O_pla_ands[30][8] ),
    .A2(net611),
    .B1(net775),
    .B2(\tms1x00.O_pla_ands[31][8] ),
    .X(_02764_));
 sky130_fd_sc_hd__o221a_1 _06279_ (.A1(\tms1x00.O_pla_ands[29][8] ),
    .A2(net884),
    .B1(net803),
    .B2(\tms1x00.O_pla_ands[28][8] ),
    .C1(net992),
    .X(_02765_));
 sky130_fd_sc_hd__o22a_1 _06280_ (.A1(\tms1x00.O_pla_ands[27][8] ),
    .A2(net855),
    .B1(net722),
    .B2(\tms1x00.O_pla_ands[26][8] ),
    .X(_02766_));
 sky130_fd_sc_hd__o211a_1 _06281_ (.A1(\tms1x00.O_pla_ands[24][8] ),
    .A2(net830),
    .B1(_02765_),
    .C1(_02766_),
    .X(_02767_));
 sky130_fd_sc_hd__o211a_1 _06282_ (.A1(\tms1x00.O_pla_ands[25][8] ),
    .A2(net748),
    .B1(_02764_),
    .C1(_02767_),
    .X(_02768_));
 sky130_fd_sc_hd__o22a_1 _06283_ (.A1(\tms1x00.O_pla_ands[21][8] ),
    .A2(net885),
    .B1(net723),
    .B2(\tms1x00.O_pla_ands[18][8] ),
    .X(_02769_));
 sky130_fd_sc_hd__o221a_1 _06284_ (.A1(\tms1x00.O_pla_ands[22][8] ),
    .A2(net610),
    .B1(net775),
    .B2(\tms1x00.O_pla_ands[23][8] ),
    .C1(_02769_),
    .X(_02770_));
 sky130_fd_sc_hd__o221a_1 _06285_ (.A1(\tms1x00.O_pla_ands[16][8] ),
    .A2(net835),
    .B1(net753),
    .B2(\tms1x00.O_pla_ands[17][8] ),
    .C1(net917),
    .X(_02771_));
 sky130_fd_sc_hd__o221a_1 _06286_ (.A1(\tms1x00.O_pla_ands[19][8] ),
    .A2(net858),
    .B1(net805),
    .B2(\tms1x00.O_pla_ands[20][8] ),
    .C1(_02771_),
    .X(_02772_));
 sky130_fd_sc_hd__a211o_4 _06287_ (.A1(_02770_),
    .A2(_02772_),
    .B1(net925),
    .C1(_02768_),
    .X(_02773_));
 sky130_fd_sc_hd__nor2_2 _06288_ (.A(net985),
    .B(_01637_),
    .Y(_02774_));
 sky130_fd_sc_hd__nand2_1 _06289_ (.A(net905),
    .B(net984),
    .Y(_02775_));
 sky130_fd_sc_hd__o22a_1 _06290_ (.A1(\tms1x00.O_pla_ands[13][8] ),
    .A2(net898),
    .B1(net735),
    .B2(\tms1x00.O_pla_ands[10][8] ),
    .X(_02776_));
 sky130_fd_sc_hd__o22a_1 _06291_ (.A1(\tms1x00.O_pla_ands[15][8] ),
    .A2(net790),
    .B1(net763),
    .B2(\tms1x00.O_pla_ands[9][8] ),
    .X(_02777_));
 sky130_fd_sc_hd__o221a_1 _06292_ (.A1(\tms1x00.O_pla_ands[14][8] ),
    .A2(net624),
    .B1(net871),
    .B2(\tms1x00.O_pla_ands[11][8] ),
    .C1(_02777_),
    .X(_02778_));
 sky130_fd_sc_hd__o211a_1 _06293_ (.A1(\tms1x00.O_pla_ands[12][8] ),
    .A2(net816),
    .B1(_02778_),
    .C1(net1000),
    .X(_02779_));
 sky130_fd_sc_hd__o211a_2 _06294_ (.A1(\tms1x00.O_pla_ands[8][8] ),
    .A2(net843),
    .B1(_02776_),
    .C1(_02779_),
    .X(_02780_));
 sky130_fd_sc_hd__o22a_1 _06295_ (.A1(\tms1x00.O_pla_ands[3][8] ),
    .A2(net868),
    .B1(net733),
    .B2(\tms1x00.O_pla_ands[2][8] ),
    .X(_02781_));
 sky130_fd_sc_hd__o221a_1 _06296_ (.A1(\tms1x00.O_pla_ands[6][8] ),
    .A2(net622),
    .B1(net765),
    .B2(\tms1x00.O_pla_ands[1][8] ),
    .C1(_02781_),
    .X(_02782_));
 sky130_fd_sc_hd__o221a_1 _06297_ (.A1(\tms1x00.O_pla_ands[5][8] ),
    .A2(net896),
    .B1(net813),
    .B2(\tms1x00.O_pla_ands[4][8] ),
    .C1(net922),
    .X(_02783_));
 sky130_fd_sc_hd__o221a_1 _06298_ (.A1(\tms1x00.O_pla_ands[0][8] ),
    .A2(net845),
    .B1(net788),
    .B2(\tms1x00.O_pla_ands[7][8] ),
    .C1(_02783_),
    .X(_02784_));
 sky130_fd_sc_hd__a211o_1 _06299_ (.A1(_02782_),
    .A2(_02784_),
    .B1(net988),
    .C1(_02780_),
    .X(_02785_));
 sky130_fd_sc_hd__or2_1 _06300_ (.A(\tms1x00.ins_pla_ors[1][8] ),
    .B(net759),
    .X(_02786_));
 sky130_fd_sc_hd__o22a_1 _06301_ (.A1(\tms1x00.ins_pla_ors[3][8] ),
    .A2(net866),
    .B1(net786),
    .B2(\tms1x00.ins_pla_ors[7][8] ),
    .X(_02787_));
 sky130_fd_sc_hd__o22a_1 _06302_ (.A1(\tms1x00.ins_pla_ors[5][8] ),
    .A2(net892),
    .B1(net840),
    .B2(\tms1x00.ins_pla_ors[0][8] ),
    .X(_02788_));
 sky130_fd_sc_hd__o221a_1 _06303_ (.A1(\tms1x00.ins_pla_ors[4][8] ),
    .A2(net810),
    .B1(net730),
    .B2(\tms1x00.ins_pla_ors[2][8] ),
    .C1(_02788_),
    .X(_02789_));
 sky130_fd_sc_hd__o211a_1 _06304_ (.A1(\tms1x00.ins_pla_ors[6][8] ),
    .A2(net619),
    .B1(_02789_),
    .C1(net919),
    .X(_02790_));
 sky130_fd_sc_hd__o22a_1 _06305_ (.A1(\tms1x00.ins_pla_ors[13][8] ),
    .A2(net881),
    .B1(net718),
    .B2(\tms1x00.ins_pla_ors[10][8] ),
    .X(_02791_));
 sky130_fd_sc_hd__o22a_1 _06306_ (.A1(\tms1x00.ins_pla_ors[11][8] ),
    .A2(net863),
    .B1(net807),
    .B2(\tms1x00.ins_pla_ors[12][8] ),
    .X(_02792_));
 sky130_fd_sc_hd__o221a_1 _06307_ (.A1(\tms1x00.ins_pla_ors[8][8] ),
    .A2(net838),
    .B1(net757),
    .B2(\tms1x00.ins_pla_ors[9][8] ),
    .C1(net996),
    .X(_02793_));
 sky130_fd_sc_hd__o221a_2 _06308_ (.A1(\tms1x00.ins_pla_ors[14][8] ),
    .A2(net606),
    .B1(net773),
    .B2(\tms1x00.ins_pla_ors[15][8] ),
    .C1(_02791_),
    .X(_02794_));
 sky130_fd_sc_hd__and3_2 _06309_ (.A(_02792_),
    .B(_02793_),
    .C(_02794_),
    .X(_02795_));
 sky130_fd_sc_hd__a31o_2 _06310_ (.A1(_02786_),
    .A2(_02787_),
    .A3(_02790_),
    .B1(_02795_),
    .X(_02796_));
 sky130_fd_sc_hd__o22a_1 _06311_ (.A1(\tms1x00.O_pla_ors[6][8] ),
    .A2(net623),
    .B1(net788),
    .B2(\tms1x00.O_pla_ors[7][8] ),
    .X(_02797_));
 sky130_fd_sc_hd__o221a_1 _06312_ (.A1(\tms1x00.O_pla_ors[0][8] ),
    .A2(net842),
    .B1(net762),
    .B2(\tms1x00.O_pla_ors[1][8] ),
    .C1(net599),
    .X(_02798_));
 sky130_fd_sc_hd__o22a_1 _06313_ (.A1(\tms1x00.O_pla_ors[3][8] ),
    .A2(net871),
    .B1(net735),
    .B2(\tms1x00.O_pla_ors[2][8] ),
    .X(_02799_));
 sky130_fd_sc_hd__o211a_1 _06314_ (.A1(\tms1x00.O_pla_ors[5][8] ),
    .A2(net898),
    .B1(_02798_),
    .C1(_02799_),
    .X(_02800_));
 sky130_fd_sc_hd__o211a_1 _06315_ (.A1(\tms1x00.O_pla_ors[4][8] ),
    .A2(net814),
    .B1(_02797_),
    .C1(_02800_),
    .X(_02801_));
 sky130_fd_sc_hd__a211o_2 _06316_ (.A1(net601),
    .A2(_02796_),
    .B1(_02801_),
    .C1(net713),
    .X(_02802_));
 sky130_fd_sc_hd__a31o_1 _06317_ (.A1(_02773_),
    .A2(_02774_),
    .A3(_02785_),
    .B1(_02802_),
    .X(_02803_));
 sky130_fd_sc_hd__o22a_1 _06318_ (.A1(\tms1x00.ins_pla_ands[6][8] ),
    .A2(net614),
    .B1(net779),
    .B2(\tms1x00.ins_pla_ands[7][8] ),
    .X(_02804_));
 sky130_fd_sc_hd__o221a_1 _06319_ (.A1(\tms1x00.ins_pla_ands[5][8] ),
    .A2(net895),
    .B1(net812),
    .B2(\tms1x00.ins_pla_ands[4][8] ),
    .C1(net921),
    .X(_02805_));
 sky130_fd_sc_hd__o22a_1 _06320_ (.A1(\tms1x00.ins_pla_ands[3][8] ),
    .A2(net859),
    .B1(net725),
    .B2(\tms1x00.ins_pla_ands[2][8] ),
    .X(_02806_));
 sky130_fd_sc_hd__o211a_1 _06321_ (.A1(\tms1x00.ins_pla_ands[1][8] ),
    .A2(net750),
    .B1(_02805_),
    .C1(_02806_),
    .X(_02807_));
 sky130_fd_sc_hd__o211a_2 _06322_ (.A1(\tms1x00.ins_pla_ands[0][8] ),
    .A2(net833),
    .B1(_02804_),
    .C1(_02807_),
    .X(_02808_));
 sky130_fd_sc_hd__o22a_1 _06323_ (.A1(\tms1x00.ins_pla_ands[11][8] ),
    .A2(net854),
    .B1(net774),
    .B2(\tms1x00.ins_pla_ands[15][8] ),
    .X(_02809_));
 sky130_fd_sc_hd__o22a_1 _06324_ (.A1(\tms1x00.ins_pla_ands[8][8] ),
    .A2(net829),
    .B1(net802),
    .B2(\tms1x00.ins_pla_ands[12][8] ),
    .X(_02810_));
 sky130_fd_sc_hd__o221a_1 _06325_ (.A1(\tms1x00.ins_pla_ands[14][8] ),
    .A2(net608),
    .B1(net720),
    .B2(\tms1x00.ins_pla_ands[10][8] ),
    .C1(_02810_),
    .X(_02811_));
 sky130_fd_sc_hd__o211a_1 _06326_ (.A1(\tms1x00.ins_pla_ands[9][8] ),
    .A2(net747),
    .B1(_02811_),
    .C1(net993),
    .X(_02812_));
 sky130_fd_sc_hd__o211a_1 _06327_ (.A1(\tms1x00.ins_pla_ands[13][8] ),
    .A2(net883),
    .B1(_02809_),
    .C1(_02812_),
    .X(_02813_));
 sky130_fd_sc_hd__o221a_1 _06328_ (.A1(\tms1x00.ins_pla_ands[21][8] ),
    .A2(net878),
    .B1(net797),
    .B2(\tms1x00.ins_pla_ands[20][8] ),
    .C1(net911),
    .X(_02814_));
 sky130_fd_sc_hd__o22a_1 _06329_ (.A1(\tms1x00.ins_pla_ands[19][8] ),
    .A2(net851),
    .B1(net715),
    .B2(\tms1x00.ins_pla_ands[18][8] ),
    .X(_02815_));
 sky130_fd_sc_hd__o221a_1 _06330_ (.A1(\tms1x00.ins_pla_ands[22][8] ),
    .A2(net604),
    .B1(net744),
    .B2(\tms1x00.ins_pla_ands[17][8] ),
    .C1(_02815_),
    .X(_02816_));
 sky130_fd_sc_hd__o221a_1 _06331_ (.A1(\tms1x00.ins_pla_ands[16][8] ),
    .A2(net825),
    .B1(net770),
    .B2(\tms1x00.ins_pla_ands[23][8] ),
    .C1(_02816_),
    .X(_02817_));
 sky130_fd_sc_hd__o22a_1 _06332_ (.A1(\tms1x00.ins_pla_ands[30][8] ),
    .A2(net602),
    .B1(net769),
    .B2(\tms1x00.ins_pla_ands[31][8] ),
    .X(_02818_));
 sky130_fd_sc_hd__o221a_1 _06333_ (.A1(\tms1x00.ins_pla_ands[29][8] ),
    .A2(net879),
    .B1(net798),
    .B2(\tms1x00.ins_pla_ands[28][8] ),
    .C1(net990),
    .X(_02819_));
 sky130_fd_sc_hd__o22a_1 _06334_ (.A1(\tms1x00.ins_pla_ands[27][8] ),
    .A2(net852),
    .B1(net717),
    .B2(\tms1x00.ins_pla_ands[26][8] ),
    .X(_02820_));
 sky130_fd_sc_hd__o211a_1 _06335_ (.A1(\tms1x00.ins_pla_ands[24][8] ),
    .A2(net823),
    .B1(_02819_),
    .C1(_02820_),
    .X(_02821_));
 sky130_fd_sc_hd__o211a_1 _06336_ (.A1(\tms1x00.ins_pla_ands[25][8] ),
    .A2(net742),
    .B1(_02818_),
    .C1(_02821_),
    .X(_02822_));
 sky130_fd_sc_hd__a21o_2 _06337_ (.A1(_02814_),
    .A2(_02817_),
    .B1(_02822_),
    .X(_02823_));
 sky130_fd_sc_hd__o21a_1 _06338_ (.A1(_02808_),
    .A2(_02813_),
    .B1(net925),
    .X(_02824_));
 sky130_fd_sc_hd__a211o_4 _06339_ (.A1(net987),
    .A2(_02823_),
    .B1(_02824_),
    .C1(net711),
    .X(_02825_));
 sky130_fd_sc_hd__a31o_1 _06340_ (.A1(net907),
    .A2(\wbs_o_buff[8] ),
    .A3(net587),
    .B1(net579),
    .X(_02826_));
 sky130_fd_sc_hd__a31o_1 _06341_ (.A1(net589),
    .A2(_02803_),
    .A3(_02825_),
    .B1(_02826_),
    .X(_02827_));
 sky130_fd_sc_hd__o21a_1 _06342_ (.A1(net128),
    .A2(_02314_),
    .B1(_02827_),
    .X(_00035_));
 sky130_fd_sc_hd__o22a_1 _06343_ (.A1(\tms1x00.O_pla_ands[30][9] ),
    .A2(net611),
    .B1(net776),
    .B2(\tms1x00.O_pla_ands[31][9] ),
    .X(_02828_));
 sky130_fd_sc_hd__o221a_1 _06344_ (.A1(\tms1x00.O_pla_ands[29][9] ),
    .A2(net884),
    .B1(net803),
    .B2(\tms1x00.O_pla_ands[28][9] ),
    .C1(net992),
    .X(_02829_));
 sky130_fd_sc_hd__o22a_1 _06345_ (.A1(\tms1x00.O_pla_ands[27][9] ),
    .A2(net855),
    .B1(net722),
    .B2(\tms1x00.O_pla_ands[26][9] ),
    .X(_02830_));
 sky130_fd_sc_hd__o211a_1 _06346_ (.A1(\tms1x00.O_pla_ands[24][9] ),
    .A2(net830),
    .B1(_02829_),
    .C1(_02830_),
    .X(_02831_));
 sky130_fd_sc_hd__o211a_1 _06347_ (.A1(\tms1x00.O_pla_ands[25][9] ),
    .A2(net748),
    .B1(_02828_),
    .C1(_02831_),
    .X(_02832_));
 sky130_fd_sc_hd__o22a_1 _06348_ (.A1(\tms1x00.O_pla_ands[22][9] ),
    .A2(net610),
    .B1(net776),
    .B2(\tms1x00.O_pla_ands[23][9] ),
    .X(_02833_));
 sky130_fd_sc_hd__o221a_1 _06349_ (.A1(\tms1x00.O_pla_ands[16][9] ),
    .A2(net835),
    .B1(net753),
    .B2(\tms1x00.O_pla_ands[17][9] ),
    .C1(net914),
    .X(_02834_));
 sky130_fd_sc_hd__o22a_1 _06350_ (.A1(\tms1x00.O_pla_ands[19][9] ),
    .A2(net858),
    .B1(net724),
    .B2(\tms1x00.O_pla_ands[18][9] ),
    .X(_02835_));
 sky130_fd_sc_hd__o211a_1 _06351_ (.A1(\tms1x00.O_pla_ands[20][9] ),
    .A2(net805),
    .B1(_02834_),
    .C1(_02835_),
    .X(_02836_));
 sky130_fd_sc_hd__o211a_1 _06352_ (.A1(\tms1x00.O_pla_ands[21][9] ),
    .A2(net885),
    .B1(_02833_),
    .C1(_02836_),
    .X(_02837_));
 sky130_fd_sc_hd__or3_4 _06353_ (.A(net925),
    .B(_02832_),
    .C(_02837_),
    .X(_02838_));
 sky130_fd_sc_hd__o22a_1 _06354_ (.A1(\tms1x00.O_pla_ands[13][9] ),
    .A2(net899),
    .B1(net735),
    .B2(\tms1x00.O_pla_ands[10][9] ),
    .X(_02839_));
 sky130_fd_sc_hd__o22a_1 _06355_ (.A1(\tms1x00.O_pla_ands[8][9] ),
    .A2(net843),
    .B1(net790),
    .B2(\tms1x00.O_pla_ands[15][9] ),
    .X(_02840_));
 sky130_fd_sc_hd__o221a_1 _06356_ (.A1(\tms1x00.O_pla_ands[14][9] ),
    .A2(net624),
    .B1(net871),
    .B2(\tms1x00.O_pla_ands[11][9] ),
    .C1(_02840_),
    .X(_02841_));
 sky130_fd_sc_hd__o211a_1 _06357_ (.A1(\tms1x00.O_pla_ands[12][9] ),
    .A2(net816),
    .B1(_02841_),
    .C1(net1000),
    .X(_02842_));
 sky130_fd_sc_hd__o211a_2 _06358_ (.A1(\tms1x00.O_pla_ands[9][9] ),
    .A2(net763),
    .B1(_02839_),
    .C1(_02842_),
    .X(_02843_));
 sky130_fd_sc_hd__o22a_1 _06359_ (.A1(\tms1x00.O_pla_ands[6][9] ),
    .A2(net622),
    .B1(net813),
    .B2(\tms1x00.O_pla_ands[4][9] ),
    .X(_02844_));
 sky130_fd_sc_hd__o22a_1 _06360_ (.A1(\tms1x00.O_pla_ands[5][9] ),
    .A2(net896),
    .B1(net845),
    .B2(\tms1x00.O_pla_ands[0][9] ),
    .X(_02845_));
 sky130_fd_sc_hd__o221a_1 _06361_ (.A1(\tms1x00.O_pla_ands[1][9] ),
    .A2(net765),
    .B1(net733),
    .B2(\tms1x00.O_pla_ands[2][9] ),
    .C1(_02845_),
    .X(_02846_));
 sky130_fd_sc_hd__o211a_1 _06362_ (.A1(\tms1x00.O_pla_ands[3][9] ),
    .A2(net868),
    .B1(_02846_),
    .C1(net921),
    .X(_02847_));
 sky130_fd_sc_hd__o211a_1 _06363_ (.A1(\tms1x00.O_pla_ands[7][9] ),
    .A2(net788),
    .B1(_02844_),
    .C1(_02847_),
    .X(_02848_));
 sky130_fd_sc_hd__or3_2 _06364_ (.A(net988),
    .B(_02843_),
    .C(_02848_),
    .X(_02849_));
 sky130_fd_sc_hd__or2_1 _06365_ (.A(\tms1x00.ins_pla_ors[0][9] ),
    .B(net841),
    .X(_02850_));
 sky130_fd_sc_hd__o22a_1 _06366_ (.A1(\tms1x00.ins_pla_ors[3][9] ),
    .A2(net866),
    .B1(net787),
    .B2(\tms1x00.ins_pla_ors[7][9] ),
    .X(_02851_));
 sky130_fd_sc_hd__o22a_1 _06367_ (.A1(\tms1x00.ins_pla_ors[5][9] ),
    .A2(net892),
    .B1(net760),
    .B2(\tms1x00.ins_pla_ors[1][9] ),
    .X(_02852_));
 sky130_fd_sc_hd__o221a_1 _06368_ (.A1(\tms1x00.ins_pla_ors[6][9] ),
    .A2(net620),
    .B1(net731),
    .B2(\tms1x00.ins_pla_ors[2][9] ),
    .C1(_02852_),
    .X(_02853_));
 sky130_fd_sc_hd__o211a_1 _06369_ (.A1(\tms1x00.ins_pla_ors[4][9] ),
    .A2(net810),
    .B1(_02853_),
    .C1(net919),
    .X(_02854_));
 sky130_fd_sc_hd__o22a_1 _06370_ (.A1(\tms1x00.ins_pla_ors[13][9] ),
    .A2(net881),
    .B1(net718),
    .B2(\tms1x00.ins_pla_ors[10][9] ),
    .X(_02855_));
 sky130_fd_sc_hd__o22a_1 _06371_ (.A1(\tms1x00.ins_pla_ors[11][9] ),
    .A2(net853),
    .B1(net799),
    .B2(\tms1x00.ins_pla_ors[12][9] ),
    .X(_02856_));
 sky130_fd_sc_hd__o221a_1 _06372_ (.A1(\tms1x00.ins_pla_ors[8][9] ),
    .A2(net827),
    .B1(net745),
    .B2(\tms1x00.ins_pla_ors[9][9] ),
    .C1(net990),
    .X(_02857_));
 sky130_fd_sc_hd__o221a_1 _06373_ (.A1(\tms1x00.ins_pla_ors[14][9] ),
    .A2(net605),
    .B1(net773),
    .B2(\tms1x00.ins_pla_ors[15][9] ),
    .C1(_02855_),
    .X(_02858_));
 sky130_fd_sc_hd__and3_4 _06374_ (.A(_02856_),
    .B(_02857_),
    .C(_02858_),
    .X(_02859_));
 sky130_fd_sc_hd__a31o_4 _06375_ (.A1(_02850_),
    .A2(_02851_),
    .A3(_02854_),
    .B1(_02859_),
    .X(_02860_));
 sky130_fd_sc_hd__o22a_1 _06376_ (.A1(\tms1x00.O_pla_ors[0][9] ),
    .A2(net844),
    .B1(net764),
    .B2(\tms1x00.O_pla_ors[1][9] ),
    .X(_02861_));
 sky130_fd_sc_hd__o22a_1 _06377_ (.A1(\tms1x00.O_pla_ors[4][9] ),
    .A2(net818),
    .B1(net792),
    .B2(\tms1x00.O_pla_ors[7][9] ),
    .X(_02862_));
 sky130_fd_sc_hd__o221a_1 _06378_ (.A1(\tms1x00.O_pla_ors[6][9] ),
    .A2(net625),
    .B1(net737),
    .B2(\tms1x00.O_pla_ors[2][9] ),
    .C1(_02862_),
    .X(_02863_));
 sky130_fd_sc_hd__o211a_1 _06379_ (.A1(\tms1x00.O_pla_ors[3][9] ),
    .A2(net872),
    .B1(_02283_),
    .C1(_02863_),
    .X(_02864_));
 sky130_fd_sc_hd__o211a_2 _06380_ (.A1(\tms1x00.O_pla_ors[5][9] ),
    .A2(net900),
    .B1(_02861_),
    .C1(_02864_),
    .X(_02865_));
 sky130_fd_sc_hd__a211o_2 _06381_ (.A1(net601),
    .A2(_02860_),
    .B1(_02865_),
    .C1(net713),
    .X(_02866_));
 sky130_fd_sc_hd__a31o_1 _06382_ (.A1(_02774_),
    .A2(_02838_),
    .A3(_02849_),
    .B1(_02866_),
    .X(_02867_));
 sky130_fd_sc_hd__o22a_1 _06383_ (.A1(\tms1x00.ins_pla_ands[0][9] ),
    .A2(net832),
    .B1(net779),
    .B2(\tms1x00.ins_pla_ands[7][9] ),
    .X(_02868_));
 sky130_fd_sc_hd__o221a_1 _06384_ (.A1(\tms1x00.ins_pla_ands[5][9] ),
    .A2(net894),
    .B1(net812),
    .B2(\tms1x00.ins_pla_ands[4][9] ),
    .C1(net921),
    .X(_02869_));
 sky130_fd_sc_hd__o22a_1 _06385_ (.A1(\tms1x00.ins_pla_ands[3][9] ),
    .A2(net859),
    .B1(net725),
    .B2(\tms1x00.ins_pla_ands[2][9] ),
    .X(_02870_));
 sky130_fd_sc_hd__o221a_1 _06386_ (.A1(\tms1x00.ins_pla_ands[6][9] ),
    .A2(net613),
    .B1(net750),
    .B2(\tms1x00.ins_pla_ands[1][9] ),
    .C1(_02870_),
    .X(_02871_));
 sky130_fd_sc_hd__and3_2 _06387_ (.A(_02868_),
    .B(_02869_),
    .C(_02871_),
    .X(_02872_));
 sky130_fd_sc_hd__or2_1 _06388_ (.A(\tms1x00.ins_pla_ands[12][9] ),
    .B(net801),
    .X(_02873_));
 sky130_fd_sc_hd__o22a_1 _06389_ (.A1(\tms1x00.ins_pla_ands[11][9] ),
    .A2(net854),
    .B1(net747),
    .B2(\tms1x00.ins_pla_ands[9][9] ),
    .X(_02874_));
 sky130_fd_sc_hd__o22a_1 _06390_ (.A1(\tms1x00.ins_pla_ands[13][9] ),
    .A2(net883),
    .B1(net774),
    .B2(\tms1x00.ins_pla_ands[15][9] ),
    .X(_02875_));
 sky130_fd_sc_hd__o221a_1 _06391_ (.A1(\tms1x00.ins_pla_ands[14][9] ),
    .A2(net608),
    .B1(net829),
    .B2(\tms1x00.ins_pla_ands[8][9] ),
    .C1(_02875_),
    .X(_02876_));
 sky130_fd_sc_hd__o211a_1 _06392_ (.A1(\tms1x00.ins_pla_ands[10][9] ),
    .A2(net720),
    .B1(_02876_),
    .C1(net993),
    .X(_02877_));
 sky130_fd_sc_hd__o22a_1 _06393_ (.A1(\tms1x00.ins_pla_ands[21][9] ),
    .A2(net878),
    .B1(net797),
    .B2(\tms1x00.ins_pla_ands[20][9] ),
    .X(_02878_));
 sky130_fd_sc_hd__o22a_1 _06394_ (.A1(\tms1x00.ins_pla_ands[23][9] ),
    .A2(net770),
    .B1(net744),
    .B2(\tms1x00.ins_pla_ands[17][9] ),
    .X(_02879_));
 sky130_fd_sc_hd__o221a_1 _06395_ (.A1(\tms1x00.ins_pla_ands[22][9] ),
    .A2(net604),
    .B1(net825),
    .B2(\tms1x00.ins_pla_ands[16][9] ),
    .C1(_02879_),
    .X(_02880_));
 sky130_fd_sc_hd__o211a_1 _06396_ (.A1(\tms1x00.ins_pla_ands[18][9] ),
    .A2(net715),
    .B1(_02880_),
    .C1(net912),
    .X(_02881_));
 sky130_fd_sc_hd__o211a_1 _06397_ (.A1(\tms1x00.ins_pla_ands[19][9] ),
    .A2(net851),
    .B1(_02878_),
    .C1(_02881_),
    .X(_02882_));
 sky130_fd_sc_hd__o22a_1 _06398_ (.A1(\tms1x00.ins_pla_ands[30][9] ),
    .A2(net602),
    .B1(net769),
    .B2(\tms1x00.ins_pla_ands[31][9] ),
    .X(_02883_));
 sky130_fd_sc_hd__o221a_1 _06399_ (.A1(\tms1x00.ins_pla_ands[29][9] ),
    .A2(net879),
    .B1(net798),
    .B2(\tms1x00.ins_pla_ands[28][9] ),
    .C1(net990),
    .X(_02884_));
 sky130_fd_sc_hd__o22a_1 _06400_ (.A1(\tms1x00.ins_pla_ands[27][9] ),
    .A2(net852),
    .B1(net717),
    .B2(\tms1x00.ins_pla_ands[26][9] ),
    .X(_02885_));
 sky130_fd_sc_hd__o211a_1 _06401_ (.A1(\tms1x00.ins_pla_ands[24][9] ),
    .A2(net823),
    .B1(_02884_),
    .C1(_02885_),
    .X(_02886_));
 sky130_fd_sc_hd__o211a_2 _06402_ (.A1(\tms1x00.ins_pla_ands[25][9] ),
    .A2(net742),
    .B1(_02883_),
    .C1(_02886_),
    .X(_02887_));
 sky130_fd_sc_hd__o21a_1 _06403_ (.A1(_02882_),
    .A2(_02887_),
    .B1(net989),
    .X(_02888_));
 sky130_fd_sc_hd__a31o_1 _06404_ (.A1(_02873_),
    .A2(_02874_),
    .A3(_02877_),
    .B1(_02872_),
    .X(_02889_));
 sky130_fd_sc_hd__a211o_4 _06405_ (.A1(net925),
    .A2(_02889_),
    .B1(_02888_),
    .C1(net711),
    .X(_02890_));
 sky130_fd_sc_hd__and2_1 _06406_ (.A(net907),
    .B(\wbs_o_buff[9] ),
    .X(_02891_));
 sky130_fd_sc_hd__a21o_1 _06407_ (.A1(_02867_),
    .A2(_02890_),
    .B1(net587),
    .X(_02892_));
 sky130_fd_sc_hd__o211a_1 _06408_ (.A1(net589),
    .A2(_02891_),
    .B1(_02892_),
    .C1(net629),
    .X(_02893_));
 sky130_fd_sc_hd__a221o_1 _06409_ (.A1(net129),
    .A2(net580),
    .B1(_02891_),
    .B2(net584),
    .C1(_02893_),
    .X(_00036_));
 sky130_fd_sc_hd__o22a_1 _06410_ (.A1(\tms1x00.ins_pla_ands[6][10] ),
    .A2(net613),
    .B1(net780),
    .B2(\tms1x00.ins_pla_ands[7][10] ),
    .X(_02894_));
 sky130_fd_sc_hd__o22a_1 _06411_ (.A1(\tms1x00.ins_pla_ands[3][10] ),
    .A2(net870),
    .B1(net732),
    .B2(\tms1x00.ins_pla_ands[2][10] ),
    .X(_02895_));
 sky130_fd_sc_hd__o221a_1 _06412_ (.A1(\tms1x00.ins_pla_ands[5][10] ),
    .A2(net894),
    .B1(net815),
    .B2(\tms1x00.ins_pla_ands[4][10] ),
    .C1(net921),
    .X(_02896_));
 sky130_fd_sc_hd__o211a_1 _06413_ (.A1(\tms1x00.ins_pla_ands[0][10] ),
    .A2(net845),
    .B1(_02895_),
    .C1(_02896_),
    .X(_02897_));
 sky130_fd_sc_hd__o211a_1 _06414_ (.A1(\tms1x00.ins_pla_ands[1][10] ),
    .A2(net750),
    .B1(_02894_),
    .C1(_02897_),
    .X(_02898_));
 sky130_fd_sc_hd__o22a_1 _06415_ (.A1(\tms1x00.ins_pla_ands[14][10] ),
    .A2(net609),
    .B1(net774),
    .B2(\tms1x00.ins_pla_ands[15][10] ),
    .X(_02899_));
 sky130_fd_sc_hd__o221a_1 _06416_ (.A1(\tms1x00.ins_pla_ands[8][10] ),
    .A2(net832),
    .B1(net751),
    .B2(\tms1x00.ins_pla_ands[9][10] ),
    .C1(net994),
    .X(_02900_));
 sky130_fd_sc_hd__o22a_1 _06417_ (.A1(\tms1x00.ins_pla_ands[11][10] ),
    .A2(net857),
    .B1(net721),
    .B2(\tms1x00.ins_pla_ands[10][10] ),
    .X(_02901_));
 sky130_fd_sc_hd__o211a_1 _06418_ (.A1(\tms1x00.ins_pla_ands[13][10] ),
    .A2(net882),
    .B1(_02900_),
    .C1(_02901_),
    .X(_02902_));
 sky130_fd_sc_hd__o211a_2 _06419_ (.A1(\tms1x00.ins_pla_ands[12][10] ),
    .A2(net801),
    .B1(_02899_),
    .C1(_02902_),
    .X(_02903_));
 sky130_fd_sc_hd__or3_2 _06420_ (.A(net988),
    .B(_02898_),
    .C(_02903_),
    .X(_02904_));
 sky130_fd_sc_hd__o22a_2 _06421_ (.A1(\tms1x00.ins_pla_ands[30][10] ),
    .A2(net602),
    .B1(net742),
    .B2(\tms1x00.ins_pla_ands[25][10] ),
    .X(_02905_));
 sky130_fd_sc_hd__o22a_1 _06422_ (.A1(\tms1x00.ins_pla_ands[27][10] ),
    .A2(net850),
    .B1(net824),
    .B2(\tms1x00.ins_pla_ands[24][10] ),
    .X(_02906_));
 sky130_fd_sc_hd__o221a_1 _06423_ (.A1(\tms1x00.ins_pla_ands[29][10] ),
    .A2(net880),
    .B1(net769),
    .B2(\tms1x00.ins_pla_ands[31][10] ),
    .C1(_02906_),
    .X(_02907_));
 sky130_fd_sc_hd__o211a_1 _06424_ (.A1(\tms1x00.ins_pla_ands[28][10] ),
    .A2(net798),
    .B1(_02907_),
    .C1(net991),
    .X(_02908_));
 sky130_fd_sc_hd__o211a_1 _06425_ (.A1(\tms1x00.ins_pla_ands[26][10] ),
    .A2(net714),
    .B1(_02905_),
    .C1(_02908_),
    .X(_02909_));
 sky130_fd_sc_hd__o22a_1 _06426_ (.A1(\tms1x00.ins_pla_ands[17][10] ),
    .A2(net744),
    .B1(net715),
    .B2(\tms1x00.ins_pla_ands[18][10] ),
    .X(_02910_));
 sky130_fd_sc_hd__o22a_1 _06427_ (.A1(\tms1x00.ins_pla_ands[16][10] ),
    .A2(net825),
    .B1(net770),
    .B2(\tms1x00.ins_pla_ands[23][10] ),
    .X(_02911_));
 sky130_fd_sc_hd__o221a_1 _06428_ (.A1(\tms1x00.ins_pla_ands[21][10] ),
    .A2(net878),
    .B1(net800),
    .B2(\tms1x00.ins_pla_ands[20][10] ),
    .C1(_02911_),
    .X(_02912_));
 sky130_fd_sc_hd__o211a_1 _06429_ (.A1(\tms1x00.ins_pla_ands[19][10] ),
    .A2(net851),
    .B1(_02912_),
    .C1(net912),
    .X(_02913_));
 sky130_fd_sc_hd__o211a_1 _06430_ (.A1(\tms1x00.ins_pla_ands[22][10] ),
    .A2(net607),
    .B1(_02910_),
    .C1(_02913_),
    .X(_02914_));
 sky130_fd_sc_hd__or3_4 _06431_ (.A(net924),
    .B(_02909_),
    .C(_02914_),
    .X(_02915_));
 sky130_fd_sc_hd__a22o_1 _06432_ (.A1(\tms1x00.ins_pla_ors[3][10] ),
    .A2(net875),
    .B1(net848),
    .B2(\tms1x00.ins_pla_ors[0][10] ),
    .X(_02916_));
 sky130_fd_sc_hd__a22o_1 _06433_ (.A1(\tms1x00.ins_pla_ors[4][10] ),
    .A2(net821),
    .B1(net794),
    .B2(\tms1x00.ins_pla_ors[7][10] ),
    .X(_02917_));
 sky130_fd_sc_hd__a221o_1 _06434_ (.A1(\tms1x00.ins_pla_ors[6][10] ),
    .A2(net627),
    .B1(net767),
    .B2(\tms1x00.ins_pla_ors[1][10] ),
    .C1(_02917_),
    .X(_02918_));
 sky130_fd_sc_hd__a211o_1 _06435_ (.A1(\tms1x00.ins_pla_ors[2][10] ),
    .A2(net740),
    .B1(_02918_),
    .C1(net998),
    .X(_02919_));
 sky130_fd_sc_hd__a211o_4 _06436_ (.A1(\tms1x00.ins_pla_ors[5][10] ),
    .A2(net903),
    .B1(_02916_),
    .C1(_02919_),
    .X(_02920_));
 sky130_fd_sc_hd__a22o_1 _06437_ (.A1(\tms1x00.ins_pla_ors[11][10] ),
    .A2(net874),
    .B1(net739),
    .B2(\tms1x00.ins_pla_ors[10][10] ),
    .X(_02921_));
 sky130_fd_sc_hd__a22o_1 _06438_ (.A1(\tms1x00.ins_pla_ors[14][10] ),
    .A2(net628),
    .B1(net795),
    .B2(\tms1x00.ins_pla_ors[15][10] ),
    .X(_02922_));
 sky130_fd_sc_hd__a221o_1 _06439_ (.A1(\tms1x00.ins_pla_ors[13][10] ),
    .A2(net902),
    .B1(net820),
    .B2(\tms1x00.ins_pla_ors[12][10] ),
    .C1(net920),
    .X(_02923_));
 sky130_fd_sc_hd__a211o_1 _06440_ (.A1(\tms1x00.ins_pla_ors[8][10] ),
    .A2(net847),
    .B1(_02921_),
    .C1(_02923_),
    .X(_02924_));
 sky130_fd_sc_hd__a211o_1 _06441_ (.A1(\tms1x00.ins_pla_ors[9][10] ),
    .A2(net766),
    .B1(_02922_),
    .C1(_02924_),
    .X(_02925_));
 sky130_fd_sc_hd__a21o_1 _06442_ (.A1(_02920_),
    .A2(_02925_),
    .B1(net984),
    .X(_02926_));
 sky130_fd_sc_hd__a22o_1 _06443_ (.A1(\tms1x00.O_pla_ors[6][10] ),
    .A2(net627),
    .B1(net794),
    .B2(\tms1x00.O_pla_ors[7][10] ),
    .X(_02927_));
 sky130_fd_sc_hd__a221o_1 _06444_ (.A1(\tms1x00.O_pla_ors[0][10] ),
    .A2(net848),
    .B1(net767),
    .B2(\tms1x00.O_pla_ors[1][10] ),
    .C1(_01637_),
    .X(_02928_));
 sky130_fd_sc_hd__a22o_1 _06445_ (.A1(\tms1x00.O_pla_ors[3][10] ),
    .A2(net875),
    .B1(net740),
    .B2(\tms1x00.O_pla_ors[2][10] ),
    .X(_02929_));
 sky130_fd_sc_hd__a211o_1 _06446_ (.A1(\tms1x00.O_pla_ors[5][10] ),
    .A2(net903),
    .B1(_02928_),
    .C1(_02929_),
    .X(_02930_));
 sky130_fd_sc_hd__a211o_4 _06447_ (.A1(\tms1x00.O_pla_ors[4][10] ),
    .A2(net821),
    .B1(_02927_),
    .C1(_02930_),
    .X(_02931_));
 sky130_fd_sc_hd__a31o_1 _06448_ (.A1(net985),
    .A2(_02926_),
    .A3(_02931_),
    .B1(net587),
    .X(_02932_));
 sky130_fd_sc_hd__a31o_1 _06449_ (.A1(net713),
    .A2(_02904_),
    .A3(_02915_),
    .B1(_02932_),
    .X(_02933_));
 sky130_fd_sc_hd__and2_1 _06450_ (.A(net906),
    .B(\wbs_o_buff[10] ),
    .X(_02934_));
 sky130_fd_sc_hd__o211a_1 _06451_ (.A1(net589),
    .A2(_02934_),
    .B1(_02933_),
    .C1(net629),
    .X(_02935_));
 sky130_fd_sc_hd__a221o_1 _06452_ (.A1(net130),
    .A2(net580),
    .B1(_02934_),
    .B2(net585),
    .C1(_02935_),
    .X(_00006_));
 sky130_fd_sc_hd__o22a_1 _06453_ (.A1(\tms1x00.ins_pla_ands[0][11] ),
    .A2(net833),
    .B1(net779),
    .B2(\tms1x00.ins_pla_ands[7][11] ),
    .X(_02936_));
 sky130_fd_sc_hd__o221a_2 _06454_ (.A1(\tms1x00.ins_pla_ands[5][11] ),
    .A2(net894),
    .B1(net812),
    .B2(\tms1x00.ins_pla_ands[4][11] ),
    .C1(net921),
    .X(_02937_));
 sky130_fd_sc_hd__o22a_1 _06455_ (.A1(\tms1x00.ins_pla_ands[3][11] ),
    .A2(net870),
    .B1(net732),
    .B2(\tms1x00.ins_pla_ands[2][11] ),
    .X(_02938_));
 sky130_fd_sc_hd__o221a_1 _06456_ (.A1(\tms1x00.ins_pla_ands[6][11] ),
    .A2(net613),
    .B1(net750),
    .B2(\tms1x00.ins_pla_ands[1][11] ),
    .C1(_02938_),
    .X(_02939_));
 sky130_fd_sc_hd__o22a_1 _06457_ (.A1(\tms1x00.ins_pla_ands[14][11] ),
    .A2(net608),
    .B1(net774),
    .B2(\tms1x00.ins_pla_ands[15][11] ),
    .X(_02940_));
 sky130_fd_sc_hd__o221a_1 _06458_ (.A1(\tms1x00.ins_pla_ands[8][11] ),
    .A2(net832),
    .B1(net751),
    .B2(\tms1x00.ins_pla_ands[9][11] ),
    .C1(net994),
    .X(_02941_));
 sky130_fd_sc_hd__o22a_1 _06459_ (.A1(\tms1x00.ins_pla_ands[11][11] ),
    .A2(net857),
    .B1(net721),
    .B2(\tms1x00.ins_pla_ands[10][11] ),
    .X(_02942_));
 sky130_fd_sc_hd__o211a_1 _06460_ (.A1(\tms1x00.ins_pla_ands[13][11] ),
    .A2(net882),
    .B1(_02941_),
    .C1(_02942_),
    .X(_02943_));
 sky130_fd_sc_hd__o211a_2 _06461_ (.A1(\tms1x00.ins_pla_ands[12][11] ),
    .A2(net801),
    .B1(_02940_),
    .C1(_02943_),
    .X(_02944_));
 sky130_fd_sc_hd__a31o_1 _06462_ (.A1(_02936_),
    .A2(_02937_),
    .A3(_02939_),
    .B1(net986),
    .X(_02945_));
 sky130_fd_sc_hd__o22a_1 _06463_ (.A1(\tms1x00.ins_pla_ands[27][11] ),
    .A2(net850),
    .B1(net714),
    .B2(\tms1x00.ins_pla_ands[26][11] ),
    .X(_02946_));
 sky130_fd_sc_hd__o22a_1 _06464_ (.A1(\tms1x00.ins_pla_ands[30][11] ),
    .A2(net602),
    .B1(net742),
    .B2(\tms1x00.ins_pla_ands[25][11] ),
    .X(_02947_));
 sky130_fd_sc_hd__o221a_1 _06465_ (.A1(\tms1x00.ins_pla_ands[29][11] ),
    .A2(net879),
    .B1(net798),
    .B2(\tms1x00.ins_pla_ands[28][11] ),
    .C1(net991),
    .X(_02948_));
 sky130_fd_sc_hd__o221a_1 _06466_ (.A1(\tms1x00.ins_pla_ands[24][11] ),
    .A2(net823),
    .B1(net771),
    .B2(\tms1x00.ins_pla_ands[31][11] ),
    .C1(_02948_),
    .X(_02949_));
 sky130_fd_sc_hd__and3_1 _06467_ (.A(_02946_),
    .B(_02947_),
    .C(_02949_),
    .X(_02950_));
 sky130_fd_sc_hd__or2_1 _06468_ (.A(\tms1x00.ins_pla_ands[21][11] ),
    .B(net878),
    .X(_02951_));
 sky130_fd_sc_hd__o221a_1 _06469_ (.A1(\tms1x00.ins_pla_ands[20][11] ),
    .A2(net800),
    .B1(net770),
    .B2(\tms1x00.ins_pla_ands[23][11] ),
    .C1(_02951_),
    .X(_02952_));
 sky130_fd_sc_hd__o22a_1 _06470_ (.A1(\tms1x00.ins_pla_ands[16][11] ),
    .A2(net826),
    .B1(net744),
    .B2(\tms1x00.ins_pla_ands[17][11] ),
    .X(_02953_));
 sky130_fd_sc_hd__o221a_1 _06471_ (.A1(\tms1x00.ins_pla_ands[22][11] ),
    .A2(net604),
    .B1(net715),
    .B2(\tms1x00.ins_pla_ands[18][11] ),
    .C1(_02953_),
    .X(_02954_));
 sky130_fd_sc_hd__o211a_1 _06472_ (.A1(\tms1x00.ins_pla_ands[19][11] ),
    .A2(net851),
    .B1(_02954_),
    .C1(net911),
    .X(_02955_));
 sky130_fd_sc_hd__a211o_2 _06473_ (.A1(_02952_),
    .A2(_02955_),
    .B1(net923),
    .C1(_02950_),
    .X(_02956_));
 sky130_fd_sc_hd__o211a_1 _06474_ (.A1(_02944_),
    .A2(_02945_),
    .B1(_02956_),
    .C1(net712),
    .X(_02957_));
 sky130_fd_sc_hd__a22o_1 _06475_ (.A1(\tms1x00.ins_pla_ors[3][11] ),
    .A2(net875),
    .B1(net767),
    .B2(\tms1x00.ins_pla_ors[1][11] ),
    .X(_02958_));
 sky130_fd_sc_hd__a22o_1 _06476_ (.A1(\tms1x00.ins_pla_ors[5][11] ),
    .A2(net903),
    .B1(net794),
    .B2(\tms1x00.ins_pla_ors[7][11] ),
    .X(_02959_));
 sky130_fd_sc_hd__a221o_2 _06477_ (.A1(\tms1x00.ins_pla_ors[6][11] ),
    .A2(net627),
    .B1(net740),
    .B2(\tms1x00.ins_pla_ors[2][11] ),
    .C1(_02959_),
    .X(_02960_));
 sky130_fd_sc_hd__a211o_1 _06478_ (.A1(\tms1x00.ins_pla_ors[0][11] ),
    .A2(net848),
    .B1(_02960_),
    .C1(net998),
    .X(_02961_));
 sky130_fd_sc_hd__a211o_2 _06479_ (.A1(\tms1x00.ins_pla_ors[4][11] ),
    .A2(net821),
    .B1(_02958_),
    .C1(_02961_),
    .X(_02962_));
 sky130_fd_sc_hd__a22o_1 _06480_ (.A1(\tms1x00.ins_pla_ors[14][11] ),
    .A2(net628),
    .B1(net795),
    .B2(\tms1x00.ins_pla_ors[15][11] ),
    .X(_02963_));
 sky130_fd_sc_hd__a221o_1 _06481_ (.A1(\tms1x00.ins_pla_ors[13][11] ),
    .A2(net902),
    .B1(net820),
    .B2(\tms1x00.ins_pla_ors[12][11] ),
    .C1(net913),
    .X(_02964_));
 sky130_fd_sc_hd__a22o_1 _06482_ (.A1(\tms1x00.ins_pla_ors[11][11] ),
    .A2(net874),
    .B1(net739),
    .B2(\tms1x00.ins_pla_ors[10][11] ),
    .X(_02965_));
 sky130_fd_sc_hd__a211o_1 _06483_ (.A1(\tms1x00.ins_pla_ors[8][11] ),
    .A2(net847),
    .B1(_02964_),
    .C1(_02965_),
    .X(_02966_));
 sky130_fd_sc_hd__a211o_2 _06484_ (.A1(\tms1x00.ins_pla_ors[9][11] ),
    .A2(net766),
    .B1(_02963_),
    .C1(_02966_),
    .X(_02967_));
 sky130_fd_sc_hd__a21o_1 _06485_ (.A1(_02962_),
    .A2(_02967_),
    .B1(net85),
    .X(_02968_));
 sky130_fd_sc_hd__a22o_1 _06486_ (.A1(\tms1x00.O_pla_ors[6][11] ),
    .A2(net627),
    .B1(net794),
    .B2(\tms1x00.O_pla_ors[7][11] ),
    .X(_02969_));
 sky130_fd_sc_hd__a221o_1 _06487_ (.A1(\tms1x00.O_pla_ors[0][11] ),
    .A2(net848),
    .B1(net767),
    .B2(\tms1x00.O_pla_ors[1][11] ),
    .C1(_01637_),
    .X(_02970_));
 sky130_fd_sc_hd__a22o_1 _06488_ (.A1(\tms1x00.O_pla_ors[3][11] ),
    .A2(net875),
    .B1(net741),
    .B2(\tms1x00.O_pla_ors[2][11] ),
    .X(_02971_));
 sky130_fd_sc_hd__a211o_1 _06489_ (.A1(\tms1x00.O_pla_ors[5][11] ),
    .A2(net903),
    .B1(_02970_),
    .C1(_02971_),
    .X(_02972_));
 sky130_fd_sc_hd__a211o_4 _06490_ (.A1(\tms1x00.O_pla_ors[4][11] ),
    .A2(net821),
    .B1(_02969_),
    .C1(_02972_),
    .X(_02973_));
 sky130_fd_sc_hd__a31o_1 _06491_ (.A1(net985),
    .A2(_02968_),
    .A3(_02973_),
    .B1(net587),
    .X(_02974_));
 sky130_fd_sc_hd__and2_1 _06492_ (.A(net907),
    .B(\wbs_o_buff[11] ),
    .X(_02975_));
 sky130_fd_sc_hd__or2_1 _06493_ (.A(net590),
    .B(_02975_),
    .X(_02976_));
 sky130_fd_sc_hd__o211a_1 _06494_ (.A1(_02957_),
    .A2(_02974_),
    .B1(_02976_),
    .C1(net629),
    .X(_02977_));
 sky130_fd_sc_hd__a221o_1 _06495_ (.A1(net131),
    .A2(net580),
    .B1(_02975_),
    .B2(net585),
    .C1(_02977_),
    .X(_00007_));
 sky130_fd_sc_hd__o22a_1 _06496_ (.A1(\tms1x00.ins_pla_ands[14][12] ),
    .A2(net608),
    .B1(net774),
    .B2(\tms1x00.ins_pla_ands[15][12] ),
    .X(_02978_));
 sky130_fd_sc_hd__o221a_2 _06497_ (.A1(\tms1x00.ins_pla_ands[8][12] ),
    .A2(net829),
    .B1(net747),
    .B2(\tms1x00.ins_pla_ands[9][12] ),
    .C1(net994),
    .X(_02979_));
 sky130_fd_sc_hd__o22a_1 _06498_ (.A1(\tms1x00.ins_pla_ands[11][12] ),
    .A2(net854),
    .B1(net720),
    .B2(\tms1x00.ins_pla_ands[10][12] ),
    .X(_02980_));
 sky130_fd_sc_hd__o211a_1 _06499_ (.A1(\tms1x00.ins_pla_ands[12][12] ),
    .A2(net802),
    .B1(_02979_),
    .C1(_02980_),
    .X(_02981_));
 sky130_fd_sc_hd__o211a_1 _06500_ (.A1(\tms1x00.ins_pla_ands[13][12] ),
    .A2(net883),
    .B1(_02978_),
    .C1(_02981_),
    .X(_02982_));
 sky130_fd_sc_hd__o22a_1 _06501_ (.A1(\tms1x00.ins_pla_ands[0][12] ),
    .A2(net833),
    .B1(net780),
    .B2(\tms1x00.ins_pla_ands[7][12] ),
    .X(_02983_));
 sky130_fd_sc_hd__o221a_2 _06502_ (.A1(\tms1x00.ins_pla_ands[5][12] ),
    .A2(net895),
    .B1(net812),
    .B2(\tms1x00.ins_pla_ands[4][12] ),
    .C1(net921),
    .X(_02984_));
 sky130_fd_sc_hd__o22a_1 _06503_ (.A1(\tms1x00.ins_pla_ands[3][12] ),
    .A2(net859),
    .B1(net725),
    .B2(\tms1x00.ins_pla_ands[2][12] ),
    .X(_02985_));
 sky130_fd_sc_hd__o221a_1 _06504_ (.A1(\tms1x00.ins_pla_ands[6][12] ),
    .A2(net613),
    .B1(net750),
    .B2(\tms1x00.ins_pla_ands[1][12] ),
    .C1(_02985_),
    .X(_02986_));
 sky130_fd_sc_hd__a31o_4 _06505_ (.A1(_02983_),
    .A2(_02984_),
    .A3(_02986_),
    .B1(net987),
    .X(_02987_));
 sky130_fd_sc_hd__o22a_1 _06506_ (.A1(\tms1x00.ins_pla_ands[20][12] ),
    .A2(net800),
    .B1(net715),
    .B2(\tms1x00.ins_pla_ands[18][12] ),
    .X(_02988_));
 sky130_fd_sc_hd__o22a_1 _06507_ (.A1(\tms1x00.ins_pla_ands[16][12] ),
    .A2(net825),
    .B1(net744),
    .B2(\tms1x00.ins_pla_ands[17][12] ),
    .X(_02989_));
 sky130_fd_sc_hd__o221a_1 _06508_ (.A1(\tms1x00.ins_pla_ands[22][12] ),
    .A2(net604),
    .B1(net851),
    .B2(\tms1x00.ins_pla_ands[19][12] ),
    .C1(_02989_),
    .X(_02990_));
 sky130_fd_sc_hd__o211a_1 _06509_ (.A1(\tms1x00.ins_pla_ands[21][12] ),
    .A2(net878),
    .B1(_02990_),
    .C1(net912),
    .X(_02991_));
 sky130_fd_sc_hd__o211a_1 _06510_ (.A1(\tms1x00.ins_pla_ands[23][12] ),
    .A2(net770),
    .B1(_02988_),
    .C1(_02991_),
    .X(_02992_));
 sky130_fd_sc_hd__o22a_2 _06511_ (.A1(\tms1x00.ins_pla_ands[27][12] ),
    .A2(net852),
    .B1(net717),
    .B2(\tms1x00.ins_pla_ands[26][12] ),
    .X(_02993_));
 sky130_fd_sc_hd__o221a_1 _06512_ (.A1(\tms1x00.ins_pla_ands[30][12] ),
    .A2(net602),
    .B1(net742),
    .B2(\tms1x00.ins_pla_ands[25][12] ),
    .C1(_02993_),
    .X(_02994_));
 sky130_fd_sc_hd__o221a_1 _06513_ (.A1(\tms1x00.ins_pla_ands[29][12] ),
    .A2(net877),
    .B1(net796),
    .B2(\tms1x00.ins_pla_ands[28][12] ),
    .C1(net990),
    .X(_02995_));
 sky130_fd_sc_hd__o221a_1 _06514_ (.A1(\tms1x00.ins_pla_ands[24][12] ),
    .A2(net824),
    .B1(net769),
    .B2(\tms1x00.ins_pla_ands[31][12] ),
    .C1(_02995_),
    .X(_02996_));
 sky130_fd_sc_hd__a21o_2 _06515_ (.A1(_02994_),
    .A2(_02996_),
    .B1(net923),
    .X(_02997_));
 sky130_fd_sc_hd__o22a_4 _06516_ (.A1(_02982_),
    .A2(_02987_),
    .B1(_02992_),
    .B2(_02997_),
    .X(_02998_));
 sky130_fd_sc_hd__a22o_1 _06517_ (.A1(\tms1x00.ins_pla_ors[3][12] ),
    .A2(net875),
    .B1(net848),
    .B2(\tms1x00.ins_pla_ors[0][12] ),
    .X(_02999_));
 sky130_fd_sc_hd__a22o_1 _06518_ (.A1(\tms1x00.ins_pla_ors[5][12] ),
    .A2(net903),
    .B1(net794),
    .B2(\tms1x00.ins_pla_ors[7][12] ),
    .X(_03000_));
 sky130_fd_sc_hd__a221o_1 _06519_ (.A1(\tms1x00.ins_pla_ors[6][12] ),
    .A2(net627),
    .B1(net740),
    .B2(\tms1x00.ins_pla_ors[2][12] ),
    .C1(_03000_),
    .X(_03001_));
 sky130_fd_sc_hd__a211o_1 _06520_ (.A1(\tms1x00.ins_pla_ors[1][12] ),
    .A2(net767),
    .B1(_03001_),
    .C1(net998),
    .X(_03002_));
 sky130_fd_sc_hd__a211o_2 _06521_ (.A1(\tms1x00.ins_pla_ors[4][12] ),
    .A2(net821),
    .B1(_02999_),
    .C1(_03002_),
    .X(_03003_));
 sky130_fd_sc_hd__a22o_1 _06522_ (.A1(\tms1x00.ins_pla_ors[11][12] ),
    .A2(net874),
    .B1(net739),
    .B2(\tms1x00.ins_pla_ors[10][12] ),
    .X(_03004_));
 sky130_fd_sc_hd__a22o_1 _06523_ (.A1(\tms1x00.ins_pla_ors[14][12] ),
    .A2(net628),
    .B1(net795),
    .B2(\tms1x00.ins_pla_ors[15][12] ),
    .X(_03005_));
 sky130_fd_sc_hd__a221o_1 _06524_ (.A1(\tms1x00.ins_pla_ors[13][12] ),
    .A2(net902),
    .B1(net820),
    .B2(\tms1x00.ins_pla_ors[12][12] ),
    .C1(net913),
    .X(_03006_));
 sky130_fd_sc_hd__a211o_1 _06525_ (.A1(\tms1x00.ins_pla_ors[9][12] ),
    .A2(net766),
    .B1(_03004_),
    .C1(_03006_),
    .X(_03007_));
 sky130_fd_sc_hd__a211o_1 _06526_ (.A1(\tms1x00.ins_pla_ors[8][12] ),
    .A2(net847),
    .B1(_03005_),
    .C1(_03007_),
    .X(_03008_));
 sky130_fd_sc_hd__a21o_1 _06527_ (.A1(_03003_),
    .A2(_03008_),
    .B1(net984),
    .X(_03009_));
 sky130_fd_sc_hd__a22o_1 _06528_ (.A1(\tms1x00.O_pla_ors[6][12] ),
    .A2(net627),
    .B1(net794),
    .B2(\tms1x00.O_pla_ors[7][12] ),
    .X(_03010_));
 sky130_fd_sc_hd__a221o_1 _06529_ (.A1(\tms1x00.O_pla_ors[0][12] ),
    .A2(net848),
    .B1(net767),
    .B2(\tms1x00.O_pla_ors[1][12] ),
    .C1(_01637_),
    .X(_03011_));
 sky130_fd_sc_hd__a22o_1 _06530_ (.A1(\tms1x00.O_pla_ors[3][12] ),
    .A2(net875),
    .B1(net740),
    .B2(\tms1x00.O_pla_ors[2][12] ),
    .X(_03012_));
 sky130_fd_sc_hd__a211o_1 _06531_ (.A1(\tms1x00.O_pla_ors[5][12] ),
    .A2(net903),
    .B1(_03011_),
    .C1(_03012_),
    .X(_03013_));
 sky130_fd_sc_hd__a211o_2 _06532_ (.A1(\tms1x00.O_pla_ors[4][12] ),
    .A2(net821),
    .B1(_03010_),
    .C1(_03013_),
    .X(_03014_));
 sky130_fd_sc_hd__a32o_1 _06533_ (.A1(net985),
    .A2(_03009_),
    .A3(_03014_),
    .B1(net713),
    .B2(_02998_),
    .X(_03015_));
 sky130_fd_sc_hd__and2_1 _06534_ (.A(net907),
    .B(\wbs_o_buff[12] ),
    .X(_03016_));
 sky130_fd_sc_hd__or2_1 _06535_ (.A(net589),
    .B(_03016_),
    .X(_03017_));
 sky130_fd_sc_hd__o211a_1 _06536_ (.A1(net587),
    .A2(_03015_),
    .B1(_03017_),
    .C1(net629),
    .X(_03018_));
 sky130_fd_sc_hd__a221o_1 _06537_ (.A1(net132),
    .A2(net579),
    .B1(_03016_),
    .B2(net585),
    .C1(_03018_),
    .X(_00008_));
 sky130_fd_sc_hd__o22a_1 _06538_ (.A1(\tms1x00.ins_pla_ands[0][13] ),
    .A2(net833),
    .B1(net780),
    .B2(\tms1x00.ins_pla_ands[7][13] ),
    .X(_03019_));
 sky130_fd_sc_hd__o221a_2 _06539_ (.A1(\tms1x00.ins_pla_ands[5][13] ),
    .A2(net895),
    .B1(net812),
    .B2(\tms1x00.ins_pla_ands[4][13] ),
    .C1(net921),
    .X(_03020_));
 sky130_fd_sc_hd__o22a_1 _06540_ (.A1(\tms1x00.ins_pla_ands[3][13] ),
    .A2(net859),
    .B1(net725),
    .B2(\tms1x00.ins_pla_ands[2][13] ),
    .X(_03021_));
 sky130_fd_sc_hd__o221a_1 _06541_ (.A1(\tms1x00.ins_pla_ands[6][13] ),
    .A2(net613),
    .B1(net751),
    .B2(\tms1x00.ins_pla_ands[1][13] ),
    .C1(_03021_),
    .X(_03022_));
 sky130_fd_sc_hd__o22a_1 _06542_ (.A1(\tms1x00.ins_pla_ands[14][13] ),
    .A2(net608),
    .B1(net774),
    .B2(\tms1x00.ins_pla_ands[15][13] ),
    .X(_03023_));
 sky130_fd_sc_hd__o221a_2 _06543_ (.A1(\tms1x00.ins_pla_ands[8][13] ),
    .A2(net829),
    .B1(net747),
    .B2(\tms1x00.ins_pla_ands[9][13] ),
    .C1(net994),
    .X(_03024_));
 sky130_fd_sc_hd__o22a_1 _06544_ (.A1(\tms1x00.ins_pla_ands[11][13] ),
    .A2(net854),
    .B1(net720),
    .B2(\tms1x00.ins_pla_ands[10][13] ),
    .X(_03025_));
 sky130_fd_sc_hd__o211a_1 _06545_ (.A1(\tms1x00.ins_pla_ands[13][13] ),
    .A2(net883),
    .B1(_03024_),
    .C1(_03025_),
    .X(_03026_));
 sky130_fd_sc_hd__o211a_2 _06546_ (.A1(\tms1x00.ins_pla_ands[12][13] ),
    .A2(net802),
    .B1(_03023_),
    .C1(_03026_),
    .X(_03027_));
 sky130_fd_sc_hd__a31o_2 _06547_ (.A1(_03019_),
    .A2(_03020_),
    .A3(_03022_),
    .B1(net987),
    .X(_03028_));
 sky130_fd_sc_hd__o22a_1 _06548_ (.A1(\tms1x00.ins_pla_ands[27][13] ),
    .A2(net852),
    .B1(net717),
    .B2(\tms1x00.ins_pla_ands[26][13] ),
    .X(_03029_));
 sky130_fd_sc_hd__o22a_1 _06549_ (.A1(\tms1x00.ins_pla_ands[30][13] ),
    .A2(net602),
    .B1(net742),
    .B2(\tms1x00.ins_pla_ands[25][13] ),
    .X(_03030_));
 sky130_fd_sc_hd__o221a_1 _06550_ (.A1(\tms1x00.ins_pla_ands[29][13] ),
    .A2(net879),
    .B1(net798),
    .B2(\tms1x00.ins_pla_ands[28][13] ),
    .C1(net990),
    .X(_03031_));
 sky130_fd_sc_hd__o221a_1 _06551_ (.A1(\tms1x00.ins_pla_ands[24][13] ),
    .A2(net823),
    .B1(net771),
    .B2(\tms1x00.ins_pla_ands[31][13] ),
    .C1(_03031_),
    .X(_03032_));
 sky130_fd_sc_hd__and3_1 _06552_ (.A(_03029_),
    .B(_03030_),
    .C(_03032_),
    .X(_03033_));
 sky130_fd_sc_hd__or2_1 _06553_ (.A(\tms1x00.ins_pla_ands[21][13] ),
    .B(net887),
    .X(_03034_));
 sky130_fd_sc_hd__o221a_1 _06554_ (.A1(\tms1x00.ins_pla_ands[20][13] ),
    .A2(net797),
    .B1(net770),
    .B2(\tms1x00.ins_pla_ands[23][13] ),
    .C1(_03034_),
    .X(_03035_));
 sky130_fd_sc_hd__o22a_1 _06555_ (.A1(\tms1x00.ins_pla_ands[16][13] ),
    .A2(net825),
    .B1(net744),
    .B2(\tms1x00.ins_pla_ands[17][13] ),
    .X(_03036_));
 sky130_fd_sc_hd__o221a_1 _06556_ (.A1(\tms1x00.ins_pla_ands[22][13] ),
    .A2(net604),
    .B1(net716),
    .B2(\tms1x00.ins_pla_ands[18][13] ),
    .C1(_03036_),
    .X(_03037_));
 sky130_fd_sc_hd__o211a_1 _06557_ (.A1(\tms1x00.ins_pla_ands[19][13] ),
    .A2(net851),
    .B1(_03037_),
    .C1(net912),
    .X(_03038_));
 sky130_fd_sc_hd__a211o_2 _06558_ (.A1(_03035_),
    .A2(_03038_),
    .B1(net924),
    .C1(_03033_),
    .X(_03039_));
 sky130_fd_sc_hd__o211a_2 _06559_ (.A1(_03027_),
    .A2(_03028_),
    .B1(_03039_),
    .C1(net712),
    .X(_03040_));
 sky130_fd_sc_hd__a221o_1 _06560_ (.A1(\tms1x00.ins_pla_ors[5][13] ),
    .A2(net903),
    .B1(net821),
    .B2(\tms1x00.ins_pla_ors[4][13] ),
    .C1(net998),
    .X(_03041_));
 sky130_fd_sc_hd__a22o_1 _06561_ (.A1(\tms1x00.ins_pla_ors[3][13] ),
    .A2(net875),
    .B1(net740),
    .B2(\tms1x00.ins_pla_ors[2][13] ),
    .X(_03042_));
 sky130_fd_sc_hd__a221o_1 _06562_ (.A1(\tms1x00.ins_pla_ors[6][13] ),
    .A2(net627),
    .B1(net767),
    .B2(\tms1x00.ins_pla_ors[1][13] ),
    .C1(_03042_),
    .X(_03043_));
 sky130_fd_sc_hd__a221o_4 _06563_ (.A1(\tms1x00.ins_pla_ors[0][13] ),
    .A2(net848),
    .B1(net794),
    .B2(\tms1x00.ins_pla_ors[7][13] ),
    .C1(_03043_),
    .X(_03044_));
 sky130_fd_sc_hd__a22o_1 _06564_ (.A1(\tms1x00.ins_pla_ors[14][13] ),
    .A2(net628),
    .B1(net795),
    .B2(\tms1x00.ins_pla_ors[15][13] ),
    .X(_03045_));
 sky130_fd_sc_hd__a221o_1 _06565_ (.A1(\tms1x00.ins_pla_ors[13][13] ),
    .A2(net902),
    .B1(net820),
    .B2(\tms1x00.ins_pla_ors[12][13] ),
    .C1(net913),
    .X(_03046_));
 sky130_fd_sc_hd__a22o_1 _06566_ (.A1(\tms1x00.ins_pla_ors[11][13] ),
    .A2(net874),
    .B1(net739),
    .B2(\tms1x00.ins_pla_ors[10][13] ),
    .X(_03047_));
 sky130_fd_sc_hd__a211o_1 _06567_ (.A1(\tms1x00.ins_pla_ors[9][13] ),
    .A2(net766),
    .B1(_03046_),
    .C1(_03047_),
    .X(_03048_));
 sky130_fd_sc_hd__a211o_4 _06568_ (.A1(\tms1x00.ins_pla_ors[8][13] ),
    .A2(net847),
    .B1(_03045_),
    .C1(_03048_),
    .X(_03049_));
 sky130_fd_sc_hd__o21a_2 _06569_ (.A1(_03041_),
    .A2(_03044_),
    .B1(_03049_),
    .X(_03050_));
 sky130_fd_sc_hd__a22o_1 _06570_ (.A1(\tms1x00.O_pla_ors[6][13] ),
    .A2(_02230_),
    .B1(_02240_),
    .B2(\tms1x00.O_pla_ors[7][13] ),
    .X(_03051_));
 sky130_fd_sc_hd__a221o_1 _06571_ (.A1(\tms1x00.O_pla_ors[0][13] ),
    .A2(net848),
    .B1(net768),
    .B2(\tms1x00.O_pla_ors[1][13] ),
    .C1(_01637_),
    .X(_03052_));
 sky130_fd_sc_hd__a22o_1 _06572_ (.A1(\tms1x00.O_pla_ors[3][13] ),
    .A2(net875),
    .B1(net740),
    .B2(\tms1x00.O_pla_ors[2][13] ),
    .X(_03053_));
 sky130_fd_sc_hd__a211o_1 _06573_ (.A1(\tms1x00.O_pla_ors[5][13] ),
    .A2(net903),
    .B1(_03052_),
    .C1(_03053_),
    .X(_03054_));
 sky130_fd_sc_hd__a211o_2 _06574_ (.A1(\tms1x00.O_pla_ors[4][13] ),
    .A2(net821),
    .B1(_03051_),
    .C1(_03054_),
    .X(_03055_));
 sky130_fd_sc_hd__o211a_1 _06575_ (.A1(net85),
    .A2(_03050_),
    .B1(_03055_),
    .C1(net985),
    .X(_03056_));
 sky130_fd_sc_hd__or3_1 _06576_ (.A(net587),
    .B(_03040_),
    .C(_03056_),
    .X(_03057_));
 sky130_fd_sc_hd__and2_1 _06577_ (.A(net910),
    .B(\wbs_o_buff[13] ),
    .X(_03058_));
 sky130_fd_sc_hd__o211a_1 _06578_ (.A1(net590),
    .A2(_03058_),
    .B1(_03057_),
    .C1(_02224_),
    .X(_03059_));
 sky130_fd_sc_hd__a221o_1 _06579_ (.A1(net133),
    .A2(_02313_),
    .B1(_03058_),
    .B2(net585),
    .C1(_03059_),
    .X(_00009_));
 sky130_fd_sc_hd__o22a_1 _06580_ (.A1(\tms1x00.ins_pla_ands[6][14] ),
    .A2(net615),
    .B1(net781),
    .B2(\tms1x00.ins_pla_ands[7][14] ),
    .X(_03060_));
 sky130_fd_sc_hd__o22a_1 _06581_ (.A1(\tms1x00.ins_pla_ands[3][14] ),
    .A2(net858),
    .B1(net724),
    .B2(\tms1x00.ins_pla_ands[2][14] ),
    .X(_03061_));
 sky130_fd_sc_hd__o221a_1 _06582_ (.A1(\tms1x00.ins_pla_ands[5][14] ),
    .A2(net896),
    .B1(net813),
    .B2(\tms1x00.ins_pla_ands[4][14] ),
    .C1(net921),
    .X(_03062_));
 sky130_fd_sc_hd__o211a_1 _06583_ (.A1(\tms1x00.ins_pla_ands[1][14] ),
    .A2(net752),
    .B1(_03061_),
    .C1(_03062_),
    .X(_03063_));
 sky130_fd_sc_hd__o211a_1 _06584_ (.A1(\tms1x00.ins_pla_ands[0][14] ),
    .A2(net835),
    .B1(_03060_),
    .C1(_03063_),
    .X(_03064_));
 sky130_fd_sc_hd__or2_1 _06585_ (.A(\tms1x00.ins_pla_ands[13][14] ),
    .B(net882),
    .X(_03065_));
 sky130_fd_sc_hd__o221a_1 _06586_ (.A1(\tms1x00.ins_pla_ands[14][14] ),
    .A2(net608),
    .B1(net829),
    .B2(\tms1x00.ins_pla_ands[8][14] ),
    .C1(_03065_),
    .X(_03066_));
 sky130_fd_sc_hd__o22a_1 _06587_ (.A1(\tms1x00.ins_pla_ands[15][14] ),
    .A2(net774),
    .B1(net720),
    .B2(\tms1x00.ins_pla_ands[10][14] ),
    .X(_03067_));
 sky130_fd_sc_hd__o221a_2 _06588_ (.A1(\tms1x00.ins_pla_ands[11][14] ),
    .A2(net854),
    .B1(net802),
    .B2(\tms1x00.ins_pla_ands[12][14] ),
    .C1(_03067_),
    .X(_03068_));
 sky130_fd_sc_hd__o211a_1 _06589_ (.A1(\tms1x00.ins_pla_ands[9][14] ),
    .A2(net751),
    .B1(_03068_),
    .C1(net994),
    .X(_03069_));
 sky130_fd_sc_hd__a211o_2 _06590_ (.A1(_03066_),
    .A2(_03069_),
    .B1(net987),
    .C1(_03064_),
    .X(_03070_));
 sky130_fd_sc_hd__o22a_1 _06591_ (.A1(\tms1x00.ins_pla_ands[30][14] ),
    .A2(net602),
    .B1(net823),
    .B2(\tms1x00.ins_pla_ands[24][14] ),
    .X(_03071_));
 sky130_fd_sc_hd__o22a_1 _06592_ (.A1(\tms1x00.ins_pla_ands[27][14] ),
    .A2(net852),
    .B1(net745),
    .B2(\tms1x00.ins_pla_ands[25][14] ),
    .X(_03072_));
 sky130_fd_sc_hd__o221a_1 _06593_ (.A1(\tms1x00.ins_pla_ands[29][14] ),
    .A2(net879),
    .B1(net772),
    .B2(\tms1x00.ins_pla_ands[31][14] ),
    .C1(_03072_),
    .X(_03073_));
 sky130_fd_sc_hd__o211a_1 _06594_ (.A1(\tms1x00.ins_pla_ands[28][14] ),
    .A2(net796),
    .B1(_03073_),
    .C1(net991),
    .X(_03074_));
 sky130_fd_sc_hd__o211a_2 _06595_ (.A1(\tms1x00.ins_pla_ands[26][14] ),
    .A2(net714),
    .B1(_03071_),
    .C1(_03074_),
    .X(_03075_));
 sky130_fd_sc_hd__o22a_1 _06596_ (.A1(\tms1x00.ins_pla_ands[23][14] ),
    .A2(net770),
    .B1(net715),
    .B2(\tms1x00.ins_pla_ands[18][14] ),
    .X(_03076_));
 sky130_fd_sc_hd__o22a_1 _06597_ (.A1(\tms1x00.ins_pla_ands[16][14] ),
    .A2(net825),
    .B1(net744),
    .B2(\tms1x00.ins_pla_ands[17][14] ),
    .X(_03077_));
 sky130_fd_sc_hd__o221a_1 _06598_ (.A1(\tms1x00.ins_pla_ands[21][14] ),
    .A2(net878),
    .B1(net797),
    .B2(\tms1x00.ins_pla_ands[20][14] ),
    .C1(_03077_),
    .X(_03078_));
 sky130_fd_sc_hd__o211a_1 _06599_ (.A1(\tms1x00.ins_pla_ands[19][14] ),
    .A2(net851),
    .B1(_03078_),
    .C1(net912),
    .X(_03079_));
 sky130_fd_sc_hd__o211a_1 _06600_ (.A1(\tms1x00.ins_pla_ands[22][14] ),
    .A2(net604),
    .B1(_03076_),
    .C1(_03079_),
    .X(_03080_));
 sky130_fd_sc_hd__or3_4 _06601_ (.A(net923),
    .B(_03075_),
    .C(_03080_),
    .X(_03081_));
 sky130_fd_sc_hd__a22o_1 _06602_ (.A1(\tms1x00.ins_pla_ors[3][14] ),
    .A2(net875),
    .B1(net794),
    .B2(\tms1x00.ins_pla_ors[7][14] ),
    .X(_03082_));
 sky130_fd_sc_hd__a22o_1 _06603_ (.A1(\tms1x00.ins_pla_ors[5][14] ),
    .A2(net903),
    .B1(net767),
    .B2(\tms1x00.ins_pla_ors[1][14] ),
    .X(_03083_));
 sky130_fd_sc_hd__a221o_1 _06604_ (.A1(\tms1x00.ins_pla_ors[6][14] ),
    .A2(net627),
    .B1(net740),
    .B2(\tms1x00.ins_pla_ors[2][14] ),
    .C1(_03083_),
    .X(_03084_));
 sky130_fd_sc_hd__a211o_1 _06605_ (.A1(\tms1x00.ins_pla_ors[0][14] ),
    .A2(net848),
    .B1(_03084_),
    .C1(net998),
    .X(_03085_));
 sky130_fd_sc_hd__a211o_2 _06606_ (.A1(\tms1x00.ins_pla_ors[4][14] ),
    .A2(net821),
    .B1(_03082_),
    .C1(_03085_),
    .X(_03086_));
 sky130_fd_sc_hd__a22o_1 _06607_ (.A1(\tms1x00.ins_pla_ors[14][14] ),
    .A2(net628),
    .B1(net795),
    .B2(\tms1x00.ins_pla_ors[15][14] ),
    .X(_03087_));
 sky130_fd_sc_hd__a221o_1 _06608_ (.A1(\tms1x00.ins_pla_ors[13][14] ),
    .A2(net902),
    .B1(net820),
    .B2(\tms1x00.ins_pla_ors[12][14] ),
    .C1(net913),
    .X(_03088_));
 sky130_fd_sc_hd__a22o_1 _06609_ (.A1(\tms1x00.ins_pla_ors[11][14] ),
    .A2(net874),
    .B1(net739),
    .B2(\tms1x00.ins_pla_ors[10][14] ),
    .X(_03089_));
 sky130_fd_sc_hd__a211o_1 _06610_ (.A1(\tms1x00.ins_pla_ors[8][14] ),
    .A2(net847),
    .B1(_03088_),
    .C1(_03089_),
    .X(_03090_));
 sky130_fd_sc_hd__a211o_1 _06611_ (.A1(\tms1x00.ins_pla_ors[9][14] ),
    .A2(net766),
    .B1(_03087_),
    .C1(_03090_),
    .X(_03091_));
 sky130_fd_sc_hd__a21o_1 _06612_ (.A1(_03086_),
    .A2(_03091_),
    .B1(net984),
    .X(_03092_));
 sky130_fd_sc_hd__a22o_1 _06613_ (.A1(\tms1x00.O_pla_ors[6][14] ),
    .A2(_02230_),
    .B1(_02240_),
    .B2(\tms1x00.O_pla_ors[7][14] ),
    .X(_03093_));
 sky130_fd_sc_hd__a221o_1 _06614_ (.A1(\tms1x00.O_pla_ors[0][14] ),
    .A2(net849),
    .B1(net768),
    .B2(\tms1x00.O_pla_ors[1][14] ),
    .C1(_01637_),
    .X(_03094_));
 sky130_fd_sc_hd__a22o_1 _06615_ (.A1(\tms1x00.O_pla_ors[3][14] ),
    .A2(net876),
    .B1(net741),
    .B2(\tms1x00.O_pla_ors[2][14] ),
    .X(_03095_));
 sky130_fd_sc_hd__a211o_1 _06616_ (.A1(\tms1x00.O_pla_ors[4][14] ),
    .A2(net822),
    .B1(_03094_),
    .C1(_03095_),
    .X(_03096_));
 sky130_fd_sc_hd__a211o_4 _06617_ (.A1(\tms1x00.O_pla_ors[5][14] ),
    .A2(net904),
    .B1(_03093_),
    .C1(_03096_),
    .X(_03097_));
 sky130_fd_sc_hd__a31o_1 _06618_ (.A1(net985),
    .A2(_03092_),
    .A3(_03097_),
    .B1(net587),
    .X(_03098_));
 sky130_fd_sc_hd__a31o_1 _06619_ (.A1(net712),
    .A2(_03070_),
    .A3(_03081_),
    .B1(_03098_),
    .X(_03099_));
 sky130_fd_sc_hd__and2_1 _06620_ (.A(net907),
    .B(\wbs_o_buff[14] ),
    .X(_03100_));
 sky130_fd_sc_hd__o211a_1 _06621_ (.A1(net589),
    .A2(_03100_),
    .B1(_03099_),
    .C1(net629),
    .X(_03101_));
 sky130_fd_sc_hd__a221o_1 _06622_ (.A1(net134),
    .A2(net579),
    .B1(_03100_),
    .B2(net585),
    .C1(_03101_),
    .X(_00010_));
 sky130_fd_sc_hd__o22a_1 _06623_ (.A1(\tms1x00.ins_pla_ands[6][15] ),
    .A2(net615),
    .B1(net781),
    .B2(\tms1x00.ins_pla_ands[7][15] ),
    .X(_03102_));
 sky130_fd_sc_hd__o221a_1 _06624_ (.A1(\tms1x00.ins_pla_ands[5][15] ),
    .A2(net896),
    .B1(net813),
    .B2(\tms1x00.ins_pla_ands[4][15] ),
    .C1(net921),
    .X(_03103_));
 sky130_fd_sc_hd__o22a_1 _06625_ (.A1(\tms1x00.ins_pla_ands[3][15] ),
    .A2(net858),
    .B1(net724),
    .B2(\tms1x00.ins_pla_ands[2][15] ),
    .X(_03104_));
 sky130_fd_sc_hd__o211a_1 _06626_ (.A1(\tms1x00.ins_pla_ands[1][15] ),
    .A2(net752),
    .B1(_03103_),
    .C1(_03104_),
    .X(_03105_));
 sky130_fd_sc_hd__o211a_1 _06627_ (.A1(\tms1x00.ins_pla_ands[0][15] ),
    .A2(net834),
    .B1(_03102_),
    .C1(_03105_),
    .X(_03106_));
 sky130_fd_sc_hd__o22a_1 _06628_ (.A1(\tms1x00.ins_pla_ands[14][15] ),
    .A2(net608),
    .B1(net774),
    .B2(\tms1x00.ins_pla_ands[15][15] ),
    .X(_03107_));
 sky130_fd_sc_hd__o221a_2 _06629_ (.A1(\tms1x00.ins_pla_ands[8][15] ),
    .A2(net832),
    .B1(net747),
    .B2(\tms1x00.ins_pla_ands[9][15] ),
    .C1(net995),
    .X(_03108_));
 sky130_fd_sc_hd__o22a_1 _06630_ (.A1(\tms1x00.ins_pla_ands[11][15] ),
    .A2(net854),
    .B1(net720),
    .B2(\tms1x00.ins_pla_ands[10][15] ),
    .X(_03109_));
 sky130_fd_sc_hd__o211a_1 _06631_ (.A1(\tms1x00.ins_pla_ands[13][15] ),
    .A2(net883),
    .B1(_03108_),
    .C1(_03109_),
    .X(_03110_));
 sky130_fd_sc_hd__o211a_2 _06632_ (.A1(\tms1x00.ins_pla_ands[12][15] ),
    .A2(net802),
    .B1(_03107_),
    .C1(_03110_),
    .X(_03111_));
 sky130_fd_sc_hd__or3_2 _06633_ (.A(net986),
    .B(_03106_),
    .C(_03111_),
    .X(_03112_));
 sky130_fd_sc_hd__o22a_1 _06634_ (.A1(\tms1x00.ins_pla_ands[30][15] ),
    .A2(net603),
    .B1(net879),
    .B2(\tms1x00.ins_pla_ands[29][15] ),
    .X(_03113_));
 sky130_fd_sc_hd__o22a_1 _06635_ (.A1(\tms1x00.ins_pla_ands[27][15] ),
    .A2(net850),
    .B1(net823),
    .B2(\tms1x00.ins_pla_ands[24][15] ),
    .X(_03114_));
 sky130_fd_sc_hd__o221a_1 _06636_ (.A1(\tms1x00.ins_pla_ands[28][15] ),
    .A2(net796),
    .B1(net769),
    .B2(\tms1x00.ins_pla_ands[31][15] ),
    .C1(_03114_),
    .X(_03115_));
 sky130_fd_sc_hd__o211a_1 _06637_ (.A1(\tms1x00.ins_pla_ands[25][15] ),
    .A2(net743),
    .B1(_03115_),
    .C1(net991),
    .X(_03116_));
 sky130_fd_sc_hd__o211a_1 _06638_ (.A1(\tms1x00.ins_pla_ands[26][15] ),
    .A2(net714),
    .B1(_03113_),
    .C1(_03116_),
    .X(_03117_));
 sky130_fd_sc_hd__o22a_1 _06639_ (.A1(\tms1x00.ins_pla_ands[21][15] ),
    .A2(net887),
    .B1(net770),
    .B2(\tms1x00.ins_pla_ands[23][15] ),
    .X(_03118_));
 sky130_fd_sc_hd__o22a_1 _06640_ (.A1(\tms1x00.ins_pla_ands[16][15] ),
    .A2(net825),
    .B1(net744),
    .B2(\tms1x00.ins_pla_ands[17][15] ),
    .X(_03119_));
 sky130_fd_sc_hd__o221a_1 _06641_ (.A1(\tms1x00.ins_pla_ands[20][15] ),
    .A2(net800),
    .B1(net715),
    .B2(\tms1x00.ins_pla_ands[18][15] ),
    .C1(_03119_),
    .X(_03120_));
 sky130_fd_sc_hd__o211a_1 _06642_ (.A1(\tms1x00.ins_pla_ands[19][15] ),
    .A2(net851),
    .B1(_03120_),
    .C1(net912),
    .X(_03121_));
 sky130_fd_sc_hd__o211a_1 _06643_ (.A1(\tms1x00.ins_pla_ands[22][15] ),
    .A2(net604),
    .B1(_03118_),
    .C1(_03121_),
    .X(_03122_));
 sky130_fd_sc_hd__or3_4 _06644_ (.A(net923),
    .B(_03117_),
    .C(_03122_),
    .X(_03123_));
 sky130_fd_sc_hd__a22o_1 _06645_ (.A1(\tms1x00.ins_pla_ors[3][15] ),
    .A2(net875),
    .B1(net794),
    .B2(\tms1x00.ins_pla_ors[7][15] ),
    .X(_03124_));
 sky130_fd_sc_hd__a22o_1 _06646_ (.A1(\tms1x00.ins_pla_ors[5][15] ),
    .A2(net903),
    .B1(net767),
    .B2(\tms1x00.ins_pla_ors[1][15] ),
    .X(_03125_));
 sky130_fd_sc_hd__a221o_1 _06647_ (.A1(\tms1x00.ins_pla_ors[6][15] ),
    .A2(net627),
    .B1(net740),
    .B2(\tms1x00.ins_pla_ors[2][15] ),
    .C1(_03125_),
    .X(_03126_));
 sky130_fd_sc_hd__a211o_1 _06648_ (.A1(\tms1x00.ins_pla_ors[0][15] ),
    .A2(net848),
    .B1(_03126_),
    .C1(net998),
    .X(_03127_));
 sky130_fd_sc_hd__a211o_2 _06649_ (.A1(\tms1x00.ins_pla_ors[4][15] ),
    .A2(net821),
    .B1(_03124_),
    .C1(_03127_),
    .X(_03128_));
 sky130_fd_sc_hd__a22o_1 _06650_ (.A1(\tms1x00.ins_pla_ors[14][15] ),
    .A2(net628),
    .B1(net795),
    .B2(\tms1x00.ins_pla_ors[15][15] ),
    .X(_03129_));
 sky130_fd_sc_hd__a221o_1 _06651_ (.A1(\tms1x00.ins_pla_ors[13][15] ),
    .A2(net902),
    .B1(net820),
    .B2(\tms1x00.ins_pla_ors[12][15] ),
    .C1(net920),
    .X(_03130_));
 sky130_fd_sc_hd__a22o_1 _06652_ (.A1(\tms1x00.ins_pla_ors[11][15] ),
    .A2(net874),
    .B1(net739),
    .B2(\tms1x00.ins_pla_ors[10][15] ),
    .X(_03131_));
 sky130_fd_sc_hd__a211o_1 _06653_ (.A1(\tms1x00.ins_pla_ors[8][15] ),
    .A2(net847),
    .B1(_03130_),
    .C1(_03131_),
    .X(_03132_));
 sky130_fd_sc_hd__a211o_1 _06654_ (.A1(\tms1x00.ins_pla_ors[9][15] ),
    .A2(net766),
    .B1(_03129_),
    .C1(_03132_),
    .X(_03133_));
 sky130_fd_sc_hd__a21o_1 _06655_ (.A1(_03128_),
    .A2(_03133_),
    .B1(net984),
    .X(_03134_));
 sky130_fd_sc_hd__a22o_1 _06656_ (.A1(\tms1x00.O_pla_ors[6][15] ),
    .A2(_02230_),
    .B1(_02240_),
    .B2(\tms1x00.O_pla_ors[7][15] ),
    .X(_03135_));
 sky130_fd_sc_hd__a221o_1 _06657_ (.A1(\tms1x00.O_pla_ors[0][15] ),
    .A2(net849),
    .B1(net768),
    .B2(\tms1x00.O_pla_ors[1][15] ),
    .C1(_01637_),
    .X(_03136_));
 sky130_fd_sc_hd__a22o_1 _06658_ (.A1(\tms1x00.O_pla_ors[3][15] ),
    .A2(net876),
    .B1(net741),
    .B2(\tms1x00.O_pla_ors[2][15] ),
    .X(_03137_));
 sky130_fd_sc_hd__a211o_1 _06659_ (.A1(\tms1x00.O_pla_ors[5][15] ),
    .A2(net904),
    .B1(_03136_),
    .C1(_03137_),
    .X(_03138_));
 sky130_fd_sc_hd__a211o_4 _06660_ (.A1(\tms1x00.O_pla_ors[4][15] ),
    .A2(net822),
    .B1(_03135_),
    .C1(_03138_),
    .X(_03139_));
 sky130_fd_sc_hd__a31o_1 _06661_ (.A1(net84),
    .A2(_03134_),
    .A3(_03139_),
    .B1(net587),
    .X(_03140_));
 sky130_fd_sc_hd__a31o_1 _06662_ (.A1(net713),
    .A2(_03112_),
    .A3(_03123_),
    .B1(_03140_),
    .X(_03141_));
 sky130_fd_sc_hd__and2_1 _06663_ (.A(net907),
    .B(\wbs_o_buff[15] ),
    .X(_03142_));
 sky130_fd_sc_hd__o211a_1 _06664_ (.A1(net589),
    .A2(_03142_),
    .B1(_03141_),
    .C1(net629),
    .X(_03143_));
 sky130_fd_sc_hd__a221o_1 _06665_ (.A1(net135),
    .A2(net580),
    .B1(_03142_),
    .B2(net584),
    .C1(_03143_),
    .X(_00011_));
 sky130_fd_sc_hd__or2_1 _06666_ (.A(\tms1x00.ins_pla_ors[12][16] ),
    .B(net807),
    .X(_03144_));
 sky130_fd_sc_hd__o221a_1 _06667_ (.A1(\tms1x00.ins_pla_ors[11][16] ),
    .A2(net862),
    .B1(net784),
    .B2(\tms1x00.ins_pla_ors[15][16] ),
    .C1(_03144_),
    .X(_03145_));
 sky130_fd_sc_hd__o22a_1 _06668_ (.A1(\tms1x00.ins_pla_ors[13][16] ),
    .A2(net890),
    .B1(net728),
    .B2(\tms1x00.ins_pla_ors[10][16] ),
    .X(_03146_));
 sky130_fd_sc_hd__o221a_1 _06669_ (.A1(\tms1x00.ins_pla_ors[14][16] ),
    .A2(net617),
    .B1(net757),
    .B2(\tms1x00.ins_pla_ors[9][16] ),
    .C1(_03146_),
    .X(_03147_));
 sky130_fd_sc_hd__o2111a_1 _06670_ (.A1(\tms1x00.ins_pla_ors[8][16] ),
    .A2(net837),
    .B1(_03145_),
    .C1(_03147_),
    .D1(net999),
    .X(_03148_));
 sky130_fd_sc_hd__o22a_1 _06671_ (.A1(\tms1x00.ins_pla_ors[6][16] ),
    .A2(net619),
    .B1(net865),
    .B2(\tms1x00.ins_pla_ors[3][16] ),
    .X(_03149_));
 sky130_fd_sc_hd__o22a_1 _06672_ (.A1(\tms1x00.ins_pla_ors[5][16] ),
    .A2(net891),
    .B1(net811),
    .B2(\tms1x00.ins_pla_ors[4][16] ),
    .X(_03150_));
 sky130_fd_sc_hd__o221a_1 _06673_ (.A1(\tms1x00.ins_pla_ors[0][16] ),
    .A2(net839),
    .B1(net787),
    .B2(\tms1x00.ins_pla_ors[7][16] ),
    .C1(_03150_),
    .X(_03151_));
 sky130_fd_sc_hd__o211a_1 _06674_ (.A1(\tms1x00.ins_pla_ors[1][16] ),
    .A2(net761),
    .B1(_03151_),
    .C1(net919),
    .X(_03152_));
 sky130_fd_sc_hd__o211a_2 _06675_ (.A1(\tms1x00.ins_pla_ors[2][16] ),
    .A2(net731),
    .B1(_03149_),
    .C1(_03152_),
    .X(_03153_));
 sky130_fd_sc_hd__o21a_1 _06676_ (.A1(_03148_),
    .A2(_03153_),
    .B1(net601),
    .X(_03154_));
 sky130_fd_sc_hd__o22a_1 _06677_ (.A1(\tms1x00.O_pla_ors[3][16] ),
    .A2(net872),
    .B1(net737),
    .B2(\tms1x00.O_pla_ors[2][16] ),
    .X(_03155_));
 sky130_fd_sc_hd__o22a_1 _06678_ (.A1(\tms1x00.O_pla_ors[6][16] ),
    .A2(net625),
    .B1(net792),
    .B2(\tms1x00.O_pla_ors[7][16] ),
    .X(_03156_));
 sky130_fd_sc_hd__o221a_1 _06679_ (.A1(\tms1x00.O_pla_ors[0][16] ),
    .A2(net844),
    .B1(net764),
    .B2(\tms1x00.O_pla_ors[1][16] ),
    .C1(_02283_),
    .X(_03157_));
 sky130_fd_sc_hd__o211a_1 _06680_ (.A1(\tms1x00.O_pla_ors[5][16] ),
    .A2(net900),
    .B1(_03155_),
    .C1(_03157_),
    .X(_03158_));
 sky130_fd_sc_hd__o211a_2 _06681_ (.A1(\tms1x00.O_pla_ors[4][16] ),
    .A2(net818),
    .B1(_03156_),
    .C1(_03158_),
    .X(_03159_));
 sky130_fd_sc_hd__a21o_1 _06682_ (.A1(net910),
    .A2(\wbs_o_buff[16] ),
    .B1(net590),
    .X(_03160_));
 sky130_fd_sc_hd__o31a_1 _06683_ (.A1(net588),
    .A2(_03154_),
    .A3(_03159_),
    .B1(_03160_),
    .X(_03161_));
 sky130_fd_sc_hd__mux2_1 _06684_ (.A0(net136),
    .A1(_03161_),
    .S(_02314_),
    .X(_00012_));
 sky130_fd_sc_hd__or2_1 _06685_ (.A(\tms1x00.ins_pla_ors[9][17] ),
    .B(net756),
    .X(_03162_));
 sky130_fd_sc_hd__o221a_1 _06686_ (.A1(\tms1x00.ins_pla_ors[13][17] ),
    .A2(net888),
    .B1(net862),
    .B2(\tms1x00.ins_pla_ors[11][17] ),
    .C1(_03162_),
    .X(_03163_));
 sky130_fd_sc_hd__o22a_1 _06687_ (.A1(\tms1x00.ins_pla_ors[8][17] ),
    .A2(net837),
    .B1(net727),
    .B2(\tms1x00.ins_pla_ors[10][17] ),
    .X(_03164_));
 sky130_fd_sc_hd__o221a_1 _06688_ (.A1(\tms1x00.ins_pla_ors[14][17] ),
    .A2(net616),
    .B1(net806),
    .B2(\tms1x00.ins_pla_ors[12][17] ),
    .C1(_03164_),
    .X(_03165_));
 sky130_fd_sc_hd__o2111a_1 _06689_ (.A1(\tms1x00.ins_pla_ors[15][17] ),
    .A2(net783),
    .B1(_03163_),
    .C1(_03165_),
    .D1(net996),
    .X(_03166_));
 sky130_fd_sc_hd__o22a_1 _06690_ (.A1(\tms1x00.ins_pla_ors[6][17] ),
    .A2(net619),
    .B1(net865),
    .B2(\tms1x00.ins_pla_ors[3][17] ),
    .X(_03167_));
 sky130_fd_sc_hd__o22a_1 _06691_ (.A1(\tms1x00.ins_pla_ors[5][17] ),
    .A2(net892),
    .B1(net785),
    .B2(\tms1x00.ins_pla_ors[7][17] ),
    .X(_03168_));
 sky130_fd_sc_hd__o221a_1 _06692_ (.A1(\tms1x00.ins_pla_ors[0][17] ),
    .A2(net839),
    .B1(net809),
    .B2(\tms1x00.ins_pla_ors[4][17] ),
    .C1(_03168_),
    .X(_03169_));
 sky130_fd_sc_hd__o211a_1 _06693_ (.A1(\tms1x00.ins_pla_ors[1][17] ),
    .A2(net758),
    .B1(_03169_),
    .C1(net919),
    .X(_03170_));
 sky130_fd_sc_hd__o211a_2 _06694_ (.A1(\tms1x00.ins_pla_ors[2][17] ),
    .A2(net731),
    .B1(_03167_),
    .C1(_03170_),
    .X(_03171_));
 sky130_fd_sc_hd__o21a_1 _06695_ (.A1(_03166_),
    .A2(_03171_),
    .B1(net601),
    .X(_03172_));
 sky130_fd_sc_hd__o22a_1 _06696_ (.A1(\tms1x00.O_pla_ors[6][17] ),
    .A2(net626),
    .B1(net789),
    .B2(\tms1x00.O_pla_ors[7][17] ),
    .X(_03173_));
 sky130_fd_sc_hd__o22a_1 _06697_ (.A1(\tms1x00.O_pla_ors[5][17] ),
    .A2(net900),
    .B1(net734),
    .B2(\tms1x00.O_pla_ors[2][17] ),
    .X(_03174_));
 sky130_fd_sc_hd__o221a_1 _06698_ (.A1(\tms1x00.O_pla_ors[0][17] ),
    .A2(net844),
    .B1(net764),
    .B2(\tms1x00.O_pla_ors[1][17] ),
    .C1(net599),
    .X(_03175_));
 sky130_fd_sc_hd__o221a_1 _06699_ (.A1(\tms1x00.O_pla_ors[3][17] ),
    .A2(net872),
    .B1(net818),
    .B2(\tms1x00.O_pla_ors[4][17] ),
    .C1(_03175_),
    .X(_03176_));
 sky130_fd_sc_hd__a31o_1 _06700_ (.A1(_03173_),
    .A2(_03174_),
    .A3(_03176_),
    .B1(net588),
    .X(_03177_));
 sky130_fd_sc_hd__a21o_1 _06701_ (.A1(net910),
    .A2(\wbs_o_buff[17] ),
    .B1(net590),
    .X(_03178_));
 sky130_fd_sc_hd__o21a_1 _06702_ (.A1(_03172_),
    .A2(_03177_),
    .B1(_03178_),
    .X(_03179_));
 sky130_fd_sc_hd__mux2_1 _06703_ (.A0(net137),
    .A1(_03179_),
    .S(_02314_),
    .X(_00013_));
 sky130_fd_sc_hd__nand2_1 _06704_ (.A(net138),
    .B(net581),
    .Y(_03180_));
 sky130_fd_sc_hd__o22a_1 _06705_ (.A1(\tms1x00.ins_pla_ors[6][18] ),
    .A2(net618),
    .B1(net891),
    .B2(\tms1x00.ins_pla_ors[5][18] ),
    .X(_03181_));
 sky130_fd_sc_hd__o22a_1 _06706_ (.A1(\tms1x00.ins_pla_ors[0][18] ),
    .A2(net841),
    .B1(net760),
    .B2(\tms1x00.ins_pla_ors[1][18] ),
    .X(_03182_));
 sky130_fd_sc_hd__o221a_1 _06707_ (.A1(\tms1x00.ins_pla_ors[7][18] ),
    .A2(net787),
    .B1(net731),
    .B2(\tms1x00.ins_pla_ors[2][18] ),
    .C1(_03182_),
    .X(_03183_));
 sky130_fd_sc_hd__o211a_2 _06708_ (.A1(\tms1x00.ins_pla_ors[3][18] ),
    .A2(net865),
    .B1(_03183_),
    .C1(net918),
    .X(_03184_));
 sky130_fd_sc_hd__o211a_1 _06709_ (.A1(\tms1x00.ins_pla_ors[4][18] ),
    .A2(net809),
    .B1(_03181_),
    .C1(_03184_),
    .X(_03185_));
 sky130_fd_sc_hd__or2_1 _06710_ (.A(\tms1x00.ins_pla_ors[10][18] ),
    .B(net727),
    .X(_03186_));
 sky130_fd_sc_hd__o221a_1 _06711_ (.A1(\tms1x00.ins_pla_ors[11][18] ),
    .A2(net863),
    .B1(net783),
    .B2(\tms1x00.ins_pla_ors[15][18] ),
    .C1(_03186_),
    .X(_03187_));
 sky130_fd_sc_hd__o22a_1 _06712_ (.A1(\tms1x00.ins_pla_ors[13][18] ),
    .A2(net888),
    .B1(net837),
    .B2(\tms1x00.ins_pla_ors[8][18] ),
    .X(_03188_));
 sky130_fd_sc_hd__o221a_1 _06713_ (.A1(\tms1x00.ins_pla_ors[14][18] ),
    .A2(net616),
    .B1(net756),
    .B2(\tms1x00.ins_pla_ors[9][18] ),
    .C1(_03188_),
    .X(_03189_));
 sky130_fd_sc_hd__o2111a_1 _06714_ (.A1(\tms1x00.ins_pla_ors[12][18] ),
    .A2(net806),
    .B1(_03187_),
    .C1(_03189_),
    .D1(net996),
    .X(_03190_));
 sky130_fd_sc_hd__o21ai_2 _06715_ (.A1(_03185_),
    .A2(_03190_),
    .B1(net601),
    .Y(_03191_));
 sky130_fd_sc_hd__o22a_1 _06716_ (.A1(\tms1x00.O_pla_ors[5][18] ),
    .A2(net899),
    .B1(net736),
    .B2(\tms1x00.O_pla_ors[2][18] ),
    .X(_03192_));
 sky130_fd_sc_hd__o221a_1 _06717_ (.A1(\tms1x00.O_pla_ors[6][18] ),
    .A2(net625),
    .B1(net791),
    .B2(\tms1x00.O_pla_ors[7][18] ),
    .C1(_03192_),
    .X(_03193_));
 sky130_fd_sc_hd__o221a_1 _06718_ (.A1(\tms1x00.O_pla_ors[0][18] ),
    .A2(net843),
    .B1(net763),
    .B2(\tms1x00.O_pla_ors[1][18] ),
    .C1(net599),
    .X(_03194_));
 sky130_fd_sc_hd__o221a_1 _06719_ (.A1(\tms1x00.O_pla_ors[3][18] ),
    .A2(net873),
    .B1(net816),
    .B2(\tms1x00.O_pla_ors[4][18] ),
    .C1(_03194_),
    .X(_03195_));
 sky130_fd_sc_hd__nand2_2 _06720_ (.A(_03193_),
    .B(_03195_),
    .Y(_03196_));
 sky130_fd_sc_hd__a21oi_1 _06721_ (.A1(net910),
    .A2(\wbs_o_buff[18] ),
    .B1(net590),
    .Y(_03197_));
 sky130_fd_sc_hd__a31o_1 _06722_ (.A1(net590),
    .A2(_03191_),
    .A3(_03196_),
    .B1(_03197_),
    .X(_03198_));
 sky130_fd_sc_hd__o21ai_1 _06723_ (.A1(net581),
    .A2(_03198_),
    .B1(_03180_),
    .Y(_00014_));
 sky130_fd_sc_hd__o22a_1 _06724_ (.A1(\tms1x00.ins_pla_ors[11][19] ),
    .A2(net852),
    .B1(net827),
    .B2(\tms1x00.ins_pla_ors[8][19] ),
    .X(_03199_));
 sky130_fd_sc_hd__o221a_1 _06725_ (.A1(\tms1x00.ins_pla_ors[9][19] ),
    .A2(net745),
    .B1(net717),
    .B2(\tms1x00.ins_pla_ors[10][19] ),
    .C1(_03199_),
    .X(_03200_));
 sky130_fd_sc_hd__or2_1 _06726_ (.A(\tms1x00.ins_pla_ors[4][19] ),
    .B(net809),
    .X(_03201_));
 sky130_fd_sc_hd__or2_1 _06727_ (.A(\tms1x00.ins_pla_ors[3][19] ),
    .B(net865),
    .X(_03202_));
 sky130_fd_sc_hd__o22a_1 _06728_ (.A1(\tms1x00.ins_pla_ors[7][19] ),
    .A2(net785),
    .B1(net731),
    .B2(\tms1x00.ins_pla_ors[2][19] ),
    .X(_03203_));
 sky130_fd_sc_hd__o221a_1 _06729_ (.A1(\tms1x00.ins_pla_ors[0][19] ),
    .A2(net839),
    .B1(net758),
    .B2(\tms1x00.ins_pla_ors[1][19] ),
    .C1(_03202_),
    .X(_03204_));
 sky130_fd_sc_hd__o221a_1 _06730_ (.A1(\tms1x00.ins_pla_ors[6][19] ),
    .A2(net618),
    .B1(net891),
    .B2(\tms1x00.ins_pla_ors[5][19] ),
    .C1(_03201_),
    .X(_03205_));
 sky130_fd_sc_hd__o221a_1 _06731_ (.A1(\tms1x00.ins_pla_ors[13][19] ),
    .A2(net880),
    .B1(net798),
    .B2(\tms1x00.ins_pla_ors[12][19] ),
    .C1(_03200_),
    .X(_03206_));
 sky130_fd_sc_hd__o221a_2 _06732_ (.A1(\tms1x00.ins_pla_ors[14][19] ),
    .A2(net605),
    .B1(net772),
    .B2(\tms1x00.ins_pla_ors[15][19] ),
    .C1(_03206_),
    .X(_03207_));
 sky130_fd_sc_hd__a31o_2 _06733_ (.A1(_03203_),
    .A2(_03204_),
    .A3(_03205_),
    .B1(net998),
    .X(_03208_));
 sky130_fd_sc_hd__o211a_1 _06734_ (.A1(net918),
    .A2(_03207_),
    .B1(_03208_),
    .C1(net601),
    .X(_03209_));
 sky130_fd_sc_hd__o22a_1 _06735_ (.A1(\tms1x00.O_pla_ors[6][19] ),
    .A2(net625),
    .B1(net818),
    .B2(\tms1x00.O_pla_ors[4][19] ),
    .X(_03210_));
 sky130_fd_sc_hd__o22a_1 _06736_ (.A1(\tms1x00.O_pla_ors[3][19] ),
    .A2(net872),
    .B1(net737),
    .B2(\tms1x00.O_pla_ors[2][19] ),
    .X(_03211_));
 sky130_fd_sc_hd__o221a_1 _06737_ (.A1(\tms1x00.O_pla_ors[5][19] ),
    .A2(net900),
    .B1(net792),
    .B2(\tms1x00.O_pla_ors[7][19] ),
    .C1(_03211_),
    .X(_03212_));
 sky130_fd_sc_hd__o211a_1 _06738_ (.A1(\tms1x00.O_pla_ors[0][19] ),
    .A2(net844),
    .B1(_02283_),
    .C1(_03212_),
    .X(_03213_));
 sky130_fd_sc_hd__o211a_2 _06739_ (.A1(\tms1x00.O_pla_ors[1][19] ),
    .A2(net764),
    .B1(_03210_),
    .C1(_03213_),
    .X(_03214_));
 sky130_fd_sc_hd__a21o_1 _06740_ (.A1(net910),
    .A2(\wbs_o_buff[19] ),
    .B1(net590),
    .X(_03215_));
 sky130_fd_sc_hd__o31a_1 _06741_ (.A1(_02228_),
    .A2(_03209_),
    .A3(_03214_),
    .B1(_03215_),
    .X(_03216_));
 sky130_fd_sc_hd__mux2_1 _06742_ (.A0(net139),
    .A1(_03216_),
    .S(_02314_),
    .X(_00015_));
 sky130_fd_sc_hd__and2_4 _06743_ (.A(_02227_),
    .B(net601),
    .X(_03217_));
 sky130_fd_sc_hd__o221a_1 _06744_ (.A1(\tms1x00.ins_pla_ors[13][20] ),
    .A2(net888),
    .B1(net806),
    .B2(\tms1x00.ins_pla_ors[12][20] ),
    .C1(net998),
    .X(_03218_));
 sky130_fd_sc_hd__o22a_1 _06745_ (.A1(\tms1x00.ins_pla_ors[11][20] ),
    .A2(net862),
    .B1(net727),
    .B2(\tms1x00.ins_pla_ors[10][20] ),
    .X(_03219_));
 sky130_fd_sc_hd__o221a_1 _06746_ (.A1(\tms1x00.ins_pla_ors[14][20] ),
    .A2(net616),
    .B1(net756),
    .B2(\tms1x00.ins_pla_ors[9][20] ),
    .C1(_03219_),
    .X(_03220_));
 sky130_fd_sc_hd__o221a_1 _06747_ (.A1(\tms1x00.ins_pla_ors[8][20] ),
    .A2(net838),
    .B1(net783),
    .B2(\tms1x00.ins_pla_ors[15][20] ),
    .C1(_03220_),
    .X(_03221_));
 sky130_fd_sc_hd__o22a_1 _06748_ (.A1(\tms1x00.ins_pla_ors[6][20] ),
    .A2(net621),
    .B1(net729),
    .B2(\tms1x00.ins_pla_ors[2][20] ),
    .X(_03222_));
 sky130_fd_sc_hd__o22a_1 _06749_ (.A1(\tms1x00.ins_pla_ors[0][20] ),
    .A2(net841),
    .B1(net785),
    .B2(\tms1x00.ins_pla_ors[7][20] ),
    .X(_03223_));
 sky130_fd_sc_hd__o221a_1 _06750_ (.A1(\tms1x00.ins_pla_ors[5][20] ),
    .A2(net891),
    .B1(net758),
    .B2(\tms1x00.ins_pla_ors[1][20] ),
    .C1(_03223_),
    .X(_03224_));
 sky130_fd_sc_hd__o211a_1 _06751_ (.A1(\tms1x00.ins_pla_ors[4][20] ),
    .A2(net811),
    .B1(_03224_),
    .C1(net918),
    .X(_03225_));
 sky130_fd_sc_hd__o211a_2 _06752_ (.A1(\tms1x00.ins_pla_ors[3][20] ),
    .A2(net864),
    .B1(_03222_),
    .C1(_03225_),
    .X(_03226_));
 sky130_fd_sc_hd__a21o_1 _06753_ (.A1(_03218_),
    .A2(_03221_),
    .B1(_03226_),
    .X(_03227_));
 sky130_fd_sc_hd__a32o_1 _06754_ (.A1(net908),
    .A2(\wbs_o_buff[20] ),
    .A3(net588),
    .B1(_03217_),
    .B2(_03227_),
    .X(_03228_));
 sky130_fd_sc_hd__a32o_1 _06755_ (.A1(net909),
    .A2(\wbs_o_buff[20] ),
    .A3(net584),
    .B1(_03228_),
    .B2(net630),
    .X(_03229_));
 sky130_fd_sc_hd__a21o_1 _06756_ (.A1(net140),
    .A2(net581),
    .B1(_03229_),
    .X(_00017_));
 sky130_fd_sc_hd__o22a_1 _06757_ (.A1(\tms1x00.ins_pla_ors[13][21] ),
    .A2(net888),
    .B1(net806),
    .B2(\tms1x00.ins_pla_ors[12][21] ),
    .X(_03230_));
 sky130_fd_sc_hd__o22a_1 _06758_ (.A1(\tms1x00.ins_pla_ors[15][21] ),
    .A2(net772),
    .B1(net745),
    .B2(\tms1x00.ins_pla_ors[9][21] ),
    .X(_03231_));
 sky130_fd_sc_hd__o221a_1 _06759_ (.A1(\tms1x00.ins_pla_ors[14][21] ),
    .A2(net605),
    .B1(net827),
    .B2(\tms1x00.ins_pla_ors[8][21] ),
    .C1(_03231_),
    .X(_03232_));
 sky130_fd_sc_hd__o211a_1 _06760_ (.A1(\tms1x00.ins_pla_ors[10][21] ),
    .A2(net717),
    .B1(_03232_),
    .C1(net997),
    .X(_03233_));
 sky130_fd_sc_hd__o211a_4 _06761_ (.A1(\tms1x00.ins_pla_ors[11][21] ),
    .A2(net862),
    .B1(_03230_),
    .C1(_03233_),
    .X(_03234_));
 sky130_fd_sc_hd__or2_1 _06762_ (.A(\tms1x00.ins_pla_ors[2][21] ),
    .B(net729),
    .X(_03235_));
 sky130_fd_sc_hd__o22a_1 _06763_ (.A1(\tms1x00.ins_pla_ors[5][21] ),
    .A2(net891),
    .B1(net864),
    .B2(\tms1x00.ins_pla_ors[3][21] ),
    .X(_03236_));
 sky130_fd_sc_hd__o22a_1 _06764_ (.A1(\tms1x00.ins_pla_ors[0][21] ),
    .A2(net839),
    .B1(net758),
    .B2(\tms1x00.ins_pla_ors[1][21] ),
    .X(_03237_));
 sky130_fd_sc_hd__o221a_1 _06765_ (.A1(\tms1x00.ins_pla_ors[6][21] ),
    .A2(net618),
    .B1(net785),
    .B2(\tms1x00.ins_pla_ors[7][21] ),
    .C1(_03237_),
    .X(_03238_));
 sky130_fd_sc_hd__o211a_1 _06766_ (.A1(\tms1x00.ins_pla_ors[4][21] ),
    .A2(net811),
    .B1(_03238_),
    .C1(net918),
    .X(_03239_));
 sky130_fd_sc_hd__a31o_1 _06767_ (.A1(_03235_),
    .A2(_03236_),
    .A3(_03239_),
    .B1(_03234_),
    .X(_03240_));
 sky130_fd_sc_hd__a32o_1 _06768_ (.A1(net908),
    .A2(\wbs_o_buff[21] ),
    .A3(net588),
    .B1(_03217_),
    .B2(_03240_),
    .X(_03241_));
 sky130_fd_sc_hd__a32o_1 _06769_ (.A1(net908),
    .A2(\wbs_o_buff[21] ),
    .A3(net584),
    .B1(_03241_),
    .B2(net630),
    .X(_03242_));
 sky130_fd_sc_hd__a21o_1 _06770_ (.A1(net141),
    .A2(net581),
    .B1(_03242_),
    .X(_00018_));
 sky130_fd_sc_hd__o22a_1 _06771_ (.A1(\tms1x00.ins_pla_ors[13][22] ),
    .A2(net888),
    .B1(net806),
    .B2(\tms1x00.ins_pla_ors[12][22] ),
    .X(_03243_));
 sky130_fd_sc_hd__o22a_1 _06772_ (.A1(\tms1x00.ins_pla_ors[11][22] ),
    .A2(net862),
    .B1(net756),
    .B2(\tms1x00.ins_pla_ors[9][22] ),
    .X(_03244_));
 sky130_fd_sc_hd__o221a_1 _06773_ (.A1(\tms1x00.ins_pla_ors[14][22] ),
    .A2(net616),
    .B1(net727),
    .B2(\tms1x00.ins_pla_ors[10][22] ),
    .C1(_03244_),
    .X(_03245_));
 sky130_fd_sc_hd__o211a_1 _06774_ (.A1(\tms1x00.ins_pla_ors[8][22] ),
    .A2(net838),
    .B1(_03245_),
    .C1(net997),
    .X(_03246_));
 sky130_fd_sc_hd__o211a_1 _06775_ (.A1(\tms1x00.ins_pla_ors[15][22] ),
    .A2(net784),
    .B1(_03243_),
    .C1(_03246_),
    .X(_03247_));
 sky130_fd_sc_hd__or2_1 _06776_ (.A(\tms1x00.ins_pla_ors[3][22] ),
    .B(net864),
    .X(_03248_));
 sky130_fd_sc_hd__o22a_1 _06777_ (.A1(\tms1x00.ins_pla_ors[4][22] ),
    .A2(net809),
    .B1(net729),
    .B2(\tms1x00.ins_pla_ors[2][22] ),
    .X(_03249_));
 sky130_fd_sc_hd__o22a_1 _06778_ (.A1(\tms1x00.ins_pla_ors[7][22] ),
    .A2(net785),
    .B1(net758),
    .B2(\tms1x00.ins_pla_ors[1][22] ),
    .X(_03250_));
 sky130_fd_sc_hd__o221a_1 _06779_ (.A1(\tms1x00.ins_pla_ors[6][22] ),
    .A2(net618),
    .B1(net839),
    .B2(\tms1x00.ins_pla_ors[0][22] ),
    .C1(_03250_),
    .X(_03251_));
 sky130_fd_sc_hd__o211a_1 _06780_ (.A1(\tms1x00.ins_pla_ors[5][22] ),
    .A2(net891),
    .B1(_03251_),
    .C1(net918),
    .X(_03252_));
 sky130_fd_sc_hd__a31o_1 _06781_ (.A1(_03248_),
    .A2(_03249_),
    .A3(_03252_),
    .B1(_03247_),
    .X(_03253_));
 sky130_fd_sc_hd__a32o_1 _06782_ (.A1(net908),
    .A2(\wbs_o_buff[22] ),
    .A3(net588),
    .B1(_03217_),
    .B2(_03253_),
    .X(_03254_));
 sky130_fd_sc_hd__a32o_1 _06783_ (.A1(net908),
    .A2(\wbs_o_buff[22] ),
    .A3(net584),
    .B1(_03254_),
    .B2(_02224_),
    .X(_03255_));
 sky130_fd_sc_hd__a21o_1 _06784_ (.A1(net142),
    .A2(net581),
    .B1(_03255_),
    .X(_00019_));
 sky130_fd_sc_hd__o22a_1 _06785_ (.A1(\tms1x00.ins_pla_ors[13][23] ),
    .A2(net888),
    .B1(net806),
    .B2(\tms1x00.ins_pla_ors[12][23] ),
    .X(_03256_));
 sky130_fd_sc_hd__o22a_1 _06786_ (.A1(\tms1x00.ins_pla_ors[8][23] ),
    .A2(net837),
    .B1(net783),
    .B2(\tms1x00.ins_pla_ors[15][23] ),
    .X(_03257_));
 sky130_fd_sc_hd__o221a_1 _06787_ (.A1(\tms1x00.ins_pla_ors[14][23] ),
    .A2(net616),
    .B1(net756),
    .B2(\tms1x00.ins_pla_ors[9][23] ),
    .C1(_03257_),
    .X(_03258_));
 sky130_fd_sc_hd__o211a_1 _06788_ (.A1(\tms1x00.ins_pla_ors[10][23] ),
    .A2(net727),
    .B1(_03258_),
    .C1(net997),
    .X(_03259_));
 sky130_fd_sc_hd__o211a_4 _06789_ (.A1(\tms1x00.ins_pla_ors[11][23] ),
    .A2(net863),
    .B1(_03256_),
    .C1(_03259_),
    .X(_03260_));
 sky130_fd_sc_hd__or2_1 _06790_ (.A(\tms1x00.ins_pla_ors[3][23] ),
    .B(net866),
    .X(_03261_));
 sky130_fd_sc_hd__o22a_1 _06791_ (.A1(\tms1x00.ins_pla_ors[6][23] ),
    .A2(net619),
    .B1(net730),
    .B2(\tms1x00.ins_pla_ors[2][23] ),
    .X(_03262_));
 sky130_fd_sc_hd__o22a_1 _06792_ (.A1(\tms1x00.ins_pla_ors[0][23] ),
    .A2(net840),
    .B1(net786),
    .B2(\tms1x00.ins_pla_ors[7][23] ),
    .X(_03263_));
 sky130_fd_sc_hd__o221a_1 _06793_ (.A1(\tms1x00.ins_pla_ors[4][23] ),
    .A2(net810),
    .B1(net759),
    .B2(\tms1x00.ins_pla_ors[1][23] ),
    .C1(_03263_),
    .X(_03264_));
 sky130_fd_sc_hd__o211a_1 _06794_ (.A1(\tms1x00.ins_pla_ors[5][23] ),
    .A2(net892),
    .B1(_03264_),
    .C1(net919),
    .X(_03265_));
 sky130_fd_sc_hd__a31o_4 _06795_ (.A1(_03261_),
    .A2(_03262_),
    .A3(_03265_),
    .B1(_03260_),
    .X(_03266_));
 sky130_fd_sc_hd__a32o_1 _06796_ (.A1(net908),
    .A2(\wbs_o_buff[23] ),
    .A3(net588),
    .B1(_03217_),
    .B2(_03266_),
    .X(_03267_));
 sky130_fd_sc_hd__a32o_1 _06797_ (.A1(net908),
    .A2(\wbs_o_buff[23] ),
    .A3(net584),
    .B1(_03267_),
    .B2(net630),
    .X(_03268_));
 sky130_fd_sc_hd__a21o_1 _06798_ (.A1(net143),
    .A2(net581),
    .B1(_03268_),
    .X(_00020_));
 sky130_fd_sc_hd__o22a_1 _06799_ (.A1(\tms1x00.ins_pla_ors[13][24] ),
    .A2(net890),
    .B1(net808),
    .B2(\tms1x00.ins_pla_ors[12][24] ),
    .X(_03269_));
 sky130_fd_sc_hd__o22a_1 _06800_ (.A1(\tms1x00.ins_pla_ors[11][24] ),
    .A2(net863),
    .B1(net784),
    .B2(\tms1x00.ins_pla_ors[15][24] ),
    .X(_03270_));
 sky130_fd_sc_hd__o221a_1 _06801_ (.A1(\tms1x00.ins_pla_ors[14][24] ),
    .A2(net617),
    .B1(net728),
    .B2(\tms1x00.ins_pla_ors[10][24] ),
    .C1(_03270_),
    .X(_03271_));
 sky130_fd_sc_hd__o211a_1 _06802_ (.A1(\tms1x00.ins_pla_ors[9][24] ),
    .A2(net757),
    .B1(_03271_),
    .C1(net997),
    .X(_03272_));
 sky130_fd_sc_hd__o211a_2 _06803_ (.A1(\tms1x00.ins_pla_ors[8][24] ),
    .A2(net838),
    .B1(_03269_),
    .C1(_03272_),
    .X(_03273_));
 sky130_fd_sc_hd__or2_1 _06804_ (.A(\tms1x00.ins_pla_ors[3][24] ),
    .B(net866),
    .X(_03274_));
 sky130_fd_sc_hd__o22a_1 _06805_ (.A1(\tms1x00.ins_pla_ors[4][24] ),
    .A2(net810),
    .B1(net730),
    .B2(\tms1x00.ins_pla_ors[2][24] ),
    .X(_03275_));
 sky130_fd_sc_hd__o22a_1 _06806_ (.A1(\tms1x00.ins_pla_ors[7][24] ),
    .A2(net787),
    .B1(net760),
    .B2(\tms1x00.ins_pla_ors[1][24] ),
    .X(_03276_));
 sky130_fd_sc_hd__o221a_2 _06807_ (.A1(\tms1x00.ins_pla_ors[6][24] ),
    .A2(net620),
    .B1(net841),
    .B2(\tms1x00.ins_pla_ors[0][24] ),
    .C1(_03276_),
    .X(_03277_));
 sky130_fd_sc_hd__o211a_1 _06808_ (.A1(\tms1x00.ins_pla_ors[5][24] ),
    .A2(net892),
    .B1(_03277_),
    .C1(net919),
    .X(_03278_));
 sky130_fd_sc_hd__a31o_1 _06809_ (.A1(_03274_),
    .A2(_03275_),
    .A3(_03278_),
    .B1(_03273_),
    .X(_03279_));
 sky130_fd_sc_hd__a32o_1 _06810_ (.A1(net910),
    .A2(\wbs_o_buff[24] ),
    .A3(net588),
    .B1(_03217_),
    .B2(_03279_),
    .X(_03280_));
 sky130_fd_sc_hd__a32o_1 _06811_ (.A1(net910),
    .A2(\wbs_o_buff[24] ),
    .A3(net584),
    .B1(_03280_),
    .B2(_02224_),
    .X(_03281_));
 sky130_fd_sc_hd__a21o_1 _06812_ (.A1(\tms1x00.status ),
    .A2(net581),
    .B1(_03281_),
    .X(_00021_));
 sky130_fd_sc_hd__or2_1 _06813_ (.A(\tms1x00.ins_pla_ors[2][25] ),
    .B(net729),
    .X(_03282_));
 sky130_fd_sc_hd__o22a_1 _06814_ (.A1(\tms1x00.ins_pla_ors[6][25] ),
    .A2(net618),
    .B1(net864),
    .B2(\tms1x00.ins_pla_ors[3][25] ),
    .X(_03283_));
 sky130_fd_sc_hd__o22a_1 _06815_ (.A1(\tms1x00.ins_pla_ors[0][25] ),
    .A2(net839),
    .B1(net758),
    .B2(\tms1x00.ins_pla_ors[1][25] ),
    .X(_03284_));
 sky130_fd_sc_hd__o221a_1 _06816_ (.A1(\tms1x00.ins_pla_ors[5][25] ),
    .A2(net891),
    .B1(net785),
    .B2(\tms1x00.ins_pla_ors[7][25] ),
    .C1(_03284_),
    .X(_03285_));
 sky130_fd_sc_hd__o211a_1 _06817_ (.A1(\tms1x00.ins_pla_ors[4][25] ),
    .A2(net809),
    .B1(_03285_),
    .C1(net918),
    .X(_03286_));
 sky130_fd_sc_hd__o22a_1 _06818_ (.A1(\tms1x00.ins_pla_ors[13][25] ),
    .A2(net888),
    .B1(net806),
    .B2(\tms1x00.ins_pla_ors[12][25] ),
    .X(_03287_));
 sky130_fd_sc_hd__o22a_1 _06819_ (.A1(\tms1x00.ins_pla_ors[15][25] ),
    .A2(net783),
    .B1(net756),
    .B2(\tms1x00.ins_pla_ors[9][25] ),
    .X(_03288_));
 sky130_fd_sc_hd__o221a_1 _06820_ (.A1(\tms1x00.ins_pla_ors[14][25] ),
    .A2(net616),
    .B1(net727),
    .B2(\tms1x00.ins_pla_ors[10][25] ),
    .C1(_03288_),
    .X(_03289_));
 sky130_fd_sc_hd__o211a_1 _06821_ (.A1(\tms1x00.ins_pla_ors[11][25] ),
    .A2(net862),
    .B1(_03289_),
    .C1(net997),
    .X(_03290_));
 sky130_fd_sc_hd__o211a_2 _06822_ (.A1(\tms1x00.ins_pla_ors[8][25] ),
    .A2(net837),
    .B1(_03287_),
    .C1(_03290_),
    .X(_03291_));
 sky130_fd_sc_hd__a31o_1 _06823_ (.A1(_03282_),
    .A2(_03283_),
    .A3(_03286_),
    .B1(_03291_),
    .X(_03292_));
 sky130_fd_sc_hd__a32o_1 _06824_ (.A1(net909),
    .A2(\wbs_o_buff[25] ),
    .A3(net588),
    .B1(_03217_),
    .B2(_03292_),
    .X(_03293_));
 sky130_fd_sc_hd__a32o_1 _06825_ (.A1(net909),
    .A2(\wbs_o_buff[25] ),
    .A3(net584),
    .B1(_03293_),
    .B2(net630),
    .X(_03294_));
 sky130_fd_sc_hd__a21o_1 _06826_ (.A1(\tms1x00.X[0] ),
    .A2(net581),
    .B1(_03294_),
    .X(_00022_));
 sky130_fd_sc_hd__o22a_1 _06827_ (.A1(\tms1x00.ins_pla_ors[13][26] ),
    .A2(net888),
    .B1(net806),
    .B2(\tms1x00.ins_pla_ors[12][26] ),
    .X(_03295_));
 sky130_fd_sc_hd__o22a_1 _06828_ (.A1(\tms1x00.ins_pla_ors[15][26] ),
    .A2(net783),
    .B1(net756),
    .B2(\tms1x00.ins_pla_ors[9][26] ),
    .X(_03296_));
 sky130_fd_sc_hd__o221a_1 _06829_ (.A1(\tms1x00.ins_pla_ors[14][26] ),
    .A2(net616),
    .B1(net727),
    .B2(\tms1x00.ins_pla_ors[10][26] ),
    .C1(_03296_),
    .X(_03297_));
 sky130_fd_sc_hd__o211a_1 _06830_ (.A1(\tms1x00.ins_pla_ors[8][26] ),
    .A2(net837),
    .B1(_03297_),
    .C1(net997),
    .X(_03298_));
 sky130_fd_sc_hd__o211a_1 _06831_ (.A1(\tms1x00.ins_pla_ors[11][26] ),
    .A2(net862),
    .B1(_03295_),
    .C1(_03298_),
    .X(_03299_));
 sky130_fd_sc_hd__or2_1 _06832_ (.A(\tms1x00.ins_pla_ors[2][26] ),
    .B(net729),
    .X(_03300_));
 sky130_fd_sc_hd__o22a_2 _06833_ (.A1(\tms1x00.ins_pla_ors[6][26] ),
    .A2(net618),
    .B1(net865),
    .B2(\tms1x00.ins_pla_ors[3][26] ),
    .X(_03301_));
 sky130_fd_sc_hd__o22a_1 _06834_ (.A1(\tms1x00.ins_pla_ors[0][26] ),
    .A2(net839),
    .B1(net758),
    .B2(\tms1x00.ins_pla_ors[1][26] ),
    .X(_03302_));
 sky130_fd_sc_hd__o221a_1 _06835_ (.A1(\tms1x00.ins_pla_ors[5][26] ),
    .A2(net891),
    .B1(net785),
    .B2(\tms1x00.ins_pla_ors[7][26] ),
    .C1(_03302_),
    .X(_03303_));
 sky130_fd_sc_hd__o211a_1 _06836_ (.A1(\tms1x00.ins_pla_ors[4][26] ),
    .A2(net809),
    .B1(_03303_),
    .C1(net918),
    .X(_03304_));
 sky130_fd_sc_hd__a31o_1 _06837_ (.A1(_03300_),
    .A2(_03301_),
    .A3(_03304_),
    .B1(_03299_),
    .X(_03305_));
 sky130_fd_sc_hd__a32o_1 _06838_ (.A1(net908),
    .A2(\wbs_o_buff[26] ),
    .A3(net588),
    .B1(_03217_),
    .B2(_03305_),
    .X(_03306_));
 sky130_fd_sc_hd__a32o_1 _06839_ (.A1(net908),
    .A2(\wbs_o_buff[26] ),
    .A3(net584),
    .B1(_03306_),
    .B2(net630),
    .X(_03307_));
 sky130_fd_sc_hd__a21o_1 _06840_ (.A1(\tms1x00.X[1] ),
    .A2(net581),
    .B1(_03307_),
    .X(_00023_));
 sky130_fd_sc_hd__or2_1 _06841_ (.A(\tms1x00.ins_pla_ors[2][27] ),
    .B(net729),
    .X(_03308_));
 sky130_fd_sc_hd__o22a_1 _06842_ (.A1(\tms1x00.ins_pla_ors[6][27] ),
    .A2(net618),
    .B1(net864),
    .B2(\tms1x00.ins_pla_ors[3][27] ),
    .X(_03309_));
 sky130_fd_sc_hd__o22a_1 _06843_ (.A1(\tms1x00.ins_pla_ors[0][27] ),
    .A2(net839),
    .B1(net758),
    .B2(\tms1x00.ins_pla_ors[1][27] ),
    .X(_03310_));
 sky130_fd_sc_hd__o221a_1 _06844_ (.A1(\tms1x00.ins_pla_ors[4][27] ),
    .A2(net809),
    .B1(net785),
    .B2(\tms1x00.ins_pla_ors[7][27] ),
    .C1(_03310_),
    .X(_03311_));
 sky130_fd_sc_hd__o211a_1 _06845_ (.A1(\tms1x00.ins_pla_ors[5][27] ),
    .A2(net891),
    .B1(_03311_),
    .C1(net918),
    .X(_03312_));
 sky130_fd_sc_hd__o22a_1 _06846_ (.A1(\tms1x00.ins_pla_ors[13][27] ),
    .A2(net889),
    .B1(net808),
    .B2(\tms1x00.ins_pla_ors[12][27] ),
    .X(_03313_));
 sky130_fd_sc_hd__o22a_1 _06847_ (.A1(\tms1x00.ins_pla_ors[15][27] ),
    .A2(net783),
    .B1(net756),
    .B2(\tms1x00.ins_pla_ors[9][27] ),
    .X(_03314_));
 sky130_fd_sc_hd__o221a_1 _06848_ (.A1(\tms1x00.ins_pla_ors[14][27] ),
    .A2(net616),
    .B1(net728),
    .B2(\tms1x00.ins_pla_ors[10][27] ),
    .C1(_03314_),
    .X(_03315_));
 sky130_fd_sc_hd__o211a_1 _06849_ (.A1(\tms1x00.ins_pla_ors[11][27] ),
    .A2(net862),
    .B1(_03315_),
    .C1(net997),
    .X(_03316_));
 sky130_fd_sc_hd__o211a_1 _06850_ (.A1(\tms1x00.ins_pla_ors[8][27] ),
    .A2(net837),
    .B1(_03313_),
    .C1(_03316_),
    .X(_03317_));
 sky130_fd_sc_hd__a31o_1 _06851_ (.A1(_03308_),
    .A2(_03309_),
    .A3(_03312_),
    .B1(_03317_),
    .X(_03318_));
 sky130_fd_sc_hd__a32o_1 _06852_ (.A1(net909),
    .A2(\wbs_o_buff[27] ),
    .A3(net588),
    .B1(_03217_),
    .B2(_03318_),
    .X(_03319_));
 sky130_fd_sc_hd__a32o_1 _06853_ (.A1(net908),
    .A2(\wbs_o_buff[27] ),
    .A3(net584),
    .B1(_03319_),
    .B2(net630),
    .X(_03320_));
 sky130_fd_sc_hd__a21o_1 _06854_ (.A1(\tms1x00.X[2] ),
    .A2(net581),
    .B1(_03320_),
    .X(_00024_));
 sky130_fd_sc_hd__nor2_8 _06855_ (.A(net74),
    .B(net590),
    .Y(_03321_));
 sky130_fd_sc_hd__o22a_1 _06856_ (.A1(\tms1x00.ins_pla_ors[15][28] ),
    .A2(net783),
    .B1(net727),
    .B2(\tms1x00.ins_pla_ors[10][28] ),
    .X(_03322_));
 sky130_fd_sc_hd__o22a_1 _06857_ (.A1(\tms1x00.ins_pla_ors[8][28] ),
    .A2(net837),
    .B1(net757),
    .B2(\tms1x00.ins_pla_ors[9][28] ),
    .X(_03323_));
 sky130_fd_sc_hd__o221a_1 _06858_ (.A1(\tms1x00.ins_pla_ors[14][28] ),
    .A2(net616),
    .B1(net806),
    .B2(\tms1x00.ins_pla_ors[12][28] ),
    .C1(_03323_),
    .X(_03324_));
 sky130_fd_sc_hd__o211a_1 _06859_ (.A1(\tms1x00.ins_pla_ors[13][28] ),
    .A2(net889),
    .B1(_03324_),
    .C1(net998),
    .X(_03325_));
 sky130_fd_sc_hd__o211a_1 _06860_ (.A1(\tms1x00.ins_pla_ors[11][28] ),
    .A2(net862),
    .B1(_03322_),
    .C1(_03325_),
    .X(_03326_));
 sky130_fd_sc_hd__or2_1 _06861_ (.A(\tms1x00.ins_pla_ors[0][28] ),
    .B(net841),
    .X(_03327_));
 sky130_fd_sc_hd__o22a_1 _06862_ (.A1(\tms1x00.ins_pla_ors[5][28] ),
    .A2(net892),
    .B1(net758),
    .B2(\tms1x00.ins_pla_ors[1][28] ),
    .X(_03328_));
 sky130_fd_sc_hd__o22a_1 _06863_ (.A1(\tms1x00.ins_pla_ors[4][28] ),
    .A2(net809),
    .B1(net785),
    .B2(\tms1x00.ins_pla_ors[7][28] ),
    .X(_03329_));
 sky130_fd_sc_hd__o221a_1 _06864_ (.A1(\tms1x00.ins_pla_ors[6][28] ),
    .A2(net618),
    .B1(net729),
    .B2(\tms1x00.ins_pla_ors[2][28] ),
    .C1(_03329_),
    .X(_03330_));
 sky130_fd_sc_hd__o211a_1 _06865_ (.A1(\tms1x00.ins_pla_ors[3][28] ),
    .A2(net864),
    .B1(_03330_),
    .C1(net918),
    .X(_03331_));
 sky130_fd_sc_hd__a31o_1 _06866_ (.A1(_03327_),
    .A2(_03328_),
    .A3(_03331_),
    .B1(_03326_),
    .X(_03332_));
 sky130_fd_sc_hd__a22o_1 _06867_ (.A1(\wbs_o_buff[28] ),
    .A2(_03321_),
    .B1(_03332_),
    .B2(_03217_),
    .X(_03333_));
 sky130_fd_sc_hd__and2_1 _06868_ (.A(_02314_),
    .B(_03333_),
    .X(_00025_));
 sky130_fd_sc_hd__or2_1 _06869_ (.A(\tms1x00.ins_pla_ors[15][29] ),
    .B(net784),
    .X(_03334_));
 sky130_fd_sc_hd__o221a_1 _06870_ (.A1(\tms1x00.ins_pla_ors[13][29] ),
    .A2(net889),
    .B1(net808),
    .B2(\tms1x00.ins_pla_ors[12][29] ),
    .C1(_03334_),
    .X(_03335_));
 sky130_fd_sc_hd__o22a_1 _06871_ (.A1(\tms1x00.ins_pla_ors[11][29] ),
    .A2(net863),
    .B1(net728),
    .B2(\tms1x00.ins_pla_ors[10][29] ),
    .X(_03336_));
 sky130_fd_sc_hd__o221a_1 _06872_ (.A1(\tms1x00.ins_pla_ors[8][29] ),
    .A2(net837),
    .B1(net756),
    .B2(\tms1x00.ins_pla_ors[9][29] ),
    .C1(_03336_),
    .X(_03337_));
 sky130_fd_sc_hd__o2111a_1 _06873_ (.A1(\tms1x00.ins_pla_ors[14][29] ),
    .A2(net616),
    .B1(_03335_),
    .C1(_03337_),
    .D1(net998),
    .X(_03338_));
 sky130_fd_sc_hd__or2_1 _06874_ (.A(\tms1x00.ins_pla_ors[0][29] ),
    .B(net839),
    .X(_03339_));
 sky130_fd_sc_hd__o22a_1 _06875_ (.A1(\tms1x00.ins_pla_ors[5][29] ),
    .A2(net891),
    .B1(net758),
    .B2(\tms1x00.ins_pla_ors[1][29] ),
    .X(_03340_));
 sky130_fd_sc_hd__o22a_1 _06876_ (.A1(\tms1x00.ins_pla_ors[3][29] ),
    .A2(net864),
    .B1(net729),
    .B2(\tms1x00.ins_pla_ors[2][29] ),
    .X(_03341_));
 sky130_fd_sc_hd__o221a_1 _06877_ (.A1(\tms1x00.ins_pla_ors[4][29] ),
    .A2(net809),
    .B1(net785),
    .B2(\tms1x00.ins_pla_ors[7][29] ),
    .C1(_03341_),
    .X(_03342_));
 sky130_fd_sc_hd__o211a_1 _06878_ (.A1(\tms1x00.ins_pla_ors[6][29] ),
    .A2(net618),
    .B1(_03342_),
    .C1(net918),
    .X(_03343_));
 sky130_fd_sc_hd__a31o_1 _06879_ (.A1(_03339_),
    .A2(_03340_),
    .A3(_03343_),
    .B1(_03338_),
    .X(_03344_));
 sky130_fd_sc_hd__a22o_1 _06880_ (.A1(\wbs_o_buff[29] ),
    .A2(_03321_),
    .B1(_03344_),
    .B2(_03217_),
    .X(_03345_));
 sky130_fd_sc_hd__and2_1 _06881_ (.A(_02314_),
    .B(_03345_),
    .X(_00026_));
 sky130_fd_sc_hd__and3_1 _06882_ (.A(\wbs_o_buff[30] ),
    .B(_02314_),
    .C(_03321_),
    .X(_00028_));
 sky130_fd_sc_hd__and3_1 _06883_ (.A(\wbs_o_buff[31] ),
    .B(_02314_),
    .C(_03321_),
    .X(_00029_));
 sky130_fd_sc_hd__nor2_4 _06884_ (.A(net74),
    .B(net582),
    .Y(_03346_));
 sky130_fd_sc_hd__a32o_1 _06885_ (.A1(net1055),
    .A2(net979),
    .A3(net582),
    .B1(_03346_),
    .B2(chip_sel_override),
    .X(_00000_));
 sky130_fd_sc_hd__a22o_1 _06886_ (.A1(net1049),
    .A2(net583),
    .B1(_03346_),
    .B2(\tms1x00.pla_override ),
    .X(_00002_));
 sky130_fd_sc_hd__a32o_1 _06887_ (.A1(net930),
    .A2(net979),
    .A3(net582),
    .B1(_03346_),
    .B2(wb_rst_override),
    .X(_00003_));
 sky130_fd_sc_hd__a32o_1 _06888_ (.A1(net1066),
    .A2(net979),
    .A3(net582),
    .B1(_03346_),
    .B2(\tms1x00.wb_step ),
    .X(_00004_));
 sky130_fd_sc_hd__a22o_1 _06889_ (.A1(net979),
    .A2(net582),
    .B1(_03346_),
    .B2(net145),
    .X(_00001_));
 sky130_fd_sc_hd__nand2_4 _06890_ (.A(net76),
    .B(valid),
    .Y(net177));
 sky130_fd_sc_hd__nor2_8 _06891_ (.A(net178),
    .B(_02226_),
    .Y(_03347_));
 sky130_fd_sc_hd__or2_4 _06892_ (.A(net178),
    .B(_02226_),
    .X(_03348_));
 sky130_fd_sc_hd__and2_4 _06893_ (.A(\tms1x00.pla_override ),
    .B(net592),
    .X(_03349_));
 sky130_fd_sc_hd__nand2_2 _06894_ (.A(\tms1x00.pla_override ),
    .B(net592),
    .Y(_03350_));
 sky130_fd_sc_hd__or3_4 _06895_ (.A(_02775_),
    .B(_03348_),
    .C(_03350_),
    .X(_03351_));
 sky130_fd_sc_hd__nor2_2 _06896_ (.A(net925),
    .B(net995),
    .Y(_03352_));
 sky130_fd_sc_hd__nand2_8 _06897_ (.A(net987),
    .B(net917),
    .Y(_03353_));
 sky130_fd_sc_hd__nor2_8 _06898_ (.A(\tms1x00.pla_override ),
    .B(net637),
    .Y(_03354_));
 sky130_fd_sc_hd__or2_4 _06899_ (.A(\tms1x00.pla_override ),
    .B(net637),
    .X(_03355_));
 sky130_fd_sc_hd__and3_4 _06900_ (.A(_02774_),
    .B(_03347_),
    .C(_03349_),
    .X(_03356_));
 sky130_fd_sc_hd__or3_4 _06901_ (.A(_02775_),
    .B(_03348_),
    .C(_03350_),
    .X(_03357_));
 sky130_fd_sc_hd__and3_4 _06902_ (.A(net739),
    .B(net598),
    .C(net359),
    .X(_03358_));
 sky130_fd_sc_hd__or3_4 _06903_ (.A(net724),
    .B(_03353_),
    .C(net357),
    .X(_03359_));
 sky130_fd_sc_hd__or2_1 _06904_ (.A(\tms1x00.O_pla_ands[18][0] ),
    .B(_03358_),
    .X(_03360_));
 sky130_fd_sc_hd__o211a_1 _06905_ (.A1(net977),
    .A2(_03359_),
    .B1(_03360_),
    .C1(net473),
    .X(_00037_));
 sky130_fd_sc_hd__or2_1 _06906_ (.A(\tms1x00.O_pla_ands[18][1] ),
    .B(_03358_),
    .X(_03361_));
 sky130_fd_sc_hd__o211a_1 _06907_ (.A1(net929),
    .A2(_03359_),
    .B1(_03361_),
    .C1(net473),
    .X(_00038_));
 sky130_fd_sc_hd__or2_1 _06908_ (.A(\tms1x00.O_pla_ands[18][2] ),
    .B(_03358_),
    .X(_03362_));
 sky130_fd_sc_hd__o211a_1 _06909_ (.A1(net1063),
    .A2(_03359_),
    .B1(_03362_),
    .C1(net474),
    .X(_00039_));
 sky130_fd_sc_hd__or2_1 _06910_ (.A(\tms1x00.O_pla_ands[18][3] ),
    .B(_03358_),
    .X(_03363_));
 sky130_fd_sc_hd__o211a_1 _06911_ (.A1(net1056),
    .A2(_03359_),
    .B1(_03363_),
    .C1(net473),
    .X(_00040_));
 sky130_fd_sc_hd__or2_1 _06912_ (.A(\tms1x00.O_pla_ands[18][4] ),
    .B(_03358_),
    .X(_03364_));
 sky130_fd_sc_hd__o211a_1 _06913_ (.A1(net1048),
    .A2(_03359_),
    .B1(_03364_),
    .C1(net473),
    .X(_00041_));
 sky130_fd_sc_hd__a21o_1 _06914_ (.A1(net1040),
    .A2(_03358_),
    .B1(net534),
    .X(_03365_));
 sky130_fd_sc_hd__a21o_1 _06915_ (.A1(\tms1x00.O_pla_ands[18][5] ),
    .A2(_03359_),
    .B1(_03365_),
    .X(_00042_));
 sky130_fd_sc_hd__or2_1 _06916_ (.A(\tms1x00.O_pla_ands[18][6] ),
    .B(_03358_),
    .X(_03366_));
 sky130_fd_sc_hd__o211a_1 _06917_ (.A1(net1031),
    .A2(_03359_),
    .B1(_03366_),
    .C1(net473),
    .X(_00043_));
 sky130_fd_sc_hd__or2_1 _06918_ (.A(\tms1x00.O_pla_ands[18][7] ),
    .B(_03358_),
    .X(_03367_));
 sky130_fd_sc_hd__o211a_1 _06919_ (.A1(net1025),
    .A2(_03359_),
    .B1(_03367_),
    .C1(net473),
    .X(_00044_));
 sky130_fd_sc_hd__a21o_1 _06920_ (.A1(net1017),
    .A2(_03358_),
    .B1(net534),
    .X(_03368_));
 sky130_fd_sc_hd__a21o_1 _06921_ (.A1(\tms1x00.O_pla_ands[18][8] ),
    .A2(_03359_),
    .B1(_03368_),
    .X(_00045_));
 sky130_fd_sc_hd__or2_1 _06922_ (.A(\tms1x00.O_pla_ands[18][9] ),
    .B(_03358_),
    .X(_03369_));
 sky130_fd_sc_hd__o211a_1 _06923_ (.A1(net1009),
    .A2(_03359_),
    .B1(_03369_),
    .C1(net474),
    .X(_00046_));
 sky130_fd_sc_hd__or3_4 _06924_ (.A(net803),
    .B(net361),
    .C(_03353_),
    .X(_03370_));
 sky130_fd_sc_hd__mux2_1 _06925_ (.A0(net977),
    .A1(\tms1x00.O_pla_ands[20][0] ),
    .S(_03370_),
    .X(_00047_));
 sky130_fd_sc_hd__mux2_1 _06926_ (.A0(net927),
    .A1(\tms1x00.O_pla_ands[20][1] ),
    .S(_03370_),
    .X(_00048_));
 sky130_fd_sc_hd__mux2_1 _06927_ (.A0(net1063),
    .A1(\tms1x00.O_pla_ands[20][2] ),
    .S(_03370_),
    .X(_00049_));
 sky130_fd_sc_hd__mux2_1 _06928_ (.A0(net1056),
    .A1(\tms1x00.O_pla_ands[20][3] ),
    .S(_03370_),
    .X(_00050_));
 sky130_fd_sc_hd__mux2_1 _06929_ (.A0(net1048),
    .A1(\tms1x00.O_pla_ands[20][4] ),
    .S(_03370_),
    .X(_00051_));
 sky130_fd_sc_hd__mux2_1 _06930_ (.A0(net1040),
    .A1(\tms1x00.O_pla_ands[20][5] ),
    .S(_03370_),
    .X(_00052_));
 sky130_fd_sc_hd__mux2_1 _06931_ (.A0(net1031),
    .A1(\tms1x00.O_pla_ands[20][6] ),
    .S(_03370_),
    .X(_00053_));
 sky130_fd_sc_hd__mux2_1 _06932_ (.A0(net1025),
    .A1(\tms1x00.O_pla_ands[20][7] ),
    .S(_03370_),
    .X(_00054_));
 sky130_fd_sc_hd__mux2_1 _06933_ (.A0(net1017),
    .A1(\tms1x00.O_pla_ands[20][8] ),
    .S(_03370_),
    .X(_00055_));
 sky130_fd_sc_hd__mux2_1 _06934_ (.A0(net1009),
    .A1(\tms1x00.O_pla_ands[20][9] ),
    .S(_03370_),
    .X(_00056_));
 sky130_fd_sc_hd__xnor2_4 _06935_ (.A(\tms1x00.wb_step ),
    .B(\tms1x00.wb_step_state ),
    .Y(_03371_));
 sky130_fd_sc_hd__and2_4 _06936_ (.A(net145),
    .B(_03371_),
    .X(_03372_));
 sky130_fd_sc_hd__nand2_8 _06937_ (.A(net145),
    .B(_03371_),
    .Y(_03373_));
 sky130_fd_sc_hd__nor2_8 _06938_ (.A(net591),
    .B(_03372_),
    .Y(_03374_));
 sky130_fd_sc_hd__or2_2 _06939_ (.A(net698),
    .B(net702),
    .X(_03375_));
 sky130_fd_sc_hd__nand2_4 _06940_ (.A(net688),
    .B(net693),
    .Y(_03376_));
 sky130_fd_sc_hd__and4_4 _06941_ (.A(_01623_),
    .B(_01624_),
    .C(_01625_),
    .D(_01626_),
    .X(_03377_));
 sky130_fd_sc_hd__or4_4 _06942_ (.A(net671),
    .B(net675),
    .C(\tms1x00.ins_arg[2] ),
    .D(net684),
    .X(_03378_));
 sky130_fd_sc_hd__and2b_2 _06943_ (.A_N(_02011_),
    .B(_03376_),
    .X(_03379_));
 sky130_fd_sc_hd__inv_2 _06944_ (.A(_03379_),
    .Y(_03380_));
 sky130_fd_sc_hd__or3_1 _06945_ (.A(\tms1x00.ins_arg[2] ),
    .B(net684),
    .C(net688),
    .X(_03381_));
 sky130_fd_sc_hd__a21o_4 _06946_ (.A1(_01624_),
    .A2(_03381_),
    .B1(net671),
    .X(_03382_));
 sky130_fd_sc_hd__a22o_1 _06947_ (.A1(\tms1x00.K_latch[0] ),
    .A2(_03377_),
    .B1(_03379_),
    .B2(_03375_),
    .X(_03383_));
 sky130_fd_sc_hd__mux2_4 _06948_ (.A0(net688),
    .A1(_03383_),
    .S(_03382_),
    .X(_03384_));
 sky130_fd_sc_hd__mux2_1 _06949_ (.A0(_01628_),
    .A1(net6),
    .S(_03375_),
    .X(_03385_));
 sky130_fd_sc_hd__and2_1 _06950_ (.A(_02012_),
    .B(_03385_),
    .X(_03386_));
 sky130_fd_sc_hd__a221o_4 _06951_ (.A1(\tms1x00.A[0] ),
    .A2(_02009_),
    .B1(_03384_),
    .B2(_01991_),
    .C1(_03386_),
    .X(_03387_));
 sky130_fd_sc_hd__mux2_1 _06952_ (.A0(net153),
    .A1(_03387_),
    .S(_03374_),
    .X(_00057_));
 sky130_fd_sc_hd__nor2_2 _06953_ (.A(_01629_),
    .B(net702),
    .Y(_03388_));
 sky130_fd_sc_hd__a2bb2o_1 _06954_ (.A1_N(_03380_),
    .A2_N(_03388_),
    .B1(\tms1x00.K_latch[1] ),
    .B2(_03377_),
    .X(_03389_));
 sky130_fd_sc_hd__mux2_4 _06955_ (.A0(net693),
    .A1(_03389_),
    .S(_03382_),
    .X(_03390_));
 sky130_fd_sc_hd__nand2_1 _06956_ (.A(net693),
    .B(_03388_),
    .Y(_03391_));
 sky130_fd_sc_hd__o211a_1 _06957_ (.A1(net7),
    .A2(_03388_),
    .B1(_03391_),
    .C1(_02012_),
    .X(_03392_));
 sky130_fd_sc_hd__a221o_4 _06958_ (.A1(\tms1x00.A[1] ),
    .A2(_02009_),
    .B1(_03390_),
    .B2(_01991_),
    .C1(_03392_),
    .X(_03393_));
 sky130_fd_sc_hd__mux2_1 _06959_ (.A0(net154),
    .A1(_03393_),
    .S(_03374_),
    .X(_00058_));
 sky130_fd_sc_hd__nand2_4 _06960_ (.A(_01629_),
    .B(net702),
    .Y(_03394_));
 sky130_fd_sc_hd__a22o_1 _06961_ (.A1(\tms1x00.K_latch[2] ),
    .A2(_03377_),
    .B1(_03379_),
    .B2(_03394_),
    .X(_03395_));
 sky130_fd_sc_hd__mux2_4 _06962_ (.A0(net699),
    .A1(_03395_),
    .S(_03382_),
    .X(_03396_));
 sky130_fd_sc_hd__mux2_1 _06963_ (.A0(_01628_),
    .A1(net8),
    .S(_03394_),
    .X(_03397_));
 sky130_fd_sc_hd__a22o_1 _06964_ (.A1(_01991_),
    .A2(_03396_),
    .B1(_03397_),
    .B2(_02012_),
    .X(_03398_));
 sky130_fd_sc_hd__a21o_2 _06965_ (.A1(\tms1x00.A[2] ),
    .A2(_02009_),
    .B1(_03398_),
    .X(_03399_));
 sky130_fd_sc_hd__mux2_1 _06966_ (.A0(net155),
    .A1(_03399_),
    .S(_03374_),
    .X(_00059_));
 sky130_fd_sc_hd__nand2_4 _06967_ (.A(net699),
    .B(net702),
    .Y(_03400_));
 sky130_fd_sc_hd__a22o_1 _06968_ (.A1(\tms1x00.K_latch[3] ),
    .A2(_03377_),
    .B1(_03379_),
    .B2(_03400_),
    .X(_03401_));
 sky130_fd_sc_hd__mux2_4 _06969_ (.A0(net702),
    .A1(_03401_),
    .S(_03382_),
    .X(_03402_));
 sky130_fd_sc_hd__and2_1 _06970_ (.A(net9),
    .B(_03400_),
    .X(_03403_));
 sky130_fd_sc_hd__nor2_1 _06971_ (.A(net693),
    .B(_03400_),
    .Y(_03404_));
 sky130_fd_sc_hd__o21a_1 _06972_ (.A1(_03403_),
    .A2(_03404_),
    .B1(_02012_),
    .X(_03405_));
 sky130_fd_sc_hd__a221o_4 _06973_ (.A1(\tms1x00.A[3] ),
    .A2(_02009_),
    .B1(_03402_),
    .B2(_01991_),
    .C1(_03405_),
    .X(_03406_));
 sky130_fd_sc_hd__mux2_1 _06974_ (.A0(net156),
    .A1(_03406_),
    .S(_03374_),
    .X(_00060_));
 sky130_fd_sc_hd__and3_4 _06975_ (.A(net874),
    .B(net598),
    .C(net359),
    .X(_03407_));
 sky130_fd_sc_hd__or3_4 _06976_ (.A(net858),
    .B(_03353_),
    .C(net357),
    .X(_03408_));
 sky130_fd_sc_hd__or2_1 _06977_ (.A(\tms1x00.O_pla_ands[19][0] ),
    .B(_03407_),
    .X(_03409_));
 sky130_fd_sc_hd__o211a_1 _06978_ (.A1(net977),
    .A2(_03408_),
    .B1(_03409_),
    .C1(net473),
    .X(_00061_));
 sky130_fd_sc_hd__or2_1 _06979_ (.A(\tms1x00.O_pla_ands[19][1] ),
    .B(_03407_),
    .X(_03410_));
 sky130_fd_sc_hd__o211a_1 _06980_ (.A1(net929),
    .A2(_03408_),
    .B1(_03410_),
    .C1(net473),
    .X(_00062_));
 sky130_fd_sc_hd__or2_1 _06981_ (.A(\tms1x00.O_pla_ands[19][2] ),
    .B(_03407_),
    .X(_03411_));
 sky130_fd_sc_hd__o211a_1 _06982_ (.A1(net1064),
    .A2(_03408_),
    .B1(_03411_),
    .C1(net474),
    .X(_00063_));
 sky130_fd_sc_hd__or2_1 _06983_ (.A(\tms1x00.O_pla_ands[19][3] ),
    .B(_03407_),
    .X(_03412_));
 sky130_fd_sc_hd__o211a_1 _06984_ (.A1(net1056),
    .A2(_03408_),
    .B1(_03412_),
    .C1(net473),
    .X(_00064_));
 sky130_fd_sc_hd__or2_1 _06985_ (.A(\tms1x00.O_pla_ands[19][4] ),
    .B(_03407_),
    .X(_03413_));
 sky130_fd_sc_hd__o211a_1 _06986_ (.A1(net1048),
    .A2(_03408_),
    .B1(_03413_),
    .C1(net474),
    .X(_00065_));
 sky130_fd_sc_hd__or2_1 _06987_ (.A(\tms1x00.O_pla_ands[19][5] ),
    .B(_03407_),
    .X(_03414_));
 sky130_fd_sc_hd__o211a_1 _06988_ (.A1(net1040),
    .A2(_03408_),
    .B1(_03414_),
    .C1(net474),
    .X(_00066_));
 sky130_fd_sc_hd__or2_1 _06989_ (.A(\tms1x00.O_pla_ands[19][6] ),
    .B(_03407_),
    .X(_03415_));
 sky130_fd_sc_hd__o211a_1 _06990_ (.A1(net1031),
    .A2(_03408_),
    .B1(_03415_),
    .C1(net473),
    .X(_00067_));
 sky130_fd_sc_hd__a21o_1 _06991_ (.A1(net1025),
    .A2(_03407_),
    .B1(net534),
    .X(_03416_));
 sky130_fd_sc_hd__a21o_1 _06992_ (.A1(\tms1x00.O_pla_ands[19][7] ),
    .A2(_03408_),
    .B1(_03416_),
    .X(_00068_));
 sky130_fd_sc_hd__a21o_1 _06993_ (.A1(net1017),
    .A2(_03407_),
    .B1(net534),
    .X(_03417_));
 sky130_fd_sc_hd__a21o_1 _06994_ (.A1(\tms1x00.O_pla_ands[19][8] ),
    .A2(_03408_),
    .B1(_03417_),
    .X(_00069_));
 sky130_fd_sc_hd__or2_1 _06995_ (.A(\tms1x00.O_pla_ands[19][9] ),
    .B(_03407_),
    .X(_03418_));
 sky130_fd_sc_hd__o211a_1 _06996_ (.A1(net1009),
    .A2(_03408_),
    .B1(_03418_),
    .C1(net474),
    .X(_00070_));
 sky130_fd_sc_hd__nand4_1 _06997_ (.A(net996),
    .B(net600),
    .C(_03347_),
    .D(_03349_),
    .Y(_03419_));
 sky130_fd_sc_hd__nor2_8 _06998_ (.A(net799),
    .B(net356),
    .Y(_03420_));
 sky130_fd_sc_hd__or2_4 _06999_ (.A(net807),
    .B(net356),
    .X(_03421_));
 sky130_fd_sc_hd__nor2_4 _07000_ (.A(net519),
    .B(_03420_),
    .Y(_03422_));
 sky130_fd_sc_hd__nand2_4 _07001_ (.A(net481),
    .B(_03421_),
    .Y(_03423_));
 sky130_fd_sc_hd__and2_2 _07002_ (.A(net930),
    .B(net462),
    .X(_03424_));
 sky130_fd_sc_hd__nor2_2 _07003_ (.A(net705),
    .B(net491),
    .Y(_03425_));
 sky130_fd_sc_hd__nand2_4 _07004_ (.A(_01638_),
    .B(net557),
    .Y(_03426_));
 sky130_fd_sc_hd__or2_4 _07005_ (.A(net397),
    .B(net396),
    .X(_03427_));
 sky130_fd_sc_hd__mux2_1 _07006_ (.A0(\tms1x00.ins_pla_ors[12][1] ),
    .A1(net354),
    .S(net234),
    .X(_00071_));
 sky130_fd_sc_hd__and2_4 _07007_ (.A(net1066),
    .B(net461),
    .X(_03428_));
 sky130_fd_sc_hd__or2_4 _07008_ (.A(net390),
    .B(_03428_),
    .X(_03429_));
 sky130_fd_sc_hd__mux2_1 _07009_ (.A0(\tms1x00.ins_pla_ors[12][2] ),
    .A1(_03429_),
    .S(net234),
    .X(_00072_));
 sky130_fd_sc_hd__and2_4 _07010_ (.A(net1058),
    .B(net461),
    .X(_03430_));
 sky130_fd_sc_hd__nor2_4 _07011_ (.A(_01638_),
    .B(net490),
    .Y(_03431_));
 sky130_fd_sc_hd__nand2_8 _07012_ (.A(net705),
    .B(net535),
    .Y(_03432_));
 sky130_fd_sc_hd__or2_4 _07013_ (.A(_03430_),
    .B(net374),
    .X(_03433_));
 sky130_fd_sc_hd__mux2_1 _07014_ (.A0(\tms1x00.ins_pla_ors[12][3] ),
    .A1(_03433_),
    .S(net234),
    .X(_00073_));
 sky130_fd_sc_hd__and2_4 _07015_ (.A(net1033),
    .B(net462),
    .X(_03434_));
 sky130_fd_sc_hd__or2_4 _07016_ (.A(net392),
    .B(_03434_),
    .X(_03435_));
 sky130_fd_sc_hd__mux2_1 _07017_ (.A0(\tms1x00.ins_pla_ors[12][6] ),
    .A1(_03435_),
    .S(net234),
    .X(_00074_));
 sky130_fd_sc_hd__and2_1 _07018_ (.A(net1026),
    .B(net478),
    .X(_03436_));
 sky130_fd_sc_hd__or2_4 _07019_ (.A(net391),
    .B(net368),
    .X(_03437_));
 sky130_fd_sc_hd__mux2_1 _07020_ (.A0(\tms1x00.ins_pla_ors[12][7] ),
    .A1(_03437_),
    .S(net234),
    .X(_00075_));
 sky130_fd_sc_hd__and2_4 _07021_ (.A(net1018),
    .B(net462),
    .X(_03438_));
 sky130_fd_sc_hd__or2_4 _07022_ (.A(net389),
    .B(_03438_),
    .X(_03439_));
 sky130_fd_sc_hd__mux2_1 _07023_ (.A0(\tms1x00.ins_pla_ors[12][8] ),
    .A1(net353),
    .S(net234),
    .X(_00076_));
 sky130_fd_sc_hd__a221o_1 _07024_ (.A1(net953),
    .A2(_03420_),
    .B1(_03422_),
    .B2(\tms1x00.ins_pla_ors[12][14] ),
    .C1(net375),
    .X(_00077_));
 sky130_fd_sc_hd__or2_1 _07025_ (.A(net942),
    .B(net541),
    .X(_03440_));
 sky130_fd_sc_hd__and2_2 _07026_ (.A(net385),
    .B(_03440_),
    .X(_03441_));
 sky130_fd_sc_hd__mux2_1 _07027_ (.A0(\tms1x00.ins_pla_ors[12][16] ),
    .A1(_03441_),
    .S(net234),
    .X(_00078_));
 sky130_fd_sc_hd__and2_1 _07028_ (.A(net940),
    .B(net480),
    .X(_03442_));
 sky130_fd_sc_hd__or2_1 _07029_ (.A(net381),
    .B(_03442_),
    .X(_03443_));
 sky130_fd_sc_hd__mux2_1 _07030_ (.A0(\tms1x00.ins_pla_ors[12][17] ),
    .A1(_03443_),
    .S(_03423_),
    .X(_00079_));
 sky130_fd_sc_hd__or2_4 _07031_ (.A(net938),
    .B(net541),
    .X(_03444_));
 sky130_fd_sc_hd__a22o_1 _07032_ (.A1(\tms1x00.ins_pla_ors[12][18] ),
    .A2(net338),
    .B1(net234),
    .B2(_03444_),
    .X(_03445_));
 sky130_fd_sc_hd__and2_1 _07033_ (.A(net385),
    .B(_03445_),
    .X(_00080_));
 sky130_fd_sc_hd__and2_1 _07034_ (.A(net1077),
    .B(net462),
    .X(_03446_));
 sky130_fd_sc_hd__a221o_1 _07035_ (.A1(\tms1x00.ins_pla_ors[12][21] ),
    .A2(_03422_),
    .B1(_03446_),
    .B2(_03420_),
    .C1(net389),
    .X(_00081_));
 sky130_fd_sc_hd__or2_4 _07036_ (.A(net1072),
    .B(net539),
    .X(_03447_));
 sky130_fd_sc_hd__and2_1 _07037_ (.A(net385),
    .B(_03447_),
    .X(_03448_));
 sky130_fd_sc_hd__mux2_1 _07038_ (.A0(\tms1x00.ins_pla_ors[12][26] ),
    .A1(_03448_),
    .S(net234),
    .X(_00082_));
 sky130_fd_sc_hd__and2_4 _07039_ (.A(net108),
    .B(net480),
    .X(_03449_));
 sky130_fd_sc_hd__or2_4 _07040_ (.A(net393),
    .B(_03449_),
    .X(_03450_));
 sky130_fd_sc_hd__mux2_1 _07041_ (.A0(\tms1x00.ins_pla_ors[12][28] ),
    .A1(_03450_),
    .S(_03423_),
    .X(_00083_));
 sky130_fd_sc_hd__and2_2 _07042_ (.A(net109),
    .B(net481),
    .X(_03451_));
 sky130_fd_sc_hd__or2_4 _07043_ (.A(net395),
    .B(_03451_),
    .X(_03452_));
 sky130_fd_sc_hd__mux2_1 _07044_ (.A0(\tms1x00.ins_pla_ors[12][29] ),
    .A1(_03452_),
    .S(_03423_),
    .X(_00084_));
 sky130_fd_sc_hd__nor2_4 _07045_ (.A(net605),
    .B(net355),
    .Y(_03453_));
 sky130_fd_sc_hd__or2_4 _07046_ (.A(net605),
    .B(net355),
    .X(_03454_));
 sky130_fd_sc_hd__nor2_1 _07047_ (.A(net522),
    .B(net337),
    .Y(_03455_));
 sky130_fd_sc_hd__and2_4 _07048_ (.A(net979),
    .B(net461),
    .X(_03456_));
 sky130_fd_sc_hd__o22a_1 _07049_ (.A1(\tms1x00.ins_pla_ors[14][0] ),
    .A2(net337),
    .B1(net231),
    .B2(_03456_),
    .X(_00085_));
 sky130_fd_sc_hd__o22a_1 _07050_ (.A1(\tms1x00.ins_pla_ors[14][1] ),
    .A2(net337),
    .B1(net233),
    .B2(net397),
    .X(_00086_));
 sky130_fd_sc_hd__o22a_1 _07051_ (.A1(\tms1x00.ins_pla_ors[14][3] ),
    .A2(net337),
    .B1(net231),
    .B2(_03430_),
    .X(_00087_));
 sky130_fd_sc_hd__and2_4 _07052_ (.A(net1041),
    .B(net461),
    .X(_03457_));
 sky130_fd_sc_hd__o22a_1 _07053_ (.A1(\tms1x00.ins_pla_ors[14][5] ),
    .A2(net336),
    .B1(net232),
    .B2(net366),
    .X(_00088_));
 sky130_fd_sc_hd__o22a_1 _07054_ (.A1(\tms1x00.ins_pla_ors[14][6] ),
    .A2(net336),
    .B1(net232),
    .B2(_03434_),
    .X(_00089_));
 sky130_fd_sc_hd__o22a_1 _07055_ (.A1(\tms1x00.ins_pla_ors[14][7] ),
    .A2(net337),
    .B1(net231),
    .B2(net367),
    .X(_00090_));
 sky130_fd_sc_hd__o22a_1 _07056_ (.A1(\tms1x00.ins_pla_ors[14][8] ),
    .A2(net337),
    .B1(net231),
    .B2(_03438_),
    .X(_00091_));
 sky130_fd_sc_hd__and2_2 _07057_ (.A(net1010),
    .B(net462),
    .X(_03458_));
 sky130_fd_sc_hd__o22a_1 _07058_ (.A1(\tms1x00.ins_pla_ors[14][9] ),
    .A2(net337),
    .B1(net231),
    .B2(net365),
    .X(_00092_));
 sky130_fd_sc_hd__and2_4 _07059_ (.A(net972),
    .B(net461),
    .X(_03459_));
 sky130_fd_sc_hd__o22a_1 _07060_ (.A1(\tms1x00.ins_pla_ors[14][10] ),
    .A2(net337),
    .B1(net231),
    .B2(_03459_),
    .X(_00093_));
 sky130_fd_sc_hd__and2_4 _07061_ (.A(net968),
    .B(net461),
    .X(_03460_));
 sky130_fd_sc_hd__o22a_1 _07062_ (.A1(\tms1x00.ins_pla_ors[14][11] ),
    .A2(net337),
    .B1(net231),
    .B2(_03460_),
    .X(_00094_));
 sky130_fd_sc_hd__mux2_1 _07063_ (.A0(net953),
    .A1(\tms1x00.ins_pla_ors[14][14] ),
    .S(_03454_),
    .X(_03461_));
 sky130_fd_sc_hd__or2_1 _07064_ (.A(net520),
    .B(_03461_),
    .X(_00095_));
 sky130_fd_sc_hd__or2_1 _07065_ (.A(\tms1x00.ins_pla_ors[14][15] ),
    .B(net336),
    .X(_03462_));
 sky130_fd_sc_hd__o211a_1 _07066_ (.A1(net948),
    .A2(_03454_),
    .B1(_03462_),
    .C1(net479),
    .X(_00096_));
 sky130_fd_sc_hd__o22a_1 _07067_ (.A1(\tms1x00.ins_pla_ors[14][17] ),
    .A2(net336),
    .B1(net232),
    .B2(_03442_),
    .X(_00097_));
 sky130_fd_sc_hd__or2_1 _07068_ (.A(\tms1x00.ins_pla_ors[14][18] ),
    .B(net336),
    .X(_03463_));
 sky130_fd_sc_hd__o211a_1 _07069_ (.A1(net938),
    .A2(_03454_),
    .B1(_03463_),
    .C1(net479),
    .X(_00098_));
 sky130_fd_sc_hd__and2_1 _07070_ (.A(net937),
    .B(net462),
    .X(_03464_));
 sky130_fd_sc_hd__o22a_1 _07071_ (.A1(\tms1x00.ins_pla_ors[14][19] ),
    .A2(net337),
    .B1(net233),
    .B2(_03464_),
    .X(_00099_));
 sky130_fd_sc_hd__or2_1 _07072_ (.A(\tms1x00.ins_pla_ors[14][20] ),
    .B(net336),
    .X(_03465_));
 sky130_fd_sc_hd__o211a_1 _07073_ (.A1(net1078),
    .A2(_03454_),
    .B1(_03465_),
    .C1(net480),
    .X(_00100_));
 sky130_fd_sc_hd__mux2_1 _07074_ (.A0(net1077),
    .A1(\tms1x00.ins_pla_ors[14][21] ),
    .S(_03454_),
    .X(_03466_));
 sky130_fd_sc_hd__or2_1 _07075_ (.A(net520),
    .B(_03466_),
    .X(_00101_));
 sky130_fd_sc_hd__and2_4 _07076_ (.A(net1073),
    .B(net481),
    .X(_03467_));
 sky130_fd_sc_hd__o22a_1 _07077_ (.A1(\tms1x00.ins_pla_ors[14][24] ),
    .A2(_03453_),
    .B1(net232),
    .B2(_03467_),
    .X(_00102_));
 sky130_fd_sc_hd__or2_1 _07078_ (.A(\tms1x00.ins_pla_ors[14][26] ),
    .B(net336),
    .X(_03468_));
 sky130_fd_sc_hd__o211a_1 _07079_ (.A1(net1072),
    .A2(_03454_),
    .B1(_03468_),
    .C1(net479),
    .X(_00103_));
 sky130_fd_sc_hd__o22a_1 _07080_ (.A1(\tms1x00.ins_pla_ors[14][28] ),
    .A2(net336),
    .B1(net232),
    .B2(_03449_),
    .X(_00104_));
 sky130_fd_sc_hd__and3_4 _07081_ (.A(net713),
    .B(_03347_),
    .C(_03349_),
    .X(_03469_));
 sky130_fd_sc_hd__or3_4 _07082_ (.A(net711),
    .B(_03348_),
    .C(_03350_),
    .X(_03470_));
 sky130_fd_sc_hd__nor2_2 _07083_ (.A(net923),
    .B(net911),
    .Y(_03471_));
 sky130_fd_sc_hd__nand2_1 _07084_ (.A(net987),
    .B(net994),
    .Y(_03472_));
 sky130_fd_sc_hd__and3_4 _07085_ (.A(net739),
    .B(net350),
    .C(_03471_),
    .X(_03473_));
 sky130_fd_sc_hd__nor2_4 _07086_ (.A(net522),
    .B(_03473_),
    .Y(_03474_));
 sky130_fd_sc_hd__or2_4 _07087_ (.A(net512),
    .B(_03473_),
    .X(_03475_));
 sky130_fd_sc_hd__or2_4 _07088_ (.A(net374),
    .B(_03456_),
    .X(_03476_));
 sky130_fd_sc_hd__mux2_1 _07089_ (.A0(\tms1x00.ins_pla_ands[26][0] ),
    .A1(_03476_),
    .S(_03475_),
    .X(_00105_));
 sky130_fd_sc_hd__or2_4 _07090_ (.A(_03428_),
    .B(net374),
    .X(_03477_));
 sky130_fd_sc_hd__mux2_1 _07091_ (.A0(\tms1x00.ins_pla_ands[26][2] ),
    .A1(_03477_),
    .S(_03475_),
    .X(_00106_));
 sky130_fd_sc_hd__and2_4 _07092_ (.A(net1049),
    .B(net461),
    .X(_03478_));
 sky130_fd_sc_hd__or2_4 _07093_ (.A(net374),
    .B(_03478_),
    .X(_03479_));
 sky130_fd_sc_hd__mux2_1 _07094_ (.A0(\tms1x00.ins_pla_ands[26][4] ),
    .A1(_03479_),
    .S(_03475_),
    .X(_00107_));
 sky130_fd_sc_hd__or2_4 _07095_ (.A(net377),
    .B(_03434_),
    .X(_03480_));
 sky130_fd_sc_hd__mux2_1 _07096_ (.A0(\tms1x00.ins_pla_ands[26][6] ),
    .A1(_03480_),
    .S(_03475_),
    .X(_00108_));
 sky130_fd_sc_hd__a221o_1 _07097_ (.A1(_03438_),
    .A2(_03473_),
    .B1(_03474_),
    .B2(\tms1x00.ins_pla_ands[26][8] ),
    .C1(net374),
    .X(_00109_));
 sky130_fd_sc_hd__or2_1 _07098_ (.A(net390),
    .B(net364),
    .X(_03481_));
 sky130_fd_sc_hd__mux2_1 _07099_ (.A0(\tms1x00.ins_pla_ands[26][9] ),
    .A1(_03481_),
    .S(_03475_),
    .X(_00110_));
 sky130_fd_sc_hd__or2_4 _07100_ (.A(net374),
    .B(_03459_),
    .X(_03482_));
 sky130_fd_sc_hd__mux2_1 _07101_ (.A0(\tms1x00.ins_pla_ands[26][10] ),
    .A1(_03482_),
    .S(_03475_),
    .X(_00111_));
 sky130_fd_sc_hd__or2_2 _07102_ (.A(net390),
    .B(_03460_),
    .X(_03483_));
 sky130_fd_sc_hd__mux2_1 _07103_ (.A0(\tms1x00.ins_pla_ands[26][11] ),
    .A1(net347),
    .S(_03475_),
    .X(_00112_));
 sky130_fd_sc_hd__and2_4 _07104_ (.A(net965),
    .B(net461),
    .X(_03484_));
 sky130_fd_sc_hd__or2_4 _07105_ (.A(net374),
    .B(_03484_),
    .X(_03485_));
 sky130_fd_sc_hd__mux2_1 _07106_ (.A0(\tms1x00.ins_pla_ands[26][12] ),
    .A1(_03485_),
    .S(_03475_),
    .X(_00113_));
 sky130_fd_sc_hd__and2_4 _07107_ (.A(net959),
    .B(net462),
    .X(_03486_));
 sky130_fd_sc_hd__or2_4 _07108_ (.A(net389),
    .B(_03486_),
    .X(_03487_));
 sky130_fd_sc_hd__mux2_1 _07109_ (.A0(\tms1x00.ins_pla_ands[26][13] ),
    .A1(_03487_),
    .S(_03475_),
    .X(_00114_));
 sky130_fd_sc_hd__nor2_1 _07110_ (.A(net772),
    .B(net355),
    .Y(_03488_));
 sky130_fd_sc_hd__or2_4 _07111_ (.A(net772),
    .B(net355),
    .X(_03489_));
 sky130_fd_sc_hd__nor2_1 _07112_ (.A(net522),
    .B(net332),
    .Y(_03490_));
 sky130_fd_sc_hd__o22a_1 _07113_ (.A1(\tms1x00.ins_pla_ors[15][0] ),
    .A2(net332),
    .B1(net228),
    .B2(_03456_),
    .X(_00115_));
 sky130_fd_sc_hd__o22a_1 _07114_ (.A1(\tms1x00.ins_pla_ors[15][1] ),
    .A2(net333),
    .B1(net228),
    .B2(_03424_),
    .X(_00116_));
 sky130_fd_sc_hd__o22a_1 _07115_ (.A1(\tms1x00.ins_pla_ors[15][2] ),
    .A2(net333),
    .B1(net229),
    .B2(_03428_),
    .X(_00117_));
 sky130_fd_sc_hd__o22a_1 _07116_ (.A1(\tms1x00.ins_pla_ors[15][3] ),
    .A2(net332),
    .B1(net229),
    .B2(_03430_),
    .X(_00118_));
 sky130_fd_sc_hd__o22a_1 _07117_ (.A1(\tms1x00.ins_pla_ors[15][4] ),
    .A2(net332),
    .B1(net229),
    .B2(_03478_),
    .X(_00119_));
 sky130_fd_sc_hd__o22a_1 _07118_ (.A1(\tms1x00.ins_pla_ors[15][5] ),
    .A2(net333),
    .B1(net228),
    .B2(_03457_),
    .X(_00120_));
 sky130_fd_sc_hd__o22a_1 _07119_ (.A1(\tms1x00.ins_pla_ors[15][6] ),
    .A2(net334),
    .B1(net230),
    .B2(_03434_),
    .X(_00121_));
 sky130_fd_sc_hd__o22a_1 _07120_ (.A1(\tms1x00.ins_pla_ors[15][8] ),
    .A2(net333),
    .B1(net229),
    .B2(_03438_),
    .X(_00122_));
 sky130_fd_sc_hd__o22a_1 _07121_ (.A1(\tms1x00.ins_pla_ors[15][9] ),
    .A2(net332),
    .B1(net228),
    .B2(net365),
    .X(_00123_));
 sky130_fd_sc_hd__o22a_1 _07122_ (.A1(\tms1x00.ins_pla_ors[15][10] ),
    .A2(net332),
    .B1(net228),
    .B2(_03459_),
    .X(_00124_));
 sky130_fd_sc_hd__o22a_1 _07123_ (.A1(\tms1x00.ins_pla_ors[15][11] ),
    .A2(net333),
    .B1(net229),
    .B2(_03460_),
    .X(_00125_));
 sky130_fd_sc_hd__o22a_1 _07124_ (.A1(\tms1x00.ins_pla_ors[15][12] ),
    .A2(net332),
    .B1(net228),
    .B2(_03484_),
    .X(_00126_));
 sky130_fd_sc_hd__o22a_1 _07125_ (.A1(\tms1x00.ins_pla_ors[15][13] ),
    .A2(net332),
    .B1(net228),
    .B2(net363),
    .X(_00127_));
 sky130_fd_sc_hd__or2_1 _07126_ (.A(\tms1x00.ins_pla_ors[15][14] ),
    .B(net332),
    .X(_03491_));
 sky130_fd_sc_hd__o211a_1 _07127_ (.A1(net953),
    .A2(_03489_),
    .B1(_03491_),
    .C1(net462),
    .X(_00128_));
 sky130_fd_sc_hd__or2_1 _07128_ (.A(\tms1x00.ins_pla_ors[15][15] ),
    .B(net334),
    .X(_03492_));
 sky130_fd_sc_hd__o211a_1 _07129_ (.A1(net948),
    .A2(_03489_),
    .B1(_03492_),
    .C1(net479),
    .X(_00129_));
 sky130_fd_sc_hd__or2_1 _07130_ (.A(\tms1x00.ins_pla_ors[15][16] ),
    .B(net334),
    .X(_03493_));
 sky130_fd_sc_hd__o211a_1 _07131_ (.A1(net942),
    .A2(_03489_),
    .B1(_03493_),
    .C1(net480),
    .X(_00130_));
 sky130_fd_sc_hd__o22a_1 _07132_ (.A1(\tms1x00.ins_pla_ors[15][17] ),
    .A2(net335),
    .B1(net230),
    .B2(_03442_),
    .X(_00131_));
 sky130_fd_sc_hd__or2_1 _07133_ (.A(\tms1x00.ins_pla_ors[15][18] ),
    .B(net334),
    .X(_03494_));
 sky130_fd_sc_hd__o211a_1 _07134_ (.A1(net938),
    .A2(_03489_),
    .B1(_03494_),
    .C1(net479),
    .X(_00132_));
 sky130_fd_sc_hd__o22a_1 _07135_ (.A1(\tms1x00.ins_pla_ors[15][19] ),
    .A2(net333),
    .B1(net228),
    .B2(_03464_),
    .X(_00133_));
 sky130_fd_sc_hd__or2_1 _07136_ (.A(\tms1x00.ins_pla_ors[15][20] ),
    .B(net334),
    .X(_03495_));
 sky130_fd_sc_hd__o211a_1 _07137_ (.A1(net1078),
    .A2(_03489_),
    .B1(_03495_),
    .C1(net480),
    .X(_00134_));
 sky130_fd_sc_hd__o22a_1 _07138_ (.A1(\tms1x00.ins_pla_ors[15][21] ),
    .A2(net332),
    .B1(net228),
    .B2(_03446_),
    .X(_00135_));
 sky130_fd_sc_hd__or2_1 _07139_ (.A(\tms1x00.ins_pla_ors[15][22] ),
    .B(net334),
    .X(_03496_));
 sky130_fd_sc_hd__o211a_1 _07140_ (.A1(net1075),
    .A2(_03489_),
    .B1(_03496_),
    .C1(net479),
    .X(_00136_));
 sky130_fd_sc_hd__and2_2 _07141_ (.A(net1074),
    .B(net479),
    .X(_03497_));
 sky130_fd_sc_hd__o22a_1 _07142_ (.A1(\tms1x00.ins_pla_ors[15][23] ),
    .A2(net334),
    .B1(net230),
    .B2(_03497_),
    .X(_00137_));
 sky130_fd_sc_hd__and2_4 _07143_ (.A(net105),
    .B(net480),
    .X(_03498_));
 sky130_fd_sc_hd__o22a_1 _07144_ (.A1(\tms1x00.ins_pla_ors[15][25] ),
    .A2(net334),
    .B1(net230),
    .B2(_03498_),
    .X(_00138_));
 sky130_fd_sc_hd__or2_1 _07145_ (.A(\tms1x00.ins_pla_ors[15][26] ),
    .B(net334),
    .X(_03499_));
 sky130_fd_sc_hd__o211a_1 _07146_ (.A1(net1072),
    .A2(_03489_),
    .B1(_03499_),
    .C1(net479),
    .X(_00139_));
 sky130_fd_sc_hd__and2_4 _07147_ (.A(net107),
    .B(net480),
    .X(_03500_));
 sky130_fd_sc_hd__o22a_1 _07148_ (.A1(\tms1x00.ins_pla_ors[15][27] ),
    .A2(net335),
    .B1(net230),
    .B2(_03500_),
    .X(_00140_));
 sky130_fd_sc_hd__o22a_1 _07149_ (.A1(\tms1x00.ins_pla_ors[15][28] ),
    .A2(net334),
    .B1(net230),
    .B2(_03449_),
    .X(_00141_));
 sky130_fd_sc_hd__o22a_1 _07150_ (.A1(\tms1x00.ins_pla_ors[15][29] ),
    .A2(net335),
    .B1(net230),
    .B2(_03451_),
    .X(_00142_));
 sky130_fd_sc_hd__nand4_4 _07151_ (.A(net913),
    .B(net600),
    .C(_03347_),
    .D(_03349_),
    .Y(_03501_));
 sky130_fd_sc_hd__nor2_8 _07152_ (.A(net810),
    .B(net345),
    .Y(_03502_));
 sky130_fd_sc_hd__or2_4 _07153_ (.A(net809),
    .B(net345),
    .X(_03503_));
 sky130_fd_sc_hd__mux2_1 _07154_ (.A0(net982),
    .A1(\tms1x00.ins_pla_ors[4][0] ),
    .S(net331),
    .X(_03504_));
 sky130_fd_sc_hd__or2_1 _07155_ (.A(net552),
    .B(_03504_),
    .X(_00143_));
 sky130_fd_sc_hd__mux2_1 _07156_ (.A0(net934),
    .A1(\tms1x00.ins_pla_ors[4][1] ),
    .S(net330),
    .X(_03505_));
 sky130_fd_sc_hd__or2_1 _07157_ (.A(net541),
    .B(_03505_),
    .X(_00144_));
 sky130_fd_sc_hd__mux2_1 _07158_ (.A0(net1070),
    .A1(\tms1x00.ins_pla_ors[4][2] ),
    .S(net331),
    .X(_03506_));
 sky130_fd_sc_hd__or2_1 _07159_ (.A(net554),
    .B(_03506_),
    .X(_00145_));
 sky130_fd_sc_hd__mux2_1 _07160_ (.A0(net1062),
    .A1(\tms1x00.ins_pla_ors[4][3] ),
    .S(net330),
    .X(_03507_));
 sky130_fd_sc_hd__or2_1 _07161_ (.A(net542),
    .B(_03507_),
    .X(_00146_));
 sky130_fd_sc_hd__mux2_1 _07162_ (.A0(net1053),
    .A1(\tms1x00.ins_pla_ors[4][4] ),
    .S(net330),
    .X(_03508_));
 sky130_fd_sc_hd__or2_1 _07163_ (.A(net542),
    .B(_03508_),
    .X(_00147_));
 sky130_fd_sc_hd__mux2_1 _07164_ (.A0(net1029),
    .A1(\tms1x00.ins_pla_ors[4][7] ),
    .S(net331),
    .X(_03509_));
 sky130_fd_sc_hd__or2_1 _07165_ (.A(net554),
    .B(_03509_),
    .X(_00148_));
 sky130_fd_sc_hd__or2_1 _07166_ (.A(\tms1x00.ins_pla_ors[4][9] ),
    .B(_03502_),
    .X(_03510_));
 sky130_fd_sc_hd__o211a_1 _07167_ (.A1(net1013),
    .A2(net331),
    .B1(_03510_),
    .C1(net487),
    .X(_00149_));
 sky130_fd_sc_hd__mux2_1 _07168_ (.A0(net975),
    .A1(\tms1x00.ins_pla_ors[4][10] ),
    .S(net331),
    .X(_03511_));
 sky130_fd_sc_hd__or2_1 _07169_ (.A(net552),
    .B(_03511_),
    .X(_00150_));
 sky130_fd_sc_hd__mux2_1 _07170_ (.A0(net966),
    .A1(\tms1x00.ins_pla_ors[4][12] ),
    .S(net330),
    .X(_03512_));
 sky130_fd_sc_hd__or2_1 _07171_ (.A(net544),
    .B(_03512_),
    .X(_00151_));
 sky130_fd_sc_hd__mux2_1 _07172_ (.A0(net961),
    .A1(\tms1x00.ins_pla_ors[4][13] ),
    .S(net331),
    .X(_03513_));
 sky130_fd_sc_hd__or2_1 _07173_ (.A(net542),
    .B(_03513_),
    .X(_00152_));
 sky130_fd_sc_hd__or2_1 _07174_ (.A(\tms1x00.ins_pla_ors[4][15] ),
    .B(_03502_),
    .X(_03514_));
 sky130_fd_sc_hd__o211a_1 _07175_ (.A1(net948),
    .A2(net330),
    .B1(_03514_),
    .C1(net482),
    .X(_00153_));
 sky130_fd_sc_hd__or2_1 _07176_ (.A(\tms1x00.ins_pla_ors[4][19] ),
    .B(_03502_),
    .X(_03515_));
 sky130_fd_sc_hd__o211a_1 _07177_ (.A1(net935),
    .A2(net331),
    .B1(_03515_),
    .C1(net487),
    .X(_00154_));
 sky130_fd_sc_hd__or2_1 _07178_ (.A(\tms1x00.ins_pla_ors[4][20] ),
    .B(_03502_),
    .X(_03516_));
 sky130_fd_sc_hd__o211a_1 _07179_ (.A1(net1078),
    .A2(_03503_),
    .B1(_03516_),
    .C1(net483),
    .X(_00155_));
 sky130_fd_sc_hd__mux2_1 _07180_ (.A0(net1077),
    .A1(\tms1x00.ins_pla_ors[4][21] ),
    .S(_03503_),
    .X(_03517_));
 sky130_fd_sc_hd__or2_1 _07181_ (.A(net545),
    .B(_03517_),
    .X(_00156_));
 sky130_fd_sc_hd__mux2_1 _07182_ (.A0(net1075),
    .A1(\tms1x00.ins_pla_ors[4][22] ),
    .S(net330),
    .X(_03518_));
 sky130_fd_sc_hd__or2_1 _07183_ (.A(net538),
    .B(_03518_),
    .X(_00157_));
 sky130_fd_sc_hd__or2_1 _07184_ (.A(\tms1x00.ins_pla_ors[4][23] ),
    .B(_03502_),
    .X(_03519_));
 sky130_fd_sc_hd__o211a_1 _07185_ (.A1(net1074),
    .A2(net331),
    .B1(_03519_),
    .C1(net487),
    .X(_00158_));
 sky130_fd_sc_hd__mux2_1 _07186_ (.A0(_03437_),
    .A1(\tms1x00.ins_pla_ors[15][7] ),
    .S(net228),
    .X(_00159_));
 sky130_fd_sc_hd__or2_1 _07187_ (.A(net381),
    .B(_03467_),
    .X(_03520_));
 sky130_fd_sc_hd__mux2_1 _07188_ (.A0(_03520_),
    .A1(\tms1x00.ins_pla_ors[15][24] ),
    .S(net230),
    .X(_00160_));
 sky130_fd_sc_hd__nor2_8 _07189_ (.A(net827),
    .B(net355),
    .Y(_03521_));
 sky130_fd_sc_hd__or2_1 _07190_ (.A(net827),
    .B(net355),
    .X(_03522_));
 sky130_fd_sc_hd__nor2_8 _07191_ (.A(net375),
    .B(_03521_),
    .Y(_03523_));
 sky130_fd_sc_hd__inv_2 _07192_ (.A(_03523_),
    .Y(_03524_));
 sky130_fd_sc_hd__a221o_1 _07193_ (.A1(_03484_),
    .A2(_03521_),
    .B1(_03523_),
    .B2(\tms1x00.ins_pla_ors[8][12] ),
    .C1(net389),
    .X(_00161_));
 sky130_fd_sc_hd__o221a_1 _07194_ (.A1(net960),
    .A2(net327),
    .B1(_03524_),
    .B2(\tms1x00.ins_pla_ors[8][13] ),
    .C1(net384),
    .X(_00162_));
 sky130_fd_sc_hd__mux2_1 _07195_ (.A0(net948),
    .A1(\tms1x00.ins_pla_ors[8][15] ),
    .S(net328),
    .X(_03525_));
 sky130_fd_sc_hd__a21o_1 _07196_ (.A1(net479),
    .A2(_03525_),
    .B1(net374),
    .X(_00163_));
 sky130_fd_sc_hd__a221o_1 _07197_ (.A1(net937),
    .A2(_03521_),
    .B1(_03523_),
    .B2(\tms1x00.ins_pla_ors[8][19] ),
    .C1(net389),
    .X(_00164_));
 sky130_fd_sc_hd__a221o_1 _07198_ (.A1(net1075),
    .A2(_03521_),
    .B1(_03523_),
    .B2(\tms1x00.ins_pla_ors[8][22] ),
    .C1(net393),
    .X(_00165_));
 sky130_fd_sc_hd__a221o_1 _07199_ (.A1(net107),
    .A2(_03521_),
    .B1(_03523_),
    .B2(\tms1x00.ins_pla_ors[8][27] ),
    .C1(net393),
    .X(_00166_));
 sky130_fd_sc_hd__a221o_1 _07200_ (.A1(net108),
    .A2(_03521_),
    .B1(_03523_),
    .B2(\tms1x00.ins_pla_ors[8][28] ),
    .C1(net393),
    .X(_00167_));
 sky130_fd_sc_hd__a221o_1 _07201_ (.A1(net109),
    .A2(_03521_),
    .B1(_03523_),
    .B2(\tms1x00.ins_pla_ors[8][29] ),
    .C1(net393),
    .X(_00168_));
 sky130_fd_sc_hd__nor2_4 _07202_ (.A(net880),
    .B(net355),
    .Y(_03526_));
 sky130_fd_sc_hd__or2_4 _07203_ (.A(net888),
    .B(net356),
    .X(_03527_));
 sky130_fd_sc_hd__nor2_8 _07204_ (.A(net519),
    .B(net325),
    .Y(_03528_));
 sky130_fd_sc_hd__nand2_2 _07205_ (.A(net481),
    .B(_03527_),
    .Y(_03529_));
 sky130_fd_sc_hd__o22a_1 _07206_ (.A1(net982),
    .A2(_03527_),
    .B1(net225),
    .B2(\tms1x00.ins_pla_ors[13][0] ),
    .X(_00169_));
 sky130_fd_sc_hd__o22a_1 _07207_ (.A1(net1022),
    .A2(_03527_),
    .B1(net225),
    .B2(\tms1x00.ins_pla_ors[13][8] ),
    .X(_00170_));
 sky130_fd_sc_hd__a22o_1 _07208_ (.A1(net1010),
    .A2(net325),
    .B1(net227),
    .B2(\tms1x00.ins_pla_ors[13][9] ),
    .X(_00171_));
 sky130_fd_sc_hd__o22a_1 _07209_ (.A1(net968),
    .A2(_03527_),
    .B1(net225),
    .B2(\tms1x00.ins_pla_ors[13][11] ),
    .X(_00172_));
 sky130_fd_sc_hd__a22o_1 _07210_ (.A1(net953),
    .A2(net325),
    .B1(net227),
    .B2(\tms1x00.ins_pla_ors[13][14] ),
    .X(_00173_));
 sky130_fd_sc_hd__or2_1 _07211_ (.A(net948),
    .B(net521),
    .X(_03530_));
 sky130_fd_sc_hd__o22a_1 _07212_ (.A1(net948),
    .A2(_03527_),
    .B1(net225),
    .B2(\tms1x00.ins_pla_ors[13][15] ),
    .X(_00174_));
 sky130_fd_sc_hd__a22o_1 _07213_ (.A1(net942),
    .A2(net325),
    .B1(net227),
    .B2(\tms1x00.ins_pla_ors[13][16] ),
    .X(_00175_));
 sky130_fd_sc_hd__o22a_1 _07214_ (.A1(net938),
    .A2(_03527_),
    .B1(net226),
    .B2(\tms1x00.ins_pla_ors[13][18] ),
    .X(_00176_));
 sky130_fd_sc_hd__o22a_1 _07215_ (.A1(net1078),
    .A2(_03527_),
    .B1(net226),
    .B2(\tms1x00.ins_pla_ors[13][20] ),
    .X(_00177_));
 sky130_fd_sc_hd__a22o_1 _07216_ (.A1(net1077),
    .A2(net325),
    .B1(net227),
    .B2(\tms1x00.ins_pla_ors[13][21] ),
    .X(_00178_));
 sky130_fd_sc_hd__a22o_1 _07217_ (.A1(net105),
    .A2(net325),
    .B1(net227),
    .B2(\tms1x00.ins_pla_ors[13][25] ),
    .X(_00179_));
 sky130_fd_sc_hd__a22o_1 _07218_ (.A1(net1072),
    .A2(net325),
    .B1(net227),
    .B2(\tms1x00.ins_pla_ors[13][26] ),
    .X(_00180_));
 sky130_fd_sc_hd__a22o_1 _07219_ (.A1(net107),
    .A2(net325),
    .B1(net227),
    .B2(\tms1x00.ins_pla_ors[13][27] ),
    .X(_00181_));
 sky130_fd_sc_hd__a22o_1 _07220_ (.A1(net108),
    .A2(net326),
    .B1(net227),
    .B2(\tms1x00.ins_pla_ors[13][28] ),
    .X(_00182_));
 sky130_fd_sc_hd__a22o_1 _07221_ (.A1(net109),
    .A2(net326),
    .B1(_03528_),
    .B2(\tms1x00.ins_pla_ors[13][29] ),
    .X(_00183_));
 sky130_fd_sc_hd__nor2_4 _07222_ (.A(net852),
    .B(net355),
    .Y(_03531_));
 sky130_fd_sc_hd__nor2_2 _07223_ (.A(net522),
    .B(net323),
    .Y(_03532_));
 sky130_fd_sc_hd__mux2_1 _07224_ (.A0(_03476_),
    .A1(\tms1x00.ins_pla_ors[11][0] ),
    .S(net224),
    .X(_00184_));
 sky130_fd_sc_hd__or2_4 _07225_ (.A(_03424_),
    .B(net378),
    .X(_03533_));
 sky130_fd_sc_hd__mux2_1 _07226_ (.A0(net344),
    .A1(\tms1x00.ins_pla_ors[11][1] ),
    .S(net222),
    .X(_00185_));
 sky130_fd_sc_hd__or2_4 _07227_ (.A(net390),
    .B(_03430_),
    .X(_03534_));
 sky130_fd_sc_hd__mux2_1 _07228_ (.A0(_03534_),
    .A1(\tms1x00.ins_pla_ors[11][3] ),
    .S(net223),
    .X(_00186_));
 sky130_fd_sc_hd__or2_4 _07229_ (.A(net390),
    .B(_03478_),
    .X(_03535_));
 sky130_fd_sc_hd__mux2_1 _07230_ (.A0(_03535_),
    .A1(\tms1x00.ins_pla_ors[11][4] ),
    .S(net224),
    .X(_00187_));
 sky130_fd_sc_hd__mux2_1 _07231_ (.A0(_03480_),
    .A1(\tms1x00.ins_pla_ors[11][6] ),
    .S(net224),
    .X(_00188_));
 sky130_fd_sc_hd__or2_4 _07232_ (.A(net376),
    .B(net368),
    .X(_03536_));
 sky130_fd_sc_hd__mux2_1 _07233_ (.A0(_03536_),
    .A1(\tms1x00.ins_pla_ors[11][7] ),
    .S(net224),
    .X(_00189_));
 sky130_fd_sc_hd__mux2_1 _07234_ (.A0(_03487_),
    .A1(\tms1x00.ins_pla_ors[11][13] ),
    .S(net222),
    .X(_00190_));
 sky130_fd_sc_hd__a21o_2 _07235_ (.A1(net953),
    .A2(net461),
    .B1(net389),
    .X(_03537_));
 sky130_fd_sc_hd__mux2_1 _07236_ (.A0(_03537_),
    .A1(\tms1x00.ins_pla_ors[11][14] ),
    .S(net222),
    .X(_00191_));
 sky130_fd_sc_hd__a21o_1 _07237_ (.A1(net945),
    .A2(net323),
    .B1(net521),
    .X(_03538_));
 sky130_fd_sc_hd__a22o_1 _07238_ (.A1(\tms1x00.ins_pla_ors[11][15] ),
    .A2(net222),
    .B1(_03538_),
    .B2(_03432_),
    .X(_00192_));
 sky130_fd_sc_hd__a21o_1 _07239_ (.A1(net942),
    .A2(net324),
    .B1(net541),
    .X(_03539_));
 sky130_fd_sc_hd__a22o_1 _07240_ (.A1(\tms1x00.ins_pla_ors[11][16] ),
    .A2(net224),
    .B1(_03539_),
    .B2(net373),
    .X(_00193_));
 sky130_fd_sc_hd__or2_1 _07241_ (.A(net393),
    .B(_03442_),
    .X(_03540_));
 sky130_fd_sc_hd__mux2_1 _07242_ (.A0(_03540_),
    .A1(\tms1x00.ins_pla_ors[11][17] ),
    .S(net223),
    .X(_00194_));
 sky130_fd_sc_hd__and2_1 _07243_ (.A(net373),
    .B(_03444_),
    .X(_03541_));
 sky130_fd_sc_hd__mux2_1 _07244_ (.A0(_03541_),
    .A1(\tms1x00.ins_pla_ors[11][18] ),
    .S(net223),
    .X(_00195_));
 sky130_fd_sc_hd__or2_1 _07245_ (.A(net375),
    .B(_03464_),
    .X(_03542_));
 sky130_fd_sc_hd__mux2_1 _07246_ (.A0(_03542_),
    .A1(\tms1x00.ins_pla_ors[11][19] ),
    .S(net222),
    .X(_00196_));
 sky130_fd_sc_hd__a221o_1 _07247_ (.A1(_03446_),
    .A2(net323),
    .B1(net222),
    .B2(\tms1x00.ins_pla_ors[11][21] ),
    .C1(net375),
    .X(_00197_));
 sky130_fd_sc_hd__a21o_1 _07248_ (.A1(net1075),
    .A2(net479),
    .B1(net374),
    .X(_03543_));
 sky130_fd_sc_hd__mux2_1 _07249_ (.A0(_03543_),
    .A1(\tms1x00.ins_pla_ors[11][22] ),
    .S(net223),
    .X(_00198_));
 sky130_fd_sc_hd__a221o_1 _07250_ (.A1(_03498_),
    .A2(net324),
    .B1(net223),
    .B2(\tms1x00.ins_pla_ors[11][25] ),
    .C1(net381),
    .X(_00199_));
 sky130_fd_sc_hd__a21o_1 _07251_ (.A1(net1072),
    .A2(net324),
    .B1(net537),
    .X(_03544_));
 sky130_fd_sc_hd__a22o_1 _07252_ (.A1(\tms1x00.ins_pla_ors[11][26] ),
    .A2(net223),
    .B1(_03544_),
    .B2(net373),
    .X(_00200_));
 sky130_fd_sc_hd__nor2_8 _07253_ (.A(net864),
    .B(net346),
    .Y(_03545_));
 sky130_fd_sc_hd__or2_4 _07254_ (.A(net864),
    .B(net346),
    .X(_03546_));
 sky130_fd_sc_hd__mux2_1 _07255_ (.A0(net982),
    .A1(\tms1x00.ins_pla_ors[3][0] ),
    .S(net321),
    .X(_03547_));
 sky130_fd_sc_hd__or2_1 _07256_ (.A(net553),
    .B(_03547_),
    .X(_00201_));
 sky130_fd_sc_hd__mux2_1 _07257_ (.A0(net934),
    .A1(\tms1x00.ins_pla_ors[3][1] ),
    .S(net320),
    .X(_03548_));
 sky130_fd_sc_hd__or2_1 _07258_ (.A(net549),
    .B(_03548_),
    .X(_00202_));
 sky130_fd_sc_hd__mux2_1 _07259_ (.A0(net1053),
    .A1(\tms1x00.ins_pla_ors[3][4] ),
    .S(_03546_),
    .X(_03549_));
 sky130_fd_sc_hd__or2_1 _07260_ (.A(net554),
    .B(_03549_),
    .X(_00203_));
 sky130_fd_sc_hd__mux2_1 _07261_ (.A0(net1044),
    .A1(\tms1x00.ins_pla_ors[3][5] ),
    .S(net321),
    .X(_03550_));
 sky130_fd_sc_hd__or2_1 _07262_ (.A(net551),
    .B(_03550_),
    .X(_00204_));
 sky130_fd_sc_hd__mux2_1 _07263_ (.A0(net1037),
    .A1(\tms1x00.ins_pla_ors[3][6] ),
    .S(net322),
    .X(_03551_));
 sky130_fd_sc_hd__or2_1 _07264_ (.A(net550),
    .B(_03551_),
    .X(_00205_));
 sky130_fd_sc_hd__mux2_1 _07265_ (.A0(net1022),
    .A1(\tms1x00.ins_pla_ors[3][8] ),
    .S(net320),
    .X(_03552_));
 sky130_fd_sc_hd__or2_1 _07266_ (.A(net542),
    .B(_03552_),
    .X(_00206_));
 sky130_fd_sc_hd__mux2_1 _07267_ (.A0(net1013),
    .A1(\tms1x00.ins_pla_ors[3][9] ),
    .S(net322),
    .X(_03553_));
 sky130_fd_sc_hd__or2_1 _07268_ (.A(net552),
    .B(_03553_),
    .X(_00207_));
 sky130_fd_sc_hd__mux2_1 _07269_ (.A0(net975),
    .A1(\tms1x00.ins_pla_ors[3][10] ),
    .S(net322),
    .X(_03554_));
 sky130_fd_sc_hd__or2_1 _07270_ (.A(net552),
    .B(_03554_),
    .X(_00208_));
 sky130_fd_sc_hd__mux2_1 _07271_ (.A0(net970),
    .A1(\tms1x00.ins_pla_ors[3][11] ),
    .S(net320),
    .X(_03555_));
 sky130_fd_sc_hd__or2_1 _07272_ (.A(net541),
    .B(_03555_),
    .X(_00209_));
 sky130_fd_sc_hd__or2_1 _07273_ (.A(\tms1x00.ins_pla_ors[3][13] ),
    .B(_03545_),
    .X(_03556_));
 sky130_fd_sc_hd__o211a_1 _07274_ (.A1(net961),
    .A2(net322),
    .B1(_03556_),
    .C1(net486),
    .X(_00210_));
 sky130_fd_sc_hd__mux2_1 _07275_ (.A0(net948),
    .A1(\tms1x00.ins_pla_ors[3][15] ),
    .S(net320),
    .X(_03557_));
 sky130_fd_sc_hd__or2_1 _07276_ (.A(net544),
    .B(_03557_),
    .X(_00211_));
 sky130_fd_sc_hd__mux2_1 _07277_ (.A0(net943),
    .A1(\tms1x00.ins_pla_ors[3][16] ),
    .S(net322),
    .X(_03558_));
 sky130_fd_sc_hd__or2_1 _07278_ (.A(net552),
    .B(_03558_),
    .X(_00212_));
 sky130_fd_sc_hd__mux2_1 _07279_ (.A0(net940),
    .A1(\tms1x00.ins_pla_ors[3][17] ),
    .S(net321),
    .X(_03559_));
 sky130_fd_sc_hd__or2_1 _07280_ (.A(net550),
    .B(_03559_),
    .X(_00213_));
 sky130_fd_sc_hd__mux2_1 _07281_ (.A0(net938),
    .A1(\tms1x00.ins_pla_ors[3][18] ),
    .S(net321),
    .X(_03560_));
 sky130_fd_sc_hd__or2_1 _07282_ (.A(net547),
    .B(_03560_),
    .X(_00214_));
 sky130_fd_sc_hd__mux2_1 _07283_ (.A0(net935),
    .A1(\tms1x00.ins_pla_ors[3][19] ),
    .S(net321),
    .X(_03561_));
 sky130_fd_sc_hd__or2_1 _07284_ (.A(net550),
    .B(_03561_),
    .X(_00215_));
 sky130_fd_sc_hd__mux2_1 _07285_ (.A0(net1078),
    .A1(\tms1x00.ins_pla_ors[3][20] ),
    .S(net321),
    .X(_03562_));
 sky130_fd_sc_hd__or2_1 _07286_ (.A(net546),
    .B(_03562_),
    .X(_00216_));
 sky130_fd_sc_hd__or2_1 _07287_ (.A(\tms1x00.ins_pla_ors[3][22] ),
    .B(_03545_),
    .X(_03563_));
 sky130_fd_sc_hd__o211a_1 _07288_ (.A1(net1075),
    .A2(net320),
    .B1(_03563_),
    .C1(net482),
    .X(_00217_));
 sky130_fd_sc_hd__mux2_1 _07289_ (.A0(net1074),
    .A1(\tms1x00.ins_pla_ors[3][23] ),
    .S(net321),
    .X(_03564_));
 sky130_fd_sc_hd__or2_1 _07290_ (.A(net551),
    .B(_03564_),
    .X(_00218_));
 sky130_fd_sc_hd__mux2_1 _07291_ (.A0(net1072),
    .A1(\tms1x00.ins_pla_ors[3][26] ),
    .S(net321),
    .X(_03565_));
 sky130_fd_sc_hd__or2_1 _07292_ (.A(net548),
    .B(_03565_),
    .X(_00219_));
 sky130_fd_sc_hd__or2_1 _07293_ (.A(\tms1x00.ins_pla_ors[3][27] ),
    .B(_03545_),
    .X(_03566_));
 sky130_fd_sc_hd__o211a_1 _07294_ (.A1(net107),
    .A2(net320),
    .B1(_03566_),
    .C1(net489),
    .X(_00220_));
 sky130_fd_sc_hd__or2_1 _07295_ (.A(\tms1x00.ins_pla_ors[3][28] ),
    .B(_03545_),
    .X(_03567_));
 sky130_fd_sc_hd__o211a_1 _07296_ (.A1(net108),
    .A2(net320),
    .B1(_03567_),
    .C1(net482),
    .X(_00221_));
 sky130_fd_sc_hd__nor2_2 _07297_ (.A(net988),
    .B(net995),
    .Y(_03568_));
 sky130_fd_sc_hd__or2_1 _07298_ (.A(net987),
    .B(net995),
    .X(_03569_));
 sky130_fd_sc_hd__and3_4 _07299_ (.A(net628),
    .B(net352),
    .C(net708),
    .X(_03570_));
 sky130_fd_sc_hd__or3_4 _07300_ (.A(net615),
    .B(net349),
    .C(net707),
    .X(_03571_));
 sky130_fd_sc_hd__nor2_2 _07301_ (.A(net378),
    .B(_03570_),
    .Y(_03572_));
 sky130_fd_sc_hd__nand2_2 _07302_ (.A(net370),
    .B(_03571_),
    .Y(_03573_));
 sky130_fd_sc_hd__or2_4 _07303_ (.A(net982),
    .B(net382),
    .X(_03574_));
 sky130_fd_sc_hd__o221a_1 _07304_ (.A1(\tms1x00.ins_pla_ands[6][0] ),
    .A2(_03573_),
    .B1(_03574_),
    .B2(_03571_),
    .C1(net384),
    .X(_00222_));
 sky130_fd_sc_hd__nor2_2 _07305_ (.A(net392),
    .B(_03570_),
    .Y(_03575_));
 sky130_fd_sc_hd__nand2_2 _07306_ (.A(net384),
    .B(_03571_),
    .Y(_03576_));
 sky130_fd_sc_hd__a22o_1 _07307_ (.A1(\tms1x00.ins_pla_ands[6][1] ),
    .A2(_03572_),
    .B1(_03576_),
    .B2(net354),
    .X(_00223_));
 sky130_fd_sc_hd__a22o_1 _07308_ (.A1(\tms1x00.ins_pla_ands[6][4] ),
    .A2(_03572_),
    .B1(_03576_),
    .B2(_03535_),
    .X(_00224_));
 sky130_fd_sc_hd__or2_4 _07309_ (.A(net375),
    .B(net366),
    .X(_03577_));
 sky130_fd_sc_hd__o22a_1 _07310_ (.A1(\tms1x00.ins_pla_ands[6][5] ),
    .A2(_03573_),
    .B1(_03575_),
    .B2(_03577_),
    .X(_00225_));
 sky130_fd_sc_hd__a22o_1 _07311_ (.A1(\tms1x00.ins_pla_ands[6][6] ),
    .A2(_03572_),
    .B1(_03576_),
    .B2(_03435_),
    .X(_00226_));
 sky130_fd_sc_hd__o22a_1 _07312_ (.A1(\tms1x00.ins_pla_ands[6][7] ),
    .A2(_03573_),
    .B1(_03575_),
    .B2(_03536_),
    .X(_00227_));
 sky130_fd_sc_hd__a22o_1 _07313_ (.A1(\tms1x00.ins_pla_ands[6][8] ),
    .A2(_03572_),
    .B1(_03576_),
    .B2(net353),
    .X(_00228_));
 sky130_fd_sc_hd__or2_4 _07314_ (.A(net377),
    .B(net365),
    .X(_03578_));
 sky130_fd_sc_hd__o22a_1 _07315_ (.A1(\tms1x00.ins_pla_ands[6][9] ),
    .A2(_03573_),
    .B1(_03575_),
    .B2(_03578_),
    .X(_00229_));
 sky130_fd_sc_hd__or2_4 _07316_ (.A(net390),
    .B(_03459_),
    .X(_03579_));
 sky130_fd_sc_hd__a22o_1 _07317_ (.A1(\tms1x00.ins_pla_ands[6][10] ),
    .A2(_03572_),
    .B1(_03576_),
    .B2(_03579_),
    .X(_00230_));
 sky130_fd_sc_hd__or2_4 _07318_ (.A(net374),
    .B(_03460_),
    .X(_03580_));
 sky130_fd_sc_hd__o22a_1 _07319_ (.A1(\tms1x00.ins_pla_ands[6][11] ),
    .A2(_03573_),
    .B1(_03575_),
    .B2(_03580_),
    .X(_00231_));
 sky130_fd_sc_hd__and3_4 _07320_ (.A(net739),
    .B(net352),
    .C(net708),
    .X(_03581_));
 sky130_fd_sc_hd__or3_4 _07321_ (.A(net733),
    .B(net349),
    .C(net706),
    .X(_03582_));
 sky130_fd_sc_hd__nor2_4 _07322_ (.A(net377),
    .B(_03581_),
    .Y(_03583_));
 sky130_fd_sc_hd__nand2_1 _07323_ (.A(net373),
    .B(_03582_),
    .Y(_03584_));
 sky130_fd_sc_hd__or2_4 _07324_ (.A(net389),
    .B(_03456_),
    .X(_03585_));
 sky130_fd_sc_hd__nor2_1 _07325_ (.A(net396),
    .B(_03581_),
    .Y(_03586_));
 sky130_fd_sc_hd__nand2_4 _07326_ (.A(net384),
    .B(_03582_),
    .Y(_03587_));
 sky130_fd_sc_hd__a22o_1 _07327_ (.A1(\tms1x00.ins_pla_ands[2][0] ),
    .A2(_03583_),
    .B1(_03585_),
    .B2(_03587_),
    .X(_00232_));
 sky130_fd_sc_hd__a22o_1 _07328_ (.A1(\tms1x00.ins_pla_ands[2][2] ),
    .A2(_03583_),
    .B1(_03587_),
    .B2(_03429_),
    .X(_00233_));
 sky130_fd_sc_hd__a22o_1 _07329_ (.A1(\tms1x00.ins_pla_ands[2][4] ),
    .A2(_03583_),
    .B1(_03587_),
    .B2(_03535_),
    .X(_00234_));
 sky130_fd_sc_hd__a22o_1 _07330_ (.A1(\tms1x00.ins_pla_ands[2][7] ),
    .A2(_03583_),
    .B1(_03587_),
    .B2(_03437_),
    .X(_00235_));
 sky130_fd_sc_hd__a22o_1 _07331_ (.A1(\tms1x00.ins_pla_ands[2][10] ),
    .A2(_03583_),
    .B1(_03587_),
    .B2(_03579_),
    .X(_00236_));
 sky130_fd_sc_hd__o22a_1 _07332_ (.A1(\tms1x00.ins_pla_ands[2][11] ),
    .A2(_03584_),
    .B1(_03586_),
    .B2(_03580_),
    .X(_00237_));
 sky130_fd_sc_hd__or2_4 _07333_ (.A(net389),
    .B(_03484_),
    .X(_03588_));
 sky130_fd_sc_hd__a22o_1 _07334_ (.A1(\tms1x00.ins_pla_ands[2][12] ),
    .A2(_03583_),
    .B1(_03587_),
    .B2(_03588_),
    .X(_00238_));
 sky130_fd_sc_hd__or2_4 _07335_ (.A(net378),
    .B(_03486_),
    .X(_03589_));
 sky130_fd_sc_hd__o22a_1 _07336_ (.A1(\tms1x00.ins_pla_ands[2][13] ),
    .A2(_03584_),
    .B1(_03586_),
    .B2(_03589_),
    .X(_00239_));
 sky130_fd_sc_hd__and3_4 _07337_ (.A(net902),
    .B(net350),
    .C(_03471_),
    .X(_03590_));
 sky130_fd_sc_hd__nor2_1 _07338_ (.A(net512),
    .B(net319),
    .Y(_03591_));
 sky130_fd_sc_hd__o22a_1 _07339_ (.A1(\tms1x00.ins_pla_ands[29][0] ),
    .A2(net319),
    .B1(net220),
    .B2(_03456_),
    .X(_00240_));
 sky130_fd_sc_hd__o22a_1 _07340_ (.A1(\tms1x00.ins_pla_ands[29][1] ),
    .A2(net319),
    .B1(net221),
    .B2(net397),
    .X(_00241_));
 sky130_fd_sc_hd__o22a_1 _07341_ (.A1(\tms1x00.ins_pla_ands[29][2] ),
    .A2(net319),
    .B1(net220),
    .B2(_03428_),
    .X(_00242_));
 sky130_fd_sc_hd__o22a_1 _07342_ (.A1(\tms1x00.ins_pla_ands[29][3] ),
    .A2(net319),
    .B1(net221),
    .B2(_03430_),
    .X(_00243_));
 sky130_fd_sc_hd__o22a_1 _07343_ (.A1(\tms1x00.ins_pla_ands[29][4] ),
    .A2(_03590_),
    .B1(net220),
    .B2(_03478_),
    .X(_00244_));
 sky130_fd_sc_hd__o22a_1 _07344_ (.A1(\tms1x00.ins_pla_ands[29][5] ),
    .A2(_03590_),
    .B1(net221),
    .B2(net366),
    .X(_00245_));
 sky130_fd_sc_hd__o22a_1 _07345_ (.A1(\tms1x00.ins_pla_ands[29][6] ),
    .A2(net319),
    .B1(net221),
    .B2(_03434_),
    .X(_00246_));
 sky130_fd_sc_hd__o22a_1 _07346_ (.A1(\tms1x00.ins_pla_ands[29][7] ),
    .A2(net319),
    .B1(net221),
    .B2(net367),
    .X(_00247_));
 sky130_fd_sc_hd__o22a_1 _07347_ (.A1(\tms1x00.ins_pla_ands[29][9] ),
    .A2(net319),
    .B1(net220),
    .B2(net365),
    .X(_00248_));
 sky130_fd_sc_hd__o22a_1 _07348_ (.A1(\tms1x00.ins_pla_ands[29][11] ),
    .A2(_03590_),
    .B1(net220),
    .B2(_03460_),
    .X(_00249_));
 sky130_fd_sc_hd__o22a_1 _07349_ (.A1(\tms1x00.ins_pla_ands[29][12] ),
    .A2(net319),
    .B1(net220),
    .B2(_03484_),
    .X(_00250_));
 sky130_fd_sc_hd__mux2_1 _07350_ (.A0(\tms1x00.ins_pla_ands[29][15] ),
    .A1(net945),
    .S(net319),
    .X(_03592_));
 sky130_fd_sc_hd__and2_1 _07351_ (.A(net460),
    .B(_03592_),
    .X(_00251_));
 sky130_fd_sc_hd__and3_4 _07352_ (.A(net874),
    .B(net350),
    .C(_03471_),
    .X(_03593_));
 sky130_fd_sc_hd__nor2_1 _07353_ (.A(net522),
    .B(_03593_),
    .Y(_03594_));
 sky130_fd_sc_hd__mux2_1 _07354_ (.A0(net353),
    .A1(\tms1x00.ins_pla_ands[27][8] ),
    .S(net218),
    .X(_00252_));
 sky130_fd_sc_hd__mux2_1 _07355_ (.A0(_03483_),
    .A1(\tms1x00.ins_pla_ands[27][11] ),
    .S(net218),
    .X(_00253_));
 sky130_fd_sc_hd__mux2_1 _07356_ (.A0(_03487_),
    .A1(\tms1x00.ins_pla_ands[27][13] ),
    .S(net219),
    .X(_00254_));
 sky130_fd_sc_hd__mux2_1 _07357_ (.A0(_03537_),
    .A1(\tms1x00.ins_pla_ands[27][14] ),
    .S(net219),
    .X(_00255_));
 sky130_fd_sc_hd__and3_4 _07358_ (.A(net795),
    .B(net598),
    .C(net350),
    .X(_03595_));
 sky130_fd_sc_hd__nor2_8 _07359_ (.A(net514),
    .B(net317),
    .Y(_03596_));
 sky130_fd_sc_hd__mux2_1 _07360_ (.A0(net343),
    .A1(\tms1x00.ins_pla_ands[23][0] ),
    .S(_03596_),
    .X(_00256_));
 sky130_fd_sc_hd__mux2_1 _07361_ (.A0(net344),
    .A1(\tms1x00.ins_pla_ands[23][1] ),
    .S(_03596_),
    .X(_00257_));
 sky130_fd_sc_hd__mux2_1 _07362_ (.A0(_03482_),
    .A1(\tms1x00.ins_pla_ands[23][10] ),
    .S(_03596_),
    .X(_00258_));
 sky130_fd_sc_hd__mux2_1 _07363_ (.A0(net347),
    .A1(\tms1x00.ins_pla_ands[23][11] ),
    .S(_03596_),
    .X(_00259_));
 sky130_fd_sc_hd__and3_1 _07364_ (.A(net628),
    .B(net598),
    .C(net350),
    .X(_03597_));
 sky130_fd_sc_hd__nor2_2 _07365_ (.A(net516),
    .B(net316),
    .Y(_03598_));
 sky130_fd_sc_hd__or2_4 _07366_ (.A(net524),
    .B(net316),
    .X(_03599_));
 sky130_fd_sc_hd__mux2_1 _07367_ (.A0(\tms1x00.ins_pla_ands[22][0] ),
    .A1(_03476_),
    .S(_03599_),
    .X(_00260_));
 sky130_fd_sc_hd__mux2_1 _07368_ (.A0(\tms1x00.ins_pla_ands[22][1] ),
    .A1(net354),
    .S(_03599_),
    .X(_00261_));
 sky130_fd_sc_hd__mux2_1 _07369_ (.A0(\tms1x00.ins_pla_ands[22][2] ),
    .A1(_03477_),
    .S(_03599_),
    .X(_00262_));
 sky130_fd_sc_hd__mux2_1 _07370_ (.A0(\tms1x00.ins_pla_ands[22][3] ),
    .A1(_03534_),
    .S(_03599_),
    .X(_00263_));
 sky130_fd_sc_hd__mux2_1 _07371_ (.A0(\tms1x00.ins_pla_ands[22][4] ),
    .A1(_03535_),
    .S(_03599_),
    .X(_00264_));
 sky130_fd_sc_hd__mux2_1 _07372_ (.A0(\tms1x00.ins_pla_ands[22][5] ),
    .A1(_03577_),
    .S(_03599_),
    .X(_00265_));
 sky130_fd_sc_hd__mux2_1 _07373_ (.A0(\tms1x00.ins_pla_ands[22][11] ),
    .A1(net347),
    .S(_03599_),
    .X(_00266_));
 sky130_fd_sc_hd__and3_4 _07374_ (.A(net874),
    .B(net598),
    .C(_03469_),
    .X(_03600_));
 sky130_fd_sc_hd__nor2_8 _07375_ (.A(net517),
    .B(net315),
    .Y(_03601_));
 sky130_fd_sc_hd__o22a_1 _07376_ (.A1(\tms1x00.ins_pla_ands[19][2] ),
    .A2(_03600_),
    .B1(_03601_),
    .B2(_03428_),
    .X(_00267_));
 sky130_fd_sc_hd__mux2_1 _07377_ (.A0(\tms1x00.ins_pla_ands[19][3] ),
    .A1(net1058),
    .S(net315),
    .X(_03602_));
 sky130_fd_sc_hd__or2_1 _07378_ (.A(net516),
    .B(_03602_),
    .X(_00268_));
 sky130_fd_sc_hd__o22a_1 _07379_ (.A1(\tms1x00.ins_pla_ands[19][4] ),
    .A2(net315),
    .B1(_03601_),
    .B2(_03478_),
    .X(_00269_));
 sky130_fd_sc_hd__mux2_1 _07380_ (.A0(\tms1x00.ins_pla_ands[19][5] ),
    .A1(net1041),
    .S(_03600_),
    .X(_03603_));
 sky130_fd_sc_hd__or2_1 _07381_ (.A(net524),
    .B(_03603_),
    .X(_00270_));
 sky130_fd_sc_hd__mux2_1 _07382_ (.A0(\tms1x00.ins_pla_ands[19][6] ),
    .A1(net1033),
    .S(net315),
    .X(_03604_));
 sky130_fd_sc_hd__or2_1 _07383_ (.A(net524),
    .B(_03604_),
    .X(_00271_));
 sky130_fd_sc_hd__o22a_1 _07384_ (.A1(\tms1x00.ins_pla_ands[19][7] ),
    .A2(_03600_),
    .B1(_03601_),
    .B2(net368),
    .X(_00272_));
 sky130_fd_sc_hd__mux2_1 _07385_ (.A0(\tms1x00.ins_pla_ands[19][8] ),
    .A1(net1014),
    .S(net315),
    .X(_03605_));
 sky130_fd_sc_hd__or2_1 _07386_ (.A(net515),
    .B(_03605_),
    .X(_00273_));
 sky130_fd_sc_hd__o22a_1 _07387_ (.A1(\tms1x00.ins_pla_ands[19][9] ),
    .A2(net315),
    .B1(_03601_),
    .B2(net364),
    .X(_00274_));
 sky130_fd_sc_hd__mux2_1 _07388_ (.A0(\tms1x00.ins_pla_ands[19][12] ),
    .A1(net963),
    .S(net315),
    .X(_03606_));
 sky130_fd_sc_hd__or2_1 _07389_ (.A(net515),
    .B(_03606_),
    .X(_00275_));
 sky130_fd_sc_hd__o22a_1 _07390_ (.A1(\tms1x00.ins_pla_ands[19][13] ),
    .A2(net315),
    .B1(_03601_),
    .B2(net363),
    .X(_00276_));
 sky130_fd_sc_hd__mux2_1 _07391_ (.A0(\tms1x00.ins_pla_ands[19][14] ),
    .A1(net951),
    .S(net315),
    .X(_03607_));
 sky130_fd_sc_hd__or2_1 _07392_ (.A(net513),
    .B(_03607_),
    .X(_00277_));
 sky130_fd_sc_hd__mux2_1 _07393_ (.A0(\tms1x00.ins_pla_ands[19][15] ),
    .A1(net944),
    .S(net315),
    .X(_03608_));
 sky130_fd_sc_hd__and2_1 _07394_ (.A(net459),
    .B(_03608_),
    .X(_00278_));
 sky130_fd_sc_hd__mux2_1 _07395_ (.A0(net979),
    .A1(\tms1x00.ins_pla_ors[8][0] ),
    .S(net327),
    .X(_03609_));
 sky130_fd_sc_hd__or2_1 _07396_ (.A(net519),
    .B(_03609_),
    .X(_00279_));
 sky130_fd_sc_hd__mux2_1 _07397_ (.A0(net930),
    .A1(\tms1x00.ins_pla_ors[8][1] ),
    .S(net327),
    .X(_03610_));
 sky130_fd_sc_hd__or2_1 _07398_ (.A(net523),
    .B(_03610_),
    .X(_00280_));
 sky130_fd_sc_hd__mux2_1 _07399_ (.A0(net1070),
    .A1(\tms1x00.ins_pla_ors[8][2] ),
    .S(net328),
    .X(_03611_));
 sky130_fd_sc_hd__or2_1 _07400_ (.A(net540),
    .B(_03611_),
    .X(_00281_));
 sky130_fd_sc_hd__mux2_1 _07401_ (.A0(net1058),
    .A1(\tms1x00.ins_pla_ors[8][3] ),
    .S(net327),
    .X(_03612_));
 sky130_fd_sc_hd__or2_1 _07402_ (.A(net520),
    .B(_03612_),
    .X(_00282_));
 sky130_fd_sc_hd__mux2_1 _07403_ (.A0(net1053),
    .A1(\tms1x00.ins_pla_ors[8][4] ),
    .S(net329),
    .X(_03613_));
 sky130_fd_sc_hd__or2_1 _07404_ (.A(net543),
    .B(_03613_),
    .X(_00283_));
 sky130_fd_sc_hd__mux2_1 _07405_ (.A0(net1041),
    .A1(\tms1x00.ins_pla_ors[8][5] ),
    .S(net327),
    .X(_03614_));
 sky130_fd_sc_hd__or2_1 _07406_ (.A(net523),
    .B(_03614_),
    .X(_00284_));
 sky130_fd_sc_hd__mux2_1 _07407_ (.A0(net1037),
    .A1(\tms1x00.ins_pla_ors[8][6] ),
    .S(net328),
    .X(_03615_));
 sky130_fd_sc_hd__or2_1 _07408_ (.A(net537),
    .B(_03615_),
    .X(_00285_));
 sky130_fd_sc_hd__mux2_1 _07409_ (.A0(net1026),
    .A1(\tms1x00.ins_pla_ors[8][7] ),
    .S(net329),
    .X(_03616_));
 sky130_fd_sc_hd__or2_1 _07410_ (.A(net523),
    .B(_03616_),
    .X(_00286_));
 sky130_fd_sc_hd__mux2_1 _07411_ (.A0(net1022),
    .A1(\tms1x00.ins_pla_ors[8][8] ),
    .S(net329),
    .X(_03617_));
 sky130_fd_sc_hd__or2_1 _07412_ (.A(net540),
    .B(_03617_),
    .X(_00287_));
 sky130_fd_sc_hd__mux2_1 _07413_ (.A0(net1010),
    .A1(\tms1x00.ins_pla_ors[8][9] ),
    .S(net327),
    .X(_03618_));
 sky130_fd_sc_hd__or2_1 _07414_ (.A(net521),
    .B(_03618_),
    .X(_00288_));
 sky130_fd_sc_hd__mux2_1 _07415_ (.A0(net972),
    .A1(\tms1x00.ins_pla_ors[8][10] ),
    .S(net327),
    .X(_03619_));
 sky130_fd_sc_hd__or2_1 _07416_ (.A(net521),
    .B(_03619_),
    .X(_00289_));
 sky130_fd_sc_hd__mux2_1 _07417_ (.A0(net968),
    .A1(\tms1x00.ins_pla_ors[8][11] ),
    .S(net327),
    .X(_03620_));
 sky130_fd_sc_hd__or2_1 _07418_ (.A(net523),
    .B(_03620_),
    .X(_00290_));
 sky130_fd_sc_hd__mux2_1 _07419_ (.A0(net953),
    .A1(\tms1x00.ins_pla_ors[8][14] ),
    .S(net327),
    .X(_03621_));
 sky130_fd_sc_hd__or2_1 _07420_ (.A(net521),
    .B(_03621_),
    .X(_00291_));
 sky130_fd_sc_hd__mux2_1 _07421_ (.A0(net942),
    .A1(\tms1x00.ins_pla_ors[8][16] ),
    .S(net328),
    .X(_03622_));
 sky130_fd_sc_hd__or2_1 _07422_ (.A(net538),
    .B(_03622_),
    .X(_00292_));
 sky130_fd_sc_hd__mux2_1 _07423_ (.A0(net940),
    .A1(\tms1x00.ins_pla_ors[8][17] ),
    .S(net328),
    .X(_03623_));
 sky130_fd_sc_hd__or2_1 _07424_ (.A(net538),
    .B(_03623_),
    .X(_00293_));
 sky130_fd_sc_hd__mux2_1 _07425_ (.A0(net938),
    .A1(\tms1x00.ins_pla_ors[8][18] ),
    .S(net329),
    .X(_03624_));
 sky130_fd_sc_hd__or2_1 _07426_ (.A(net540),
    .B(_03624_),
    .X(_00294_));
 sky130_fd_sc_hd__mux2_1 _07427_ (.A0(net1078),
    .A1(\tms1x00.ins_pla_ors[8][20] ),
    .S(net328),
    .X(_03625_));
 sky130_fd_sc_hd__or2_1 _07428_ (.A(net538),
    .B(_03625_),
    .X(_00295_));
 sky130_fd_sc_hd__mux2_1 _07429_ (.A0(net1077),
    .A1(\tms1x00.ins_pla_ors[8][21] ),
    .S(net327),
    .X(_03626_));
 sky130_fd_sc_hd__or2_1 _07430_ (.A(net520),
    .B(_03626_),
    .X(_00296_));
 sky130_fd_sc_hd__mux2_1 _07431_ (.A0(net1074),
    .A1(\tms1x00.ins_pla_ors[8][23] ),
    .S(net328),
    .X(_03627_));
 sky130_fd_sc_hd__or2_1 _07432_ (.A(net537),
    .B(_03627_),
    .X(_00297_));
 sky130_fd_sc_hd__mux2_1 _07433_ (.A0(net1073),
    .A1(\tms1x00.ins_pla_ors[8][24] ),
    .S(net328),
    .X(_03628_));
 sky130_fd_sc_hd__or2_1 _07434_ (.A(net537),
    .B(_03628_),
    .X(_00298_));
 sky130_fd_sc_hd__mux2_1 _07435_ (.A0(net105),
    .A1(\tms1x00.ins_pla_ors[8][25] ),
    .S(net328),
    .X(_03629_));
 sky130_fd_sc_hd__or2_1 _07436_ (.A(net537),
    .B(_03629_),
    .X(_00299_));
 sky130_fd_sc_hd__mux2_1 _07437_ (.A0(net1072),
    .A1(\tms1x00.ins_pla_ors[8][26] ),
    .S(net328),
    .X(_03630_));
 sky130_fd_sc_hd__or2_1 _07438_ (.A(net537),
    .B(_03630_),
    .X(_00300_));
 sky130_fd_sc_hd__nor2_8 _07439_ (.A(net729),
    .B(net346),
    .Y(_03631_));
 sky130_fd_sc_hd__or2_1 _07440_ (.A(net729),
    .B(net346),
    .X(_03632_));
 sky130_fd_sc_hd__nor2_4 _07441_ (.A(net379),
    .B(_03631_),
    .Y(_03633_));
 sky130_fd_sc_hd__nand2_2 _07442_ (.A(net372),
    .B(net312),
    .Y(_03634_));
 sky130_fd_sc_hd__nand2_1 _07443_ (.A(net386),
    .B(net314),
    .Y(_03635_));
 sky130_fd_sc_hd__a22o_1 _07444_ (.A1(\tms1x00.ins_pla_ors[2][0] ),
    .A2(_03633_),
    .B1(_03635_),
    .B2(net343),
    .X(_00301_));
 sky130_fd_sc_hd__o221a_1 _07445_ (.A1(net1070),
    .A2(net312),
    .B1(_03634_),
    .B2(\tms1x00.ins_pla_ors[2][2] ),
    .C1(net386),
    .X(_00302_));
 sky130_fd_sc_hd__o221a_1 _07446_ (.A1(net1062),
    .A2(net312),
    .B1(_03634_),
    .B2(\tms1x00.ins_pla_ors[2][3] ),
    .C1(net386),
    .X(_00303_));
 sky130_fd_sc_hd__o221a_1 _07447_ (.A1(net1022),
    .A2(net313),
    .B1(_03634_),
    .B2(\tms1x00.ins_pla_ors[2][8] ),
    .C1(net386),
    .X(_00304_));
 sky130_fd_sc_hd__a221o_1 _07448_ (.A1(net940),
    .A2(_03631_),
    .B1(_03633_),
    .B2(\tms1x00.ins_pla_ors[2][17] ),
    .C1(net395),
    .X(_00305_));
 sky130_fd_sc_hd__a221o_1 _07449_ (.A1(net938),
    .A2(_03631_),
    .B1(_03633_),
    .B2(\tms1x00.ins_pla_ors[2][18] ),
    .C1(net394),
    .X(_00306_));
 sky130_fd_sc_hd__o221a_1 _07450_ (.A1(net1072),
    .A2(net314),
    .B1(_03634_),
    .B2(\tms1x00.ins_pla_ors[2][26] ),
    .C1(net386),
    .X(_00307_));
 sky130_fd_sc_hd__or2_4 _07451_ (.A(net393),
    .B(_03500_),
    .X(_03636_));
 sky130_fd_sc_hd__a22o_1 _07452_ (.A1(\tms1x00.ins_pla_ors[2][27] ),
    .A2(_03633_),
    .B1(_03635_),
    .B2(_03636_),
    .X(_00308_));
 sky130_fd_sc_hd__a22o_1 _07453_ (.A1(\tms1x00.ins_pla_ors[2][28] ),
    .A2(_03633_),
    .B1(_03635_),
    .B2(_03450_),
    .X(_00309_));
 sky130_fd_sc_hd__nor2_4 _07454_ (.A(net759),
    .B(net345),
    .Y(_03637_));
 sky130_fd_sc_hd__or2_4 _07455_ (.A(net759),
    .B(net345),
    .X(_03638_));
 sky130_fd_sc_hd__o31a_1 _07456_ (.A1(net1070),
    .A2(net379),
    .A3(net308),
    .B1(net387),
    .X(_03639_));
 sky130_fd_sc_hd__o31a_1 _07457_ (.A1(\tms1x00.ins_pla_ors[1][2] ),
    .A2(net380),
    .A3(net311),
    .B1(_03639_),
    .X(_00310_));
 sky130_fd_sc_hd__a31o_1 _07458_ (.A1(\tms1x00.ins_pla_ors[1][27] ),
    .A2(net371),
    .A3(net308),
    .B1(net394),
    .X(_03640_));
 sky130_fd_sc_hd__a21o_1 _07459_ (.A1(_03500_),
    .A2(net311),
    .B1(_03640_),
    .X(_00311_));
 sky130_fd_sc_hd__o22a_1 _07460_ (.A1(\tms1x00.ins_pla_ors[12][0] ),
    .A2(_03420_),
    .B1(_03422_),
    .B2(_03456_),
    .X(_00312_));
 sky130_fd_sc_hd__mux2_1 _07461_ (.A0(net1053),
    .A1(\tms1x00.ins_pla_ors[12][4] ),
    .S(net338),
    .X(_03641_));
 sky130_fd_sc_hd__or2_1 _07462_ (.A(net540),
    .B(_03641_),
    .X(_00313_));
 sky130_fd_sc_hd__mux2_1 _07463_ (.A0(net1041),
    .A1(\tms1x00.ins_pla_ors[12][5] ),
    .S(net338),
    .X(_03642_));
 sky130_fd_sc_hd__or2_1 _07464_ (.A(net523),
    .B(_03642_),
    .X(_00314_));
 sky130_fd_sc_hd__mux2_1 _07465_ (.A0(net1010),
    .A1(\tms1x00.ins_pla_ors[12][9] ),
    .S(net338),
    .X(_03643_));
 sky130_fd_sc_hd__or2_1 _07466_ (.A(net523),
    .B(_03643_),
    .X(_00315_));
 sky130_fd_sc_hd__mux2_1 _07467_ (.A0(net972),
    .A1(\tms1x00.ins_pla_ors[12][10] ),
    .S(net338),
    .X(_03644_));
 sky130_fd_sc_hd__or2_1 _07468_ (.A(net523),
    .B(_03644_),
    .X(_00316_));
 sky130_fd_sc_hd__mux2_1 _07469_ (.A0(net971),
    .A1(\tms1x00.ins_pla_ors[12][11] ),
    .S(net338),
    .X(_03645_));
 sky130_fd_sc_hd__or2_1 _07470_ (.A(net523),
    .B(_03645_),
    .X(_00317_));
 sky130_fd_sc_hd__o22a_1 _07471_ (.A1(\tms1x00.ins_pla_ors[12][12] ),
    .A2(_03420_),
    .B1(_03422_),
    .B2(_03484_),
    .X(_00318_));
 sky130_fd_sc_hd__mux2_1 _07472_ (.A0(net92),
    .A1(\tms1x00.ins_pla_ors[12][13] ),
    .S(net338),
    .X(_03646_));
 sky130_fd_sc_hd__or2_1 _07473_ (.A(net523),
    .B(_03646_),
    .X(_00319_));
 sky130_fd_sc_hd__a22o_1 _07474_ (.A1(\tms1x00.ins_pla_ors[12][15] ),
    .A2(net338),
    .B1(net234),
    .B2(_03530_),
    .X(_00320_));
 sky130_fd_sc_hd__mux2_1 _07475_ (.A0(net937),
    .A1(\tms1x00.ins_pla_ors[12][19] ),
    .S(net338),
    .X(_03647_));
 sky130_fd_sc_hd__or2_1 _07476_ (.A(net523),
    .B(_03647_),
    .X(_00321_));
 sky130_fd_sc_hd__mux2_1 _07477_ (.A0(net1078),
    .A1(\tms1x00.ins_pla_ors[12][20] ),
    .S(net338),
    .X(_03648_));
 sky130_fd_sc_hd__or2_1 _07478_ (.A(net538),
    .B(_03648_),
    .X(_00322_));
 sky130_fd_sc_hd__mux2_1 _07479_ (.A0(net1075),
    .A1(\tms1x00.ins_pla_ors[12][22] ),
    .S(_03421_),
    .X(_03649_));
 sky130_fd_sc_hd__or2_1 _07480_ (.A(net538),
    .B(_03649_),
    .X(_00323_));
 sky130_fd_sc_hd__mux2_1 _07481_ (.A0(net1074),
    .A1(\tms1x00.ins_pla_ors[12][23] ),
    .S(_03421_),
    .X(_03650_));
 sky130_fd_sc_hd__or2_1 _07482_ (.A(net538),
    .B(_03650_),
    .X(_00324_));
 sky130_fd_sc_hd__mux2_1 _07483_ (.A0(net1073),
    .A1(\tms1x00.ins_pla_ors[12][24] ),
    .S(_03421_),
    .X(_03651_));
 sky130_fd_sc_hd__or2_1 _07484_ (.A(net540),
    .B(_03651_),
    .X(_00325_));
 sky130_fd_sc_hd__o22a_1 _07485_ (.A1(\tms1x00.ins_pla_ors[12][25] ),
    .A2(_03420_),
    .B1(_03422_),
    .B2(_03498_),
    .X(_00326_));
 sky130_fd_sc_hd__o22a_1 _07486_ (.A1(\tms1x00.ins_pla_ors[12][27] ),
    .A2(_03420_),
    .B1(_03422_),
    .B2(_03500_),
    .X(_00327_));
 sky130_fd_sc_hd__mux2_1 _07487_ (.A0(_03477_),
    .A1(\tms1x00.ins_pla_ors[14][2] ),
    .S(net231),
    .X(_00328_));
 sky130_fd_sc_hd__mux2_1 _07488_ (.A0(_03479_),
    .A1(\tms1x00.ins_pla_ors[14][4] ),
    .S(net233),
    .X(_00329_));
 sky130_fd_sc_hd__mux2_1 _07489_ (.A0(_03485_),
    .A1(\tms1x00.ins_pla_ors[14][12] ),
    .S(net231),
    .X(_00330_));
 sky130_fd_sc_hd__mux2_1 _07490_ (.A0(_03487_),
    .A1(\tms1x00.ins_pla_ors[14][13] ),
    .S(net231),
    .X(_00331_));
 sky130_fd_sc_hd__mux2_1 _07491_ (.A0(_03441_),
    .A1(\tms1x00.ins_pla_ors[14][16] ),
    .S(net233),
    .X(_00332_));
 sky130_fd_sc_hd__mux2_1 _07492_ (.A0(_03543_),
    .A1(\tms1x00.ins_pla_ors[14][22] ),
    .S(net232),
    .X(_00333_));
 sky130_fd_sc_hd__a221o_1 _07493_ (.A1(\tms1x00.ins_pla_ors[14][23] ),
    .A2(net232),
    .B1(_03497_),
    .B2(net336),
    .C1(net393),
    .X(_00334_));
 sky130_fd_sc_hd__a221o_1 _07494_ (.A1(\tms1x00.ins_pla_ors[14][25] ),
    .A2(net232),
    .B1(_03498_),
    .B2(net336),
    .C1(net393),
    .X(_00335_));
 sky130_fd_sc_hd__mux2_1 _07495_ (.A0(_03636_),
    .A1(\tms1x00.ins_pla_ors[14][27] ),
    .S(net232),
    .X(_00336_));
 sky130_fd_sc_hd__mux2_1 _07496_ (.A0(_03452_),
    .A1(\tms1x00.ins_pla_ors[14][29] ),
    .S(net232),
    .X(_00337_));
 sky130_fd_sc_hd__or2_1 _07497_ (.A(\tms1x00.ins_pla_ors[2][1] ),
    .B(_03631_),
    .X(_03652_));
 sky130_fd_sc_hd__o211a_1 _07498_ (.A1(net934),
    .A2(net312),
    .B1(_03652_),
    .C1(net485),
    .X(_00338_));
 sky130_fd_sc_hd__or2_1 _07499_ (.A(\tms1x00.ins_pla_ors[2][4] ),
    .B(_03631_),
    .X(_03653_));
 sky130_fd_sc_hd__o211a_1 _07500_ (.A1(net1053),
    .A2(net312),
    .B1(_03653_),
    .C1(net486),
    .X(_00339_));
 sky130_fd_sc_hd__mux2_1 _07501_ (.A0(net1044),
    .A1(\tms1x00.ins_pla_ors[2][5] ),
    .S(net312),
    .X(_03654_));
 sky130_fd_sc_hd__or2_1 _07502_ (.A(net549),
    .B(_03654_),
    .X(_00340_));
 sky130_fd_sc_hd__mux2_1 _07503_ (.A0(net1037),
    .A1(\tms1x00.ins_pla_ors[2][6] ),
    .S(net313),
    .X(_03655_));
 sky130_fd_sc_hd__or2_1 _07504_ (.A(net552),
    .B(_03655_),
    .X(_00341_));
 sky130_fd_sc_hd__mux2_1 _07505_ (.A0(net1029),
    .A1(\tms1x00.ins_pla_ors[2][7] ),
    .S(net312),
    .X(_03656_));
 sky130_fd_sc_hd__or2_1 _07506_ (.A(net554),
    .B(_03656_),
    .X(_00342_));
 sky130_fd_sc_hd__or2_1 _07507_ (.A(\tms1x00.ins_pla_ors[2][9] ),
    .B(_03631_),
    .X(_03657_));
 sky130_fd_sc_hd__o211a_1 _07508_ (.A1(net1013),
    .A2(net313),
    .B1(_03657_),
    .C1(net488),
    .X(_00343_));
 sky130_fd_sc_hd__mux2_1 _07509_ (.A0(net975),
    .A1(\tms1x00.ins_pla_ors[2][10] ),
    .S(net313),
    .X(_03658_));
 sky130_fd_sc_hd__or2_1 _07510_ (.A(net549),
    .B(_03658_),
    .X(_00344_));
 sky130_fd_sc_hd__mux2_1 _07511_ (.A0(net971),
    .A1(\tms1x00.ins_pla_ors[2][11] ),
    .S(net312),
    .X(_03659_));
 sky130_fd_sc_hd__or2_1 _07512_ (.A(net549),
    .B(_03659_),
    .X(_00345_));
 sky130_fd_sc_hd__mux2_1 _07513_ (.A0(net966),
    .A1(\tms1x00.ins_pla_ors[2][12] ),
    .S(net312),
    .X(_03660_));
 sky130_fd_sc_hd__or2_1 _07514_ (.A(net549),
    .B(_03660_),
    .X(_00346_));
 sky130_fd_sc_hd__mux2_1 _07515_ (.A0(net92),
    .A1(\tms1x00.ins_pla_ors[2][13] ),
    .S(net313),
    .X(_03661_));
 sky130_fd_sc_hd__or2_1 _07516_ (.A(net553),
    .B(_03661_),
    .X(_00347_));
 sky130_fd_sc_hd__mux2_1 _07517_ (.A0(net955),
    .A1(\tms1x00.ins_pla_ors[2][14] ),
    .S(net314),
    .X(_03662_));
 sky130_fd_sc_hd__or2_1 _07518_ (.A(net546),
    .B(_03662_),
    .X(_00348_));
 sky130_fd_sc_hd__mux2_1 _07519_ (.A0(net948),
    .A1(\tms1x00.ins_pla_ors[2][15] ),
    .S(net314),
    .X(_03663_));
 sky130_fd_sc_hd__or2_1 _07520_ (.A(net544),
    .B(_03663_),
    .X(_00349_));
 sky130_fd_sc_hd__mux2_1 _07521_ (.A0(net942),
    .A1(\tms1x00.ins_pla_ors[2][16] ),
    .S(net313),
    .X(_03664_));
 sky130_fd_sc_hd__or2_1 _07522_ (.A(net550),
    .B(_03664_),
    .X(_00350_));
 sky130_fd_sc_hd__mux2_1 _07523_ (.A0(net935),
    .A1(\tms1x00.ins_pla_ors[2][19] ),
    .S(net314),
    .X(_03665_));
 sky130_fd_sc_hd__or2_1 _07524_ (.A(net547),
    .B(_03665_),
    .X(_00351_));
 sky130_fd_sc_hd__mux2_1 _07525_ (.A0(net1079),
    .A1(\tms1x00.ins_pla_ors[2][20] ),
    .S(net314),
    .X(_03666_));
 sky130_fd_sc_hd__or2_1 _07526_ (.A(net546),
    .B(_03666_),
    .X(_00352_));
 sky130_fd_sc_hd__mux2_1 _07527_ (.A0(net1077),
    .A1(\tms1x00.ins_pla_ors[2][21] ),
    .S(net314),
    .X(_03667_));
 sky130_fd_sc_hd__or2_1 _07528_ (.A(net544),
    .B(_03667_),
    .X(_00353_));
 sky130_fd_sc_hd__mux2_1 _07529_ (.A0(net1075),
    .A1(\tms1x00.ins_pla_ors[2][22] ),
    .S(net314),
    .X(_03668_));
 sky130_fd_sc_hd__or2_1 _07530_ (.A(net545),
    .B(_03668_),
    .X(_00354_));
 sky130_fd_sc_hd__mux2_1 _07531_ (.A0(net1074),
    .A1(\tms1x00.ins_pla_ors[2][23] ),
    .S(net313),
    .X(_03669_));
 sky130_fd_sc_hd__or2_1 _07532_ (.A(net550),
    .B(_03669_),
    .X(_00355_));
 sky130_fd_sc_hd__mux2_1 _07533_ (.A0(net1073),
    .A1(\tms1x00.ins_pla_ors[2][24] ),
    .S(net313),
    .X(_03670_));
 sky130_fd_sc_hd__or2_1 _07534_ (.A(net551),
    .B(_03670_),
    .X(_00356_));
 sky130_fd_sc_hd__mux2_1 _07535_ (.A0(net105),
    .A1(\tms1x00.ins_pla_ors[2][25] ),
    .S(net314),
    .X(_03671_));
 sky130_fd_sc_hd__or2_1 _07536_ (.A(net544),
    .B(_03671_),
    .X(_00357_));
 sky130_fd_sc_hd__or2_1 _07537_ (.A(\tms1x00.ins_pla_ors[2][29] ),
    .B(_03631_),
    .X(_03672_));
 sky130_fd_sc_hd__o211a_1 _07538_ (.A1(net109),
    .A2(net312),
    .B1(_03672_),
    .C1(net485),
    .X(_00358_));
 sky130_fd_sc_hd__nor2_1 _07539_ (.A(net784),
    .B(net345),
    .Y(_03673_));
 sky130_fd_sc_hd__or2_1 _07540_ (.A(net786),
    .B(net345),
    .X(_03674_));
 sky130_fd_sc_hd__mux2_1 _07541_ (.A0(net982),
    .A1(\tms1x00.ins_pla_ors[7][0] ),
    .S(net304),
    .X(_03675_));
 sky130_fd_sc_hd__or2_1 _07542_ (.A(net572),
    .B(_03675_),
    .X(_00359_));
 sky130_fd_sc_hd__mux2_1 _07543_ (.A0(net934),
    .A1(\tms1x00.ins_pla_ors[7][1] ),
    .S(net302),
    .X(_03676_));
 sky130_fd_sc_hd__or2_1 _07544_ (.A(net568),
    .B(_03676_),
    .X(_00360_));
 sky130_fd_sc_hd__mux2_1 _07545_ (.A0(net1070),
    .A1(\tms1x00.ins_pla_ors[7][2] ),
    .S(net302),
    .X(_03677_));
 sky130_fd_sc_hd__or2_1 _07546_ (.A(net568),
    .B(_03677_),
    .X(_00361_));
 sky130_fd_sc_hd__mux2_1 _07547_ (.A0(net1062),
    .A1(\tms1x00.ins_pla_ors[7][3] ),
    .S(net302),
    .X(_03678_));
 sky130_fd_sc_hd__or2_1 _07548_ (.A(net541),
    .B(_03678_),
    .X(_00362_));
 sky130_fd_sc_hd__mux2_1 _07549_ (.A0(net1053),
    .A1(\tms1x00.ins_pla_ors[7][4] ),
    .S(net304),
    .X(_03679_));
 sky130_fd_sc_hd__or2_1 _07550_ (.A(net568),
    .B(_03679_),
    .X(_00363_));
 sky130_fd_sc_hd__mux2_1 _07551_ (.A0(net1044),
    .A1(\tms1x00.ins_pla_ors[7][5] ),
    .S(net304),
    .X(_03680_));
 sky130_fd_sc_hd__or2_1 _07552_ (.A(net549),
    .B(_03680_),
    .X(_00364_));
 sky130_fd_sc_hd__mux2_1 _07553_ (.A0(net1037),
    .A1(\tms1x00.ins_pla_ors[7][6] ),
    .S(net303),
    .X(_03681_));
 sky130_fd_sc_hd__or2_1 _07554_ (.A(net550),
    .B(_03681_),
    .X(_00365_));
 sky130_fd_sc_hd__mux2_1 _07555_ (.A0(net1027),
    .A1(\tms1x00.ins_pla_ors[7][7] ),
    .S(net305),
    .X(_03682_));
 sky130_fd_sc_hd__or2_1 _07556_ (.A(net567),
    .B(_03682_),
    .X(_00366_));
 sky130_fd_sc_hd__mux2_1 _07557_ (.A0(net1021),
    .A1(\tms1x00.ins_pla_ors[7][8] ),
    .S(net305),
    .X(_03683_));
 sky130_fd_sc_hd__or2_1 _07558_ (.A(net567),
    .B(_03683_),
    .X(_00367_));
 sky130_fd_sc_hd__mux2_1 _07559_ (.A0(net1013),
    .A1(\tms1x00.ins_pla_ors[7][9] ),
    .S(net304),
    .X(_03684_));
 sky130_fd_sc_hd__or2_1 _07560_ (.A(net572),
    .B(_03684_),
    .X(_00368_));
 sky130_fd_sc_hd__mux2_1 _07561_ (.A0(net974),
    .A1(\tms1x00.ins_pla_ors[7][10] ),
    .S(net304),
    .X(_03685_));
 sky130_fd_sc_hd__or2_1 _07562_ (.A(net572),
    .B(_03685_),
    .X(_00369_));
 sky130_fd_sc_hd__mux2_1 _07563_ (.A0(net971),
    .A1(\tms1x00.ins_pla_ors[7][11] ),
    .S(net303),
    .X(_03686_));
 sky130_fd_sc_hd__or2_1 _07564_ (.A(net549),
    .B(_03686_),
    .X(_00370_));
 sky130_fd_sc_hd__mux2_1 _07565_ (.A0(net966),
    .A1(\tms1x00.ins_pla_ors[7][12] ),
    .S(net303),
    .X(_03687_));
 sky130_fd_sc_hd__or2_1 _07566_ (.A(net545),
    .B(_03687_),
    .X(_00371_));
 sky130_fd_sc_hd__mux2_1 _07567_ (.A0(net961),
    .A1(\tms1x00.ins_pla_ors[7][13] ),
    .S(net304),
    .X(_03688_));
 sky130_fd_sc_hd__or2_1 _07568_ (.A(net568),
    .B(_03688_),
    .X(_00372_));
 sky130_fd_sc_hd__mux2_1 _07569_ (.A0(net955),
    .A1(\tms1x00.ins_pla_ors[7][14] ),
    .S(net302),
    .X(_03689_));
 sky130_fd_sc_hd__or2_1 _07570_ (.A(net539),
    .B(_03689_),
    .X(_00373_));
 sky130_fd_sc_hd__mux2_1 _07571_ (.A0(net948),
    .A1(\tms1x00.ins_pla_ors[7][15] ),
    .S(net302),
    .X(_03690_));
 sky130_fd_sc_hd__or2_1 _07572_ (.A(net544),
    .B(_03690_),
    .X(_00374_));
 sky130_fd_sc_hd__mux2_1 _07573_ (.A0(net942),
    .A1(\tms1x00.ins_pla_ors[7][16] ),
    .S(net303),
    .X(_03691_));
 sky130_fd_sc_hd__or2_1 _07574_ (.A(net546),
    .B(_03691_),
    .X(_00375_));
 sky130_fd_sc_hd__mux2_1 _07575_ (.A0(net940),
    .A1(\tms1x00.ins_pla_ors[7][17] ),
    .S(net303),
    .X(_03692_));
 sky130_fd_sc_hd__or2_1 _07576_ (.A(net546),
    .B(_03692_),
    .X(_00376_));
 sky130_fd_sc_hd__mux2_1 _07577_ (.A0(net938),
    .A1(\tms1x00.ins_pla_ors[7][18] ),
    .S(net303),
    .X(_03693_));
 sky130_fd_sc_hd__or2_1 _07578_ (.A(net546),
    .B(_03693_),
    .X(_00377_));
 sky130_fd_sc_hd__mux2_1 _07579_ (.A0(net935),
    .A1(\tms1x00.ins_pla_ors[7][19] ),
    .S(net303),
    .X(_03694_));
 sky130_fd_sc_hd__or2_1 _07580_ (.A(net547),
    .B(_03694_),
    .X(_00378_));
 sky130_fd_sc_hd__mux2_1 _07581_ (.A0(net1079),
    .A1(\tms1x00.ins_pla_ors[7][20] ),
    .S(net303),
    .X(_03695_));
 sky130_fd_sc_hd__or2_1 _07582_ (.A(net546),
    .B(_03695_),
    .X(_00379_));
 sky130_fd_sc_hd__mux2_1 _07583_ (.A0(net1077),
    .A1(\tms1x00.ins_pla_ors[7][21] ),
    .S(net303),
    .X(_03696_));
 sky130_fd_sc_hd__or2_1 _07584_ (.A(net548),
    .B(_03696_),
    .X(_00380_));
 sky130_fd_sc_hd__mux2_1 _07585_ (.A0(net1076),
    .A1(\tms1x00.ins_pla_ors[7][22] ),
    .S(net302),
    .X(_03697_));
 sky130_fd_sc_hd__or2_1 _07586_ (.A(net544),
    .B(_03697_),
    .X(_00381_));
 sky130_fd_sc_hd__mux2_1 _07587_ (.A0(net1074),
    .A1(\tms1x00.ins_pla_ors[7][23] ),
    .S(net304),
    .X(_03698_));
 sky130_fd_sc_hd__or2_1 _07588_ (.A(net550),
    .B(_03698_),
    .X(_00382_));
 sky130_fd_sc_hd__mux2_1 _07589_ (.A0(net1073),
    .A1(\tms1x00.ins_pla_ors[7][24] ),
    .S(net304),
    .X(_03699_));
 sky130_fd_sc_hd__or2_1 _07590_ (.A(net552),
    .B(_03699_),
    .X(_00383_));
 sky130_fd_sc_hd__mux2_1 _07591_ (.A0(net105),
    .A1(\tms1x00.ins_pla_ors[7][25] ),
    .S(net302),
    .X(_03700_));
 sky130_fd_sc_hd__or2_1 _07592_ (.A(net539),
    .B(_03700_),
    .X(_00384_));
 sky130_fd_sc_hd__mux2_1 _07593_ (.A0(net1072),
    .A1(\tms1x00.ins_pla_ors[7][26] ),
    .S(net303),
    .X(_03701_));
 sky130_fd_sc_hd__or2_1 _07594_ (.A(net547),
    .B(_03701_),
    .X(_00385_));
 sky130_fd_sc_hd__and3_2 _07595_ (.A(net904),
    .B(net352),
    .C(net708),
    .X(_03702_));
 sky130_fd_sc_hd__or3_4 _07596_ (.A(net896),
    .B(net349),
    .C(net706),
    .X(_03703_));
 sky130_fd_sc_hd__nor2_2 _07597_ (.A(net382),
    .B(_03702_),
    .Y(_03704_));
 sky130_fd_sc_hd__nand2_2 _07598_ (.A(net373),
    .B(_03703_),
    .Y(_03705_));
 sky130_fd_sc_hd__nor2_2 _07599_ (.A(net396),
    .B(_03702_),
    .Y(_03706_));
 sky130_fd_sc_hd__nand2_2 _07600_ (.A(net385),
    .B(_03703_),
    .Y(_03707_));
 sky130_fd_sc_hd__a22o_1 _07601_ (.A1(\tms1x00.ins_pla_ands[5][0] ),
    .A2(_03704_),
    .B1(_03707_),
    .B2(net343),
    .X(_00386_));
 sky130_fd_sc_hd__o22a_1 _07602_ (.A1(\tms1x00.ins_pla_ands[5][1] ),
    .A2(_03705_),
    .B1(_03706_),
    .B2(net344),
    .X(_00387_));
 sky130_fd_sc_hd__a22o_1 _07603_ (.A1(\tms1x00.ins_pla_ands[5][2] ),
    .A2(_03704_),
    .B1(_03707_),
    .B2(_03429_),
    .X(_00388_));
 sky130_fd_sc_hd__o22a_1 _07604_ (.A1(\tms1x00.ins_pla_ands[5][3] ),
    .A2(_03705_),
    .B1(_03706_),
    .B2(_03433_),
    .X(_00389_));
 sky130_fd_sc_hd__a22o_1 _07605_ (.A1(\tms1x00.ins_pla_ands[5][6] ),
    .A2(_03704_),
    .B1(_03707_),
    .B2(_03435_),
    .X(_00390_));
 sky130_fd_sc_hd__o22a_1 _07606_ (.A1(\tms1x00.ins_pla_ands[5][7] ),
    .A2(_03705_),
    .B1(_03706_),
    .B2(_03536_),
    .X(_00391_));
 sky130_fd_sc_hd__a22o_1 _07607_ (.A1(\tms1x00.ins_pla_ands[5][8] ),
    .A2(_03704_),
    .B1(_03707_),
    .B2(_03439_),
    .X(_00392_));
 sky130_fd_sc_hd__o22a_1 _07608_ (.A1(\tms1x00.ins_pla_ands[5][9] ),
    .A2(_03705_),
    .B1(_03706_),
    .B2(_03578_),
    .X(_00393_));
 sky130_fd_sc_hd__a22o_1 _07609_ (.A1(\tms1x00.ins_pla_ands[5][10] ),
    .A2(_03704_),
    .B1(_03707_),
    .B2(_03579_),
    .X(_00394_));
 sky130_fd_sc_hd__o22a_1 _07610_ (.A1(\tms1x00.ins_pla_ands[5][11] ),
    .A2(_03705_),
    .B1(_03706_),
    .B2(_03580_),
    .X(_00395_));
 sky130_fd_sc_hd__and3_4 _07611_ (.A(net822),
    .B(net352),
    .C(net708),
    .X(_03708_));
 sky130_fd_sc_hd__or3_4 _07612_ (.A(net813),
    .B(_03470_),
    .C(net706),
    .X(_03709_));
 sky130_fd_sc_hd__nor2_2 _07613_ (.A(net382),
    .B(_03708_),
    .Y(_03710_));
 sky130_fd_sc_hd__nand2_2 _07614_ (.A(net388),
    .B(net301),
    .Y(_03711_));
 sky130_fd_sc_hd__a22o_1 _07615_ (.A1(\tms1x00.ins_pla_ands[4][0] ),
    .A2(_03710_),
    .B1(_03711_),
    .B2(_03585_),
    .X(_00396_));
 sky130_fd_sc_hd__a22o_1 _07616_ (.A1(\tms1x00.ins_pla_ands[4][3] ),
    .A2(_03710_),
    .B1(_03711_),
    .B2(_03534_),
    .X(_00397_));
 sky130_fd_sc_hd__or2_4 _07617_ (.A(net390),
    .B(net366),
    .X(_03712_));
 sky130_fd_sc_hd__a22o_1 _07618_ (.A1(\tms1x00.ins_pla_ands[4][5] ),
    .A2(_03710_),
    .B1(_03711_),
    .B2(_03712_),
    .X(_00398_));
 sky130_fd_sc_hd__a22o_1 _07619_ (.A1(\tms1x00.ins_pla_ands[4][6] ),
    .A2(_03710_),
    .B1(_03711_),
    .B2(_03435_),
    .X(_00399_));
 sky130_fd_sc_hd__a22o_1 _07620_ (.A1(\tms1x00.ins_pla_ands[4][12] ),
    .A2(_03710_),
    .B1(_03711_),
    .B2(_03588_),
    .X(_00400_));
 sky130_fd_sc_hd__a21o_1 _07621_ (.A1(net385),
    .A2(net301),
    .B1(_03589_),
    .X(_03713_));
 sky130_fd_sc_hd__o31a_1 _07622_ (.A1(\tms1x00.ins_pla_ands[4][13] ),
    .A2(net382),
    .A3(_03708_),
    .B1(_03713_),
    .X(_00401_));
 sky130_fd_sc_hd__and3_2 _07623_ (.A(net820),
    .B(net350),
    .C(_03471_),
    .X(_03714_));
 sky130_fd_sc_hd__nor2_1 _07624_ (.A(net512),
    .B(net300),
    .Y(_03715_));
 sky130_fd_sc_hd__mux2_1 _07625_ (.A0(_03481_),
    .A1(\tms1x00.ins_pla_ands[28][9] ),
    .S(net216),
    .X(_00402_));
 sky130_fd_sc_hd__mux2_1 _07626_ (.A0(_03579_),
    .A1(\tms1x00.ins_pla_ands[28][10] ),
    .S(net217),
    .X(_00403_));
 sky130_fd_sc_hd__mux2_1 _07627_ (.A0(_03487_),
    .A1(\tms1x00.ins_pla_ands[28][13] ),
    .S(net216),
    .X(_00404_));
 sky130_fd_sc_hd__mux2_1 _07628_ (.A0(_03537_),
    .A1(\tms1x00.ins_pla_ands[28][14] ),
    .S(net216),
    .X(_00405_));
 sky130_fd_sc_hd__and3_2 _07629_ (.A(net847),
    .B(net350),
    .C(_03471_),
    .X(_03716_));
 sky130_fd_sc_hd__nor2_2 _07630_ (.A(net511),
    .B(_03716_),
    .Y(_03717_));
 sky130_fd_sc_hd__or2_4 _07631_ (.A(net518),
    .B(net299),
    .X(_03718_));
 sky130_fd_sc_hd__mux2_1 _07632_ (.A0(\tms1x00.ins_pla_ands[24][0] ),
    .A1(_03476_),
    .S(_03718_),
    .X(_00406_));
 sky130_fd_sc_hd__mux2_1 _07633_ (.A0(\tms1x00.ins_pla_ands[24][1] ),
    .A1(net354),
    .S(_03718_),
    .X(_00407_));
 sky130_fd_sc_hd__mux2_1 _07634_ (.A0(\tms1x00.ins_pla_ands[24][2] ),
    .A1(_03429_),
    .S(_03718_),
    .X(_00408_));
 sky130_fd_sc_hd__mux2_1 _07635_ (.A0(\tms1x00.ins_pla_ands[24][3] ),
    .A1(_03433_),
    .S(_03718_),
    .X(_00409_));
 sky130_fd_sc_hd__mux2_1 _07636_ (.A0(\tms1x00.ins_pla_ands[24][10] ),
    .A1(_03482_),
    .S(_03718_),
    .X(_00410_));
 sky130_fd_sc_hd__mux2_1 _07637_ (.A0(\tms1x00.ins_pla_ands[24][11] ),
    .A1(net347),
    .S(_03718_),
    .X(_00411_));
 sky130_fd_sc_hd__and3_1 _07638_ (.A(net902),
    .B(net598),
    .C(net350),
    .X(_03719_));
 sky130_fd_sc_hd__nor2_8 _07639_ (.A(net511),
    .B(net298),
    .Y(_03720_));
 sky130_fd_sc_hd__mux2_1 _07640_ (.A0(net343),
    .A1(\tms1x00.ins_pla_ands[21][0] ),
    .S(_03720_),
    .X(_00412_));
 sky130_fd_sc_hd__mux2_1 _07641_ (.A0(net344),
    .A1(\tms1x00.ins_pla_ands[21][1] ),
    .S(_03720_),
    .X(_00413_));
 sky130_fd_sc_hd__mux2_1 _07642_ (.A0(net347),
    .A1(\tms1x00.ins_pla_ands[21][11] ),
    .S(_03720_),
    .X(_00414_));
 sky130_fd_sc_hd__and3_2 _07643_ (.A(net820),
    .B(net598),
    .C(_03469_),
    .X(_03721_));
 sky130_fd_sc_hd__nor2_2 _07644_ (.A(net513),
    .B(net296),
    .Y(_03722_));
 sky130_fd_sc_hd__or2_4 _07645_ (.A(net517),
    .B(_03721_),
    .X(_03723_));
 sky130_fd_sc_hd__mux2_1 _07646_ (.A0(\tms1x00.ins_pla_ands[20][0] ),
    .A1(_03476_),
    .S(_03723_),
    .X(_00415_));
 sky130_fd_sc_hd__mux2_1 _07647_ (.A0(\tms1x00.ins_pla_ands[20][1] ),
    .A1(net354),
    .S(_03723_),
    .X(_00416_));
 sky130_fd_sc_hd__mux2_1 _07648_ (.A0(\tms1x00.ins_pla_ands[20][2] ),
    .A1(_03429_),
    .S(_03723_),
    .X(_00417_));
 sky130_fd_sc_hd__mux2_1 _07649_ (.A0(\tms1x00.ins_pla_ands[20][3] ),
    .A1(_03433_),
    .S(_03723_),
    .X(_00418_));
 sky130_fd_sc_hd__mux2_1 _07650_ (.A0(\tms1x00.ins_pla_ands[20][10] ),
    .A1(_03482_),
    .S(_03723_),
    .X(_00419_));
 sky130_fd_sc_hd__mux2_1 _07651_ (.A0(\tms1x00.ins_pla_ands[20][11] ),
    .A1(net347),
    .S(_03723_),
    .X(_00420_));
 sky130_fd_sc_hd__mux2_1 _07652_ (.A0(net343),
    .A1(\tms1x00.ins_pla_ands[19][0] ),
    .S(_03601_),
    .X(_00421_));
 sky130_fd_sc_hd__mux2_1 _07653_ (.A0(net344),
    .A1(\tms1x00.ins_pla_ands[19][1] ),
    .S(_03601_),
    .X(_00422_));
 sky130_fd_sc_hd__mux2_1 _07654_ (.A0(_03482_),
    .A1(\tms1x00.ins_pla_ands[19][10] ),
    .S(_03601_),
    .X(_00423_));
 sky130_fd_sc_hd__mux2_1 _07655_ (.A0(net347),
    .A1(\tms1x00.ins_pla_ands[19][11] ),
    .S(_03601_),
    .X(_00424_));
 sky130_fd_sc_hd__o22a_1 _07656_ (.A1(\tms1x00.ins_pla_ors[11][2] ),
    .A2(net323),
    .B1(net222),
    .B2(_03428_),
    .X(_00425_));
 sky130_fd_sc_hd__o22a_1 _07657_ (.A1(\tms1x00.ins_pla_ors[11][5] ),
    .A2(net323),
    .B1(net222),
    .B2(_03457_),
    .X(_00426_));
 sky130_fd_sc_hd__mux2_1 _07658_ (.A0(\tms1x00.ins_pla_ors[11][8] ),
    .A1(net1022),
    .S(net323),
    .X(_03724_));
 sky130_fd_sc_hd__or2_1 _07659_ (.A(net525),
    .B(_03724_),
    .X(_00427_));
 sky130_fd_sc_hd__o22a_1 _07660_ (.A1(\tms1x00.ins_pla_ors[11][9] ),
    .A2(net323),
    .B1(net222),
    .B2(net365),
    .X(_00428_));
 sky130_fd_sc_hd__o22a_1 _07661_ (.A1(\tms1x00.ins_pla_ors[11][10] ),
    .A2(net323),
    .B1(net222),
    .B2(_03459_),
    .X(_00429_));
 sky130_fd_sc_hd__o22a_1 _07662_ (.A1(\tms1x00.ins_pla_ors[11][11] ),
    .A2(net323),
    .B1(net224),
    .B2(_03460_),
    .X(_00430_));
 sky130_fd_sc_hd__mux2_1 _07663_ (.A0(\tms1x00.ins_pla_ors[11][12] ),
    .A1(net965),
    .S(net323),
    .X(_03725_));
 sky130_fd_sc_hd__or2_1 _07664_ (.A(net522),
    .B(_03725_),
    .X(_00431_));
 sky130_fd_sc_hd__mux2_1 _07665_ (.A0(\tms1x00.ins_pla_ors[11][20] ),
    .A1(net1078),
    .S(net324),
    .X(_03726_));
 sky130_fd_sc_hd__or2_1 _07666_ (.A(net538),
    .B(_03726_),
    .X(_00432_));
 sky130_fd_sc_hd__o22a_1 _07667_ (.A1(\tms1x00.ins_pla_ors[11][23] ),
    .A2(net324),
    .B1(net223),
    .B2(_03497_),
    .X(_00433_));
 sky130_fd_sc_hd__o22a_1 _07668_ (.A1(\tms1x00.ins_pla_ors[11][24] ),
    .A2(net324),
    .B1(net224),
    .B2(_03467_),
    .X(_00434_));
 sky130_fd_sc_hd__o22a_1 _07669_ (.A1(\tms1x00.ins_pla_ors[11][27] ),
    .A2(net324),
    .B1(net223),
    .B2(_03500_),
    .X(_00435_));
 sky130_fd_sc_hd__o22a_1 _07670_ (.A1(\tms1x00.ins_pla_ors[11][28] ),
    .A2(net324),
    .B1(net223),
    .B2(_03449_),
    .X(_00436_));
 sky130_fd_sc_hd__o22a_1 _07671_ (.A1(\tms1x00.ins_pla_ors[11][29] ),
    .A2(net324),
    .B1(net223),
    .B2(_03451_),
    .X(_00437_));
 sky130_fd_sc_hd__and3_4 _07672_ (.A(net795),
    .B(net351),
    .C(net708),
    .X(_03727_));
 sky130_fd_sc_hd__nor2_4 _07673_ (.A(net376),
    .B(_03727_),
    .Y(_03728_));
 sky130_fd_sc_hd__or2_4 _07674_ (.A(net376),
    .B(_03727_),
    .X(_03729_));
 sky130_fd_sc_hd__nor2_2 _07675_ (.A(net391),
    .B(_03727_),
    .Y(_03730_));
 sky130_fd_sc_hd__or2_4 _07676_ (.A(net392),
    .B(_03727_),
    .X(_03731_));
 sky130_fd_sc_hd__a22o_1 _07677_ (.A1(\tms1x00.ins_pla_ands[7][0] ),
    .A2(_03728_),
    .B1(_03731_),
    .B2(net343),
    .X(_00438_));
 sky130_fd_sc_hd__o22a_1 _07678_ (.A1(\tms1x00.ins_pla_ands[7][1] ),
    .A2(_03729_),
    .B1(_03730_),
    .B2(_03533_),
    .X(_00439_));
 sky130_fd_sc_hd__o22a_1 _07679_ (.A1(\tms1x00.ins_pla_ands[7][2] ),
    .A2(_03729_),
    .B1(_03730_),
    .B2(_03477_),
    .X(_00440_));
 sky130_fd_sc_hd__a22o_1 _07680_ (.A1(\tms1x00.ins_pla_ands[7][3] ),
    .A2(_03728_),
    .B1(_03731_),
    .B2(_03534_),
    .X(_00441_));
 sky130_fd_sc_hd__a22o_1 _07681_ (.A1(\tms1x00.ins_pla_ands[7][4] ),
    .A2(_03728_),
    .B1(_03731_),
    .B2(_03535_),
    .X(_00442_));
 sky130_fd_sc_hd__o22a_1 _07682_ (.A1(\tms1x00.ins_pla_ands[7][5] ),
    .A2(_03729_),
    .B1(_03730_),
    .B2(_03577_),
    .X(_00443_));
 sky130_fd_sc_hd__a22o_1 _07683_ (.A1(\tms1x00.ins_pla_ands[7][6] ),
    .A2(_03728_),
    .B1(_03731_),
    .B2(_03435_),
    .X(_00444_));
 sky130_fd_sc_hd__o22a_1 _07684_ (.A1(\tms1x00.ins_pla_ands[7][7] ),
    .A2(_03729_),
    .B1(_03730_),
    .B2(_03536_),
    .X(_00445_));
 sky130_fd_sc_hd__a22o_1 _07685_ (.A1(\tms1x00.ins_pla_ands[7][8] ),
    .A2(_03728_),
    .B1(_03731_),
    .B2(net353),
    .X(_00446_));
 sky130_fd_sc_hd__o22a_1 _07686_ (.A1(\tms1x00.ins_pla_ands[7][9] ),
    .A2(_03729_),
    .B1(_03730_),
    .B2(_03578_),
    .X(_00447_));
 sky130_fd_sc_hd__a22o_1 _07687_ (.A1(\tms1x00.ins_pla_ands[7][10] ),
    .A2(_03728_),
    .B1(_03731_),
    .B2(_03579_),
    .X(_00448_));
 sky130_fd_sc_hd__o22a_1 _07688_ (.A1(\tms1x00.ins_pla_ands[7][11] ),
    .A2(_03729_),
    .B1(_03730_),
    .B2(_03580_),
    .X(_00449_));
 sky130_fd_sc_hd__nor2_8 _07689_ (.A(net987),
    .B(net917),
    .Y(_03732_));
 sky130_fd_sc_hd__nand2_8 _07690_ (.A(net925),
    .B(net994),
    .Y(_03733_));
 sky130_fd_sc_hd__and3_4 _07691_ (.A(net847),
    .B(net351),
    .C(net596),
    .X(_03734_));
 sky130_fd_sc_hd__or3_4 _07692_ (.A(net829),
    .B(net349),
    .C(net594),
    .X(_03735_));
 sky130_fd_sc_hd__nor2_2 _07693_ (.A(net376),
    .B(_03734_),
    .Y(_03736_));
 sky130_fd_sc_hd__nand2_2 _07694_ (.A(net370),
    .B(_03735_),
    .Y(_03737_));
 sky130_fd_sc_hd__o221a_1 _07695_ (.A1(_03574_),
    .A2(_03735_),
    .B1(_03737_),
    .B2(\tms1x00.ins_pla_ands[8][0] ),
    .C1(net383),
    .X(_00450_));
 sky130_fd_sc_hd__nor2_2 _07696_ (.A(net391),
    .B(_03734_),
    .Y(_03738_));
 sky130_fd_sc_hd__nand2_2 _07697_ (.A(net384),
    .B(_03735_),
    .Y(_03739_));
 sky130_fd_sc_hd__a22o_1 _07698_ (.A1(\tms1x00.ins_pla_ands[8][1] ),
    .A2(_03736_),
    .B1(_03739_),
    .B2(net354),
    .X(_00451_));
 sky130_fd_sc_hd__o22a_1 _07699_ (.A1(\tms1x00.ins_pla_ands[8][5] ),
    .A2(_03737_),
    .B1(_03738_),
    .B2(_03577_),
    .X(_00452_));
 sky130_fd_sc_hd__a22o_1 _07700_ (.A1(\tms1x00.ins_pla_ands[8][6] ),
    .A2(_03736_),
    .B1(_03739_),
    .B2(_03435_),
    .X(_00453_));
 sky130_fd_sc_hd__o22a_1 _07701_ (.A1(\tms1x00.ins_pla_ands[8][7] ),
    .A2(_03737_),
    .B1(_03738_),
    .B2(_03536_),
    .X(_00454_));
 sky130_fd_sc_hd__a22o_1 _07702_ (.A1(\tms1x00.ins_pla_ands[8][8] ),
    .A2(_03736_),
    .B1(_03739_),
    .B2(net353),
    .X(_00455_));
 sky130_fd_sc_hd__o22a_1 _07703_ (.A1(\tms1x00.ins_pla_ands[8][9] ),
    .A2(_03737_),
    .B1(_03738_),
    .B2(_03578_),
    .X(_00456_));
 sky130_fd_sc_hd__a22o_1 _07704_ (.A1(\tms1x00.ins_pla_ands[8][10] ),
    .A2(_03736_),
    .B1(_03739_),
    .B2(_03579_),
    .X(_00457_));
 sky130_fd_sc_hd__o22a_1 _07705_ (.A1(\tms1x00.ins_pla_ands[8][11] ),
    .A2(_03737_),
    .B1(_03738_),
    .B2(_03580_),
    .X(_00458_));
 sky130_fd_sc_hd__or2_1 _07706_ (.A(\tms1x00.ins_pla_ors[1][0] ),
    .B(net310),
    .X(_03740_));
 sky130_fd_sc_hd__o211a_1 _07707_ (.A1(net982),
    .A2(net307),
    .B1(_03740_),
    .C1(net486),
    .X(_00459_));
 sky130_fd_sc_hd__or2_1 _07708_ (.A(\tms1x00.ins_pla_ors[1][1] ),
    .B(net311),
    .X(_03741_));
 sky130_fd_sc_hd__o211a_1 _07709_ (.A1(net934),
    .A2(net308),
    .B1(_03741_),
    .C1(net485),
    .X(_00460_));
 sky130_fd_sc_hd__or2_1 _07710_ (.A(\tms1x00.ins_pla_ors[1][3] ),
    .B(net311),
    .X(_03742_));
 sky130_fd_sc_hd__o211a_1 _07711_ (.A1(net1062),
    .A2(net308),
    .B1(_03742_),
    .C1(net488),
    .X(_00461_));
 sky130_fd_sc_hd__or2_1 _07712_ (.A(\tms1x00.ins_pla_ors[1][4] ),
    .B(net311),
    .X(_03743_));
 sky130_fd_sc_hd__o211a_1 _07713_ (.A1(net1053),
    .A2(net308),
    .B1(_03743_),
    .C1(net485),
    .X(_00462_));
 sky130_fd_sc_hd__or2_1 _07714_ (.A(\tms1x00.ins_pla_ors[1][5] ),
    .B(net310),
    .X(_03744_));
 sky130_fd_sc_hd__o211a_1 _07715_ (.A1(net1044),
    .A2(net307),
    .B1(_03744_),
    .C1(net487),
    .X(_00463_));
 sky130_fd_sc_hd__or2_1 _07716_ (.A(\tms1x00.ins_pla_ors[1][6] ),
    .B(net310),
    .X(_03745_));
 sky130_fd_sc_hd__o211a_1 _07717_ (.A1(net1037),
    .A2(net307),
    .B1(_03745_),
    .C1(net486),
    .X(_00464_));
 sky130_fd_sc_hd__or2_1 _07718_ (.A(\tms1x00.ins_pla_ors[1][7] ),
    .B(net311),
    .X(_03746_));
 sky130_fd_sc_hd__o211a_1 _07719_ (.A1(net1029),
    .A2(net308),
    .B1(_03746_),
    .C1(net485),
    .X(_00465_));
 sky130_fd_sc_hd__or2_1 _07720_ (.A(\tms1x00.ins_pla_ors[1][8] ),
    .B(net311),
    .X(_03747_));
 sky130_fd_sc_hd__o211a_1 _07721_ (.A1(net1022),
    .A2(net308),
    .B1(_03747_),
    .C1(net485),
    .X(_00466_));
 sky130_fd_sc_hd__or2_1 _07722_ (.A(\tms1x00.ins_pla_ors[1][9] ),
    .B(net310),
    .X(_03748_));
 sky130_fd_sc_hd__o211a_1 _07723_ (.A1(net1013),
    .A2(net307),
    .B1(_03748_),
    .C1(net487),
    .X(_00467_));
 sky130_fd_sc_hd__or2_1 _07724_ (.A(\tms1x00.ins_pla_ors[1][10] ),
    .B(net309),
    .X(_03749_));
 sky130_fd_sc_hd__o211a_1 _07725_ (.A1(net975),
    .A2(net307),
    .B1(_03749_),
    .C1(net484),
    .X(_00468_));
 sky130_fd_sc_hd__or2_1 _07726_ (.A(\tms1x00.ins_pla_ors[1][11] ),
    .B(net311),
    .X(_03750_));
 sky130_fd_sc_hd__o211a_1 _07727_ (.A1(net970),
    .A2(net308),
    .B1(_03750_),
    .C1(net481),
    .X(_00469_));
 sky130_fd_sc_hd__or2_1 _07728_ (.A(\tms1x00.ins_pla_ors[1][12] ),
    .B(net309),
    .X(_03751_));
 sky130_fd_sc_hd__o211a_1 _07729_ (.A1(net966),
    .A2(net306),
    .B1(_03751_),
    .C1(net482),
    .X(_00470_));
 sky130_fd_sc_hd__or2_1 _07730_ (.A(\tms1x00.ins_pla_ors[1][13] ),
    .B(net310),
    .X(_03752_));
 sky130_fd_sc_hd__o211a_1 _07731_ (.A1(net961),
    .A2(net307),
    .B1(_03752_),
    .C1(net486),
    .X(_00471_));
 sky130_fd_sc_hd__or2_1 _07732_ (.A(\tms1x00.ins_pla_ors[1][14] ),
    .B(net310),
    .X(_03753_));
 sky130_fd_sc_hd__o211a_1 _07733_ (.A1(net955),
    .A2(net306),
    .B1(_03753_),
    .C1(net483),
    .X(_00472_));
 sky130_fd_sc_hd__or2_1 _07734_ (.A(\tms1x00.ins_pla_ors[1][15] ),
    .B(net309),
    .X(_03754_));
 sky130_fd_sc_hd__o211a_1 _07735_ (.A1(net950),
    .A2(net306),
    .B1(_03754_),
    .C1(net484),
    .X(_00473_));
 sky130_fd_sc_hd__or2_1 _07736_ (.A(\tms1x00.ins_pla_ors[1][16] ),
    .B(net310),
    .X(_03755_));
 sky130_fd_sc_hd__o211a_1 _07737_ (.A1(net942),
    .A2(net306),
    .B1(_03755_),
    .C1(net484),
    .X(_00474_));
 sky130_fd_sc_hd__or2_1 _07738_ (.A(\tms1x00.ins_pla_ors[1][17] ),
    .B(net309),
    .X(_03756_));
 sky130_fd_sc_hd__o211a_1 _07739_ (.A1(net940),
    .A2(net306),
    .B1(_03756_),
    .C1(net484),
    .X(_00475_));
 sky130_fd_sc_hd__or2_1 _07740_ (.A(\tms1x00.ins_pla_ors[1][18] ),
    .B(net310),
    .X(_03757_));
 sky130_fd_sc_hd__o211a_1 _07741_ (.A1(net939),
    .A2(net307),
    .B1(_03757_),
    .C1(net487),
    .X(_00476_));
 sky130_fd_sc_hd__or2_1 _07742_ (.A(\tms1x00.ins_pla_ors[1][19] ),
    .B(net309),
    .X(_03758_));
 sky130_fd_sc_hd__o211a_1 _07743_ (.A1(net935),
    .A2(net306),
    .B1(_03758_),
    .C1(net483),
    .X(_00477_));
 sky130_fd_sc_hd__or2_1 _07744_ (.A(\tms1x00.ins_pla_ors[1][20] ),
    .B(net309),
    .X(_03759_));
 sky130_fd_sc_hd__o211a_1 _07745_ (.A1(net1079),
    .A2(net306),
    .B1(_03759_),
    .C1(net483),
    .X(_00478_));
 sky130_fd_sc_hd__or2_1 _07746_ (.A(\tms1x00.ins_pla_ors[1][21] ),
    .B(net309),
    .X(_03760_));
 sky130_fd_sc_hd__o211a_1 _07747_ (.A1(net1077),
    .A2(net307),
    .B1(_03760_),
    .C1(net484),
    .X(_00479_));
 sky130_fd_sc_hd__or2_1 _07748_ (.A(\tms1x00.ins_pla_ors[1][22] ),
    .B(net311),
    .X(_03761_));
 sky130_fd_sc_hd__o211a_1 _07749_ (.A1(net1076),
    .A2(net308),
    .B1(_03761_),
    .C1(net482),
    .X(_00480_));
 sky130_fd_sc_hd__or2_1 _07750_ (.A(\tms1x00.ins_pla_ors[1][23] ),
    .B(net310),
    .X(_03762_));
 sky130_fd_sc_hd__o211a_1 _07751_ (.A1(net1074),
    .A2(net307),
    .B1(_03762_),
    .C1(net487),
    .X(_00481_));
 sky130_fd_sc_hd__or2_1 _07752_ (.A(\tms1x00.ins_pla_ors[1][24] ),
    .B(_03637_),
    .X(_03763_));
 sky130_fd_sc_hd__o211a_1 _07753_ (.A1(net1073),
    .A2(_03638_),
    .B1(_03763_),
    .C1(net486),
    .X(_00482_));
 sky130_fd_sc_hd__or2_1 _07754_ (.A(\tms1x00.ins_pla_ors[1][25] ),
    .B(net311),
    .X(_03764_));
 sky130_fd_sc_hd__o211a_1 _07755_ (.A1(net105),
    .A2(net308),
    .B1(_03764_),
    .C1(net485),
    .X(_00483_));
 sky130_fd_sc_hd__or2_1 _07756_ (.A(\tms1x00.ins_pla_ors[1][26] ),
    .B(net309),
    .X(_03765_));
 sky130_fd_sc_hd__o211a_1 _07757_ (.A1(net1072),
    .A2(net306),
    .B1(_03765_),
    .C1(net484),
    .X(_00484_));
 sky130_fd_sc_hd__or2_1 _07758_ (.A(\tms1x00.ins_pla_ors[1][28] ),
    .B(net309),
    .X(_03766_));
 sky130_fd_sc_hd__o211a_1 _07759_ (.A1(net108),
    .A2(net306),
    .B1(_03766_),
    .C1(net484),
    .X(_00485_));
 sky130_fd_sc_hd__or2_1 _07760_ (.A(\tms1x00.ins_pla_ors[1][29] ),
    .B(net309),
    .X(_03767_));
 sky130_fd_sc_hd__o211a_1 _07761_ (.A1(net109),
    .A2(net306),
    .B1(_03767_),
    .C1(net483),
    .X(_00486_));
 sky130_fd_sc_hd__mux2_1 _07762_ (.A0(\tms1x00.ins_pla_ors[13][1] ),
    .A1(net344),
    .S(net225),
    .X(_00487_));
 sky130_fd_sc_hd__mux2_1 _07763_ (.A0(\tms1x00.ins_pla_ors[13][2] ),
    .A1(_03429_),
    .S(net226),
    .X(_00488_));
 sky130_fd_sc_hd__mux2_1 _07764_ (.A0(\tms1x00.ins_pla_ors[13][3] ),
    .A1(_03534_),
    .S(net225),
    .X(_00489_));
 sky130_fd_sc_hd__mux2_1 _07765_ (.A0(\tms1x00.ins_pla_ors[13][4] ),
    .A1(_03535_),
    .S(net225),
    .X(_00490_));
 sky130_fd_sc_hd__mux2_1 _07766_ (.A0(\tms1x00.ins_pla_ors[13][5] ),
    .A1(_03712_),
    .S(net226),
    .X(_00491_));
 sky130_fd_sc_hd__mux2_1 _07767_ (.A0(\tms1x00.ins_pla_ors[13][6] ),
    .A1(_03480_),
    .S(net226),
    .X(_00492_));
 sky130_fd_sc_hd__mux2_1 _07768_ (.A0(\tms1x00.ins_pla_ors[13][7] ),
    .A1(_03536_),
    .S(net225),
    .X(_00493_));
 sky130_fd_sc_hd__mux2_1 _07769_ (.A0(\tms1x00.ins_pla_ors[13][10] ),
    .A1(_03579_),
    .S(net225),
    .X(_00494_));
 sky130_fd_sc_hd__a221o_1 _07770_ (.A1(_03484_),
    .A2(net325),
    .B1(net227),
    .B2(\tms1x00.ins_pla_ors[13][12] ),
    .C1(net389),
    .X(_00495_));
 sky130_fd_sc_hd__a221o_1 _07771_ (.A1(_03486_),
    .A2(net325),
    .B1(net227),
    .B2(\tms1x00.ins_pla_ors[13][13] ),
    .C1(net375),
    .X(_00496_));
 sky130_fd_sc_hd__mux2_1 _07772_ (.A0(\tms1x00.ins_pla_ors[13][17] ),
    .A1(_03540_),
    .S(net226),
    .X(_00497_));
 sky130_fd_sc_hd__mux2_1 _07773_ (.A0(\tms1x00.ins_pla_ors[13][19] ),
    .A1(_03542_),
    .S(net225),
    .X(_00498_));
 sky130_fd_sc_hd__a221o_1 _07774_ (.A1(net1075),
    .A2(net326),
    .B1(_03528_),
    .B2(\tms1x00.ins_pla_ors[13][22] ),
    .C1(net393),
    .X(_00499_));
 sky130_fd_sc_hd__a221o_1 _07775_ (.A1(_03497_),
    .A2(net326),
    .B1(_03528_),
    .B2(\tms1x00.ins_pla_ors[13][23] ),
    .C1(net381),
    .X(_00500_));
 sky130_fd_sc_hd__a221o_1 _07776_ (.A1(net1073),
    .A2(net326),
    .B1(_03528_),
    .B2(\tms1x00.ins_pla_ors[13][24] ),
    .C1(net395),
    .X(_00501_));
 sky130_fd_sc_hd__nor2_2 _07777_ (.A(net618),
    .B(net345),
    .Y(_03768_));
 sky130_fd_sc_hd__or2_1 _07778_ (.A(net619),
    .B(net346),
    .X(_03769_));
 sky130_fd_sc_hd__mux2_1 _07779_ (.A0(net982),
    .A1(\tms1x00.ins_pla_ors[6][0] ),
    .S(net294),
    .X(_03770_));
 sky130_fd_sc_hd__or2_1 _07780_ (.A(net552),
    .B(_03770_),
    .X(_00502_));
 sky130_fd_sc_hd__mux2_1 _07781_ (.A0(net934),
    .A1(\tms1x00.ins_pla_ors[6][1] ),
    .S(net294),
    .X(_03771_));
 sky130_fd_sc_hd__or2_1 _07782_ (.A(net567),
    .B(_03771_),
    .X(_00503_));
 sky130_fd_sc_hd__mux2_1 _07783_ (.A0(net1070),
    .A1(\tms1x00.ins_pla_ors[6][2] ),
    .S(net294),
    .X(_03772_));
 sky130_fd_sc_hd__or2_1 _07784_ (.A(net567),
    .B(_03772_),
    .X(_00504_));
 sky130_fd_sc_hd__mux2_1 _07785_ (.A0(net1062),
    .A1(\tms1x00.ins_pla_ors[6][3] ),
    .S(net294),
    .X(_03773_));
 sky130_fd_sc_hd__or2_1 _07786_ (.A(net541),
    .B(_03773_),
    .X(_00505_));
 sky130_fd_sc_hd__mux2_1 _07787_ (.A0(net1053),
    .A1(\tms1x00.ins_pla_ors[6][4] ),
    .S(net294),
    .X(_03774_));
 sky130_fd_sc_hd__or2_1 _07788_ (.A(net568),
    .B(_03774_),
    .X(_00506_));
 sky130_fd_sc_hd__mux2_1 _07789_ (.A0(net1044),
    .A1(\tms1x00.ins_pla_ors[6][5] ),
    .S(net294),
    .X(_03775_));
 sky130_fd_sc_hd__or2_1 _07790_ (.A(net554),
    .B(_03775_),
    .X(_00507_));
 sky130_fd_sc_hd__mux2_1 _07791_ (.A0(net1037),
    .A1(\tms1x00.ins_pla_ors[6][6] ),
    .S(net293),
    .X(_03776_));
 sky130_fd_sc_hd__or2_1 _07792_ (.A(net550),
    .B(_03776_),
    .X(_00508_));
 sky130_fd_sc_hd__mux2_1 _07793_ (.A0(net1013),
    .A1(\tms1x00.ins_pla_ors[6][9] ),
    .S(net294),
    .X(_03777_));
 sky130_fd_sc_hd__or2_1 _07794_ (.A(net552),
    .B(_03777_),
    .X(_00509_));
 sky130_fd_sc_hd__mux2_1 _07795_ (.A0(net974),
    .A1(\tms1x00.ins_pla_ors[6][10] ),
    .S(net294),
    .X(_03778_));
 sky130_fd_sc_hd__or2_1 _07796_ (.A(net552),
    .B(_03778_),
    .X(_00510_));
 sky130_fd_sc_hd__mux2_1 _07797_ (.A0(net971),
    .A1(\tms1x00.ins_pla_ors[6][11] ),
    .S(net293),
    .X(_03779_));
 sky130_fd_sc_hd__or2_1 _07798_ (.A(net549),
    .B(_03779_),
    .X(_00511_));
 sky130_fd_sc_hd__mux2_1 _07799_ (.A0(net961),
    .A1(\tms1x00.ins_pla_ors[6][13] ),
    .S(net295),
    .X(_03780_));
 sky130_fd_sc_hd__or2_1 _07800_ (.A(net553),
    .B(_03780_),
    .X(_00512_));
 sky130_fd_sc_hd__mux2_1 _07801_ (.A0(net955),
    .A1(\tms1x00.ins_pla_ors[6][14] ),
    .S(net295),
    .X(_03781_));
 sky130_fd_sc_hd__or2_1 _07802_ (.A(net547),
    .B(_03781_),
    .X(_00513_));
 sky130_fd_sc_hd__mux2_1 _07803_ (.A0(net950),
    .A1(\tms1x00.ins_pla_ors[6][15] ),
    .S(net293),
    .X(_03782_));
 sky130_fd_sc_hd__or2_1 _07804_ (.A(net547),
    .B(_03782_),
    .X(_00514_));
 sky130_fd_sc_hd__mux2_1 _07805_ (.A0(net940),
    .A1(\tms1x00.ins_pla_ors[6][17] ),
    .S(net293),
    .X(_03783_));
 sky130_fd_sc_hd__or2_1 _07806_ (.A(net547),
    .B(_03783_),
    .X(_00515_));
 sky130_fd_sc_hd__mux2_1 _07807_ (.A0(net935),
    .A1(\tms1x00.ins_pla_ors[6][19] ),
    .S(net293),
    .X(_03784_));
 sky130_fd_sc_hd__or2_1 _07808_ (.A(net546),
    .B(_03784_),
    .X(_00516_));
 sky130_fd_sc_hd__mux2_1 _07809_ (.A0(net1079),
    .A1(\tms1x00.ins_pla_ors[6][20] ),
    .S(net293),
    .X(_03785_));
 sky130_fd_sc_hd__or2_1 _07810_ (.A(net546),
    .B(_03785_),
    .X(_00517_));
 sky130_fd_sc_hd__mux2_1 _07811_ (.A0(net101),
    .A1(\tms1x00.ins_pla_ors[6][21] ),
    .S(net295),
    .X(_03786_));
 sky130_fd_sc_hd__or2_1 _07812_ (.A(net548),
    .B(_03786_),
    .X(_00518_));
 sky130_fd_sc_hd__mux2_1 _07813_ (.A0(net1076),
    .A1(\tms1x00.ins_pla_ors[6][22] ),
    .S(net293),
    .X(_03787_));
 sky130_fd_sc_hd__or2_1 _07814_ (.A(net544),
    .B(_03787_),
    .X(_00519_));
 sky130_fd_sc_hd__mux2_1 _07815_ (.A0(net103),
    .A1(\tms1x00.ins_pla_ors[6][23] ),
    .S(net294),
    .X(_03788_));
 sky130_fd_sc_hd__or2_1 _07816_ (.A(net551),
    .B(_03788_),
    .X(_00520_));
 sky130_fd_sc_hd__mux2_1 _07817_ (.A0(net1073),
    .A1(\tms1x00.ins_pla_ors[6][24] ),
    .S(net294),
    .X(_03789_));
 sky130_fd_sc_hd__or2_1 _07818_ (.A(net553),
    .B(_03789_),
    .X(_00521_));
 sky130_fd_sc_hd__nor2_8 _07819_ (.A(net717),
    .B(net355),
    .Y(_03790_));
 sky130_fd_sc_hd__nor2_1 _07820_ (.A(net519),
    .B(net291),
    .Y(_03791_));
 sky130_fd_sc_hd__inv_2 _07821_ (.A(net212),
    .Y(_03792_));
 sky130_fd_sc_hd__a22o_1 _07822_ (.A1(net979),
    .A2(net292),
    .B1(net213),
    .B2(\tms1x00.ins_pla_ors[10][0] ),
    .X(_00522_));
 sky130_fd_sc_hd__a22o_1 _07823_ (.A1(net1066),
    .A2(net292),
    .B1(net212),
    .B2(\tms1x00.ins_pla_ors[10][2] ),
    .X(_00523_));
 sky130_fd_sc_hd__a22o_1 _07824_ (.A1(net1049),
    .A2(net291),
    .B1(net212),
    .B2(\tms1x00.ins_pla_ors[10][4] ),
    .X(_00524_));
 sky130_fd_sc_hd__a22o_1 _07825_ (.A1(net1037),
    .A2(net292),
    .B1(net214),
    .B2(\tms1x00.ins_pla_ors[10][6] ),
    .X(_00525_));
 sky130_fd_sc_hd__a22o_1 _07826_ (.A1(net1022),
    .A2(net291),
    .B1(net213),
    .B2(\tms1x00.ins_pla_ors[10][8] ),
    .X(_00526_));
 sky130_fd_sc_hd__o32a_1 _07827_ (.A1(net1010),
    .A2(net718),
    .A3(net356),
    .B1(_03792_),
    .B2(\tms1x00.ins_pla_ors[10][9] ),
    .X(_00527_));
 sky130_fd_sc_hd__a22o_1 _07828_ (.A1(net972),
    .A2(net292),
    .B1(net212),
    .B2(\tms1x00.ins_pla_ors[10][10] ),
    .X(_00528_));
 sky130_fd_sc_hd__a22o_1 _07829_ (.A1(net968),
    .A2(net291),
    .B1(net213),
    .B2(\tms1x00.ins_pla_ors[10][11] ),
    .X(_00529_));
 sky130_fd_sc_hd__a22o_1 _07830_ (.A1(net965),
    .A2(net291),
    .B1(net212),
    .B2(\tms1x00.ins_pla_ors[10][12] ),
    .X(_00530_));
 sky130_fd_sc_hd__a22o_1 _07831_ (.A1(net960),
    .A2(net291),
    .B1(net212),
    .B2(\tms1x00.ins_pla_ors[10][13] ),
    .X(_00531_));
 sky130_fd_sc_hd__a22o_1 _07832_ (.A1(net953),
    .A2(net291),
    .B1(net212),
    .B2(\tms1x00.ins_pla_ors[10][14] ),
    .X(_00532_));
 sky130_fd_sc_hd__a22o_1 _07833_ (.A1(net948),
    .A2(net291),
    .B1(net212),
    .B2(\tms1x00.ins_pla_ors[10][15] ),
    .X(_00533_));
 sky130_fd_sc_hd__a22o_1 _07834_ (.A1(net942),
    .A2(net292),
    .B1(net215),
    .B2(\tms1x00.ins_pla_ors[10][16] ),
    .X(_00534_));
 sky130_fd_sc_hd__a22o_1 _07835_ (.A1(net938),
    .A2(net292),
    .B1(net215),
    .B2(\tms1x00.ins_pla_ors[10][18] ),
    .X(_00535_));
 sky130_fd_sc_hd__a22o_1 _07836_ (.A1(net1078),
    .A2(net292),
    .B1(net214),
    .B2(\tms1x00.ins_pla_ors[10][20] ),
    .X(_00536_));
 sky130_fd_sc_hd__a22o_1 _07837_ (.A1(net1077),
    .A2(net291),
    .B1(net212),
    .B2(\tms1x00.ins_pla_ors[10][21] ),
    .X(_00537_));
 sky130_fd_sc_hd__a22o_1 _07838_ (.A1(net1075),
    .A2(net292),
    .B1(net214),
    .B2(\tms1x00.ins_pla_ors[10][22] ),
    .X(_00538_));
 sky130_fd_sc_hd__a22o_1 _07839_ (.A1(net1074),
    .A2(net292),
    .B1(net214),
    .B2(\tms1x00.ins_pla_ors[10][23] ),
    .X(_00539_));
 sky130_fd_sc_hd__a22o_1 _07840_ (.A1(net105),
    .A2(_03790_),
    .B1(net214),
    .B2(\tms1x00.ins_pla_ors[10][25] ),
    .X(_00540_));
 sky130_fd_sc_hd__a22o_1 _07841_ (.A1(net107),
    .A2(_03790_),
    .B1(net214),
    .B2(\tms1x00.ins_pla_ors[10][27] ),
    .X(_00541_));
 sky130_fd_sc_hd__a22o_1 _07842_ (.A1(net109),
    .A2(_03790_),
    .B1(net215),
    .B2(\tms1x00.ins_pla_ors[10][29] ),
    .X(_00542_));
 sky130_fd_sc_hd__mux2_1 _07843_ (.A0(net353),
    .A1(\tms1x00.ins_pla_ands[29][8] ),
    .S(net220),
    .X(_00543_));
 sky130_fd_sc_hd__mux2_1 _07844_ (.A0(_03579_),
    .A1(\tms1x00.ins_pla_ands[29][10] ),
    .S(net220),
    .X(_00544_));
 sky130_fd_sc_hd__mux2_1 _07845_ (.A0(_03487_),
    .A1(\tms1x00.ins_pla_ands[29][13] ),
    .S(net220),
    .X(_00545_));
 sky130_fd_sc_hd__mux2_1 _07846_ (.A0(_03537_),
    .A1(\tms1x00.ins_pla_ands[29][14] ),
    .S(net220),
    .X(_00546_));
 sky130_fd_sc_hd__and3_4 _07847_ (.A(net766),
    .B(net350),
    .C(_03471_),
    .X(_03793_));
 sky130_fd_sc_hd__nor2_8 _07848_ (.A(net511),
    .B(net290),
    .Y(_03794_));
 sky130_fd_sc_hd__mux2_1 _07849_ (.A0(net343),
    .A1(\tms1x00.ins_pla_ands[25][0] ),
    .S(_03794_),
    .X(_00547_));
 sky130_fd_sc_hd__mux2_1 _07850_ (.A0(net344),
    .A1(\tms1x00.ins_pla_ands[25][1] ),
    .S(_03794_),
    .X(_00548_));
 sky130_fd_sc_hd__mux2_1 _07851_ (.A0(_03482_),
    .A1(\tms1x00.ins_pla_ands[25][10] ),
    .S(_03794_),
    .X(_00549_));
 sky130_fd_sc_hd__mux2_1 _07852_ (.A0(net347),
    .A1(\tms1x00.ins_pla_ands[25][11] ),
    .S(_03794_),
    .X(_00550_));
 sky130_fd_sc_hd__nor2_1 _07853_ (.A(net840),
    .B(net345),
    .Y(_03795_));
 sky130_fd_sc_hd__or2_1 _07854_ (.A(net839),
    .B(net346),
    .X(_03796_));
 sky130_fd_sc_hd__or2_1 _07855_ (.A(\tms1x00.ins_pla_ors[0][0] ),
    .B(net289),
    .X(_03797_));
 sky130_fd_sc_hd__o211a_1 _07856_ (.A1(net982),
    .A2(net285),
    .B1(_03797_),
    .C1(net486),
    .X(_00551_));
 sky130_fd_sc_hd__or2_1 _07857_ (.A(\tms1x00.ins_pla_ors[0][1] ),
    .B(net288),
    .X(_03798_));
 sky130_fd_sc_hd__o211a_1 _07858_ (.A1(net934),
    .A2(net284),
    .B1(_03798_),
    .C1(net485),
    .X(_00552_));
 sky130_fd_sc_hd__or2_1 _07859_ (.A(\tms1x00.ins_pla_ors[0][2] ),
    .B(net288),
    .X(_03799_));
 sky130_fd_sc_hd__o211a_1 _07860_ (.A1(net1070),
    .A2(net284),
    .B1(_03799_),
    .C1(net485),
    .X(_00553_));
 sky130_fd_sc_hd__or2_1 _07861_ (.A(\tms1x00.ins_pla_ors[0][3] ),
    .B(net288),
    .X(_03800_));
 sky130_fd_sc_hd__o211a_1 _07862_ (.A1(net1060),
    .A2(net284),
    .B1(_03800_),
    .C1(net488),
    .X(_00554_));
 sky130_fd_sc_hd__or2_1 _07863_ (.A(\tms1x00.ins_pla_ors[0][4] ),
    .B(net288),
    .X(_03801_));
 sky130_fd_sc_hd__o211a_1 _07864_ (.A1(net1053),
    .A2(net284),
    .B1(_03801_),
    .C1(net488),
    .X(_00555_));
 sky130_fd_sc_hd__or2_1 _07865_ (.A(\tms1x00.ins_pla_ors[0][7] ),
    .B(net288),
    .X(_03802_));
 sky130_fd_sc_hd__o211a_1 _07866_ (.A1(net1029),
    .A2(net284),
    .B1(_03802_),
    .C1(net488),
    .X(_00556_));
 sky130_fd_sc_hd__or2_1 _07867_ (.A(\tms1x00.ins_pla_ors[0][8] ),
    .B(net288),
    .X(_03803_));
 sky130_fd_sc_hd__o211a_1 _07868_ (.A1(net1022),
    .A2(net284),
    .B1(_03803_),
    .C1(net485),
    .X(_00557_));
 sky130_fd_sc_hd__or2_1 _07869_ (.A(\tms1x00.ins_pla_ors[0][9] ),
    .B(net288),
    .X(_03804_));
 sky130_fd_sc_hd__o211a_1 _07870_ (.A1(net1013),
    .A2(net285),
    .B1(_03804_),
    .C1(net486),
    .X(_00558_));
 sky130_fd_sc_hd__mux2_1 _07871_ (.A0(net970),
    .A1(\tms1x00.ins_pla_ors[0][11] ),
    .S(net284),
    .X(_03805_));
 sky130_fd_sc_hd__or2_1 _07872_ (.A(net567),
    .B(_03805_),
    .X(_00559_));
 sky130_fd_sc_hd__or2_1 _07873_ (.A(\tms1x00.ins_pla_ors[0][13] ),
    .B(net289),
    .X(_03806_));
 sky130_fd_sc_hd__o211a_1 _07874_ (.A1(net961),
    .A2(net285),
    .B1(_03806_),
    .C1(net486),
    .X(_00560_));
 sky130_fd_sc_hd__or2_1 _07875_ (.A(\tms1x00.ins_pla_ors[0][14] ),
    .B(net289),
    .X(_03807_));
 sky130_fd_sc_hd__o211a_1 _07876_ (.A1(net955),
    .A2(net286),
    .B1(_03807_),
    .C1(net483),
    .X(_00561_));
 sky130_fd_sc_hd__or2_1 _07877_ (.A(\tms1x00.ins_pla_ors[0][15] ),
    .B(net289),
    .X(_03808_));
 sky130_fd_sc_hd__o211a_1 _07878_ (.A1(net950),
    .A2(net284),
    .B1(_03808_),
    .C1(net487),
    .X(_00562_));
 sky130_fd_sc_hd__or2_1 _07879_ (.A(\tms1x00.ins_pla_ors[0][16] ),
    .B(net289),
    .X(_03809_));
 sky130_fd_sc_hd__o211a_1 _07880_ (.A1(net942),
    .A2(net286),
    .B1(_03809_),
    .C1(net483),
    .X(_00563_));
 sky130_fd_sc_hd__or2_1 _07881_ (.A(\tms1x00.ins_pla_ors[0][17] ),
    .B(net289),
    .X(_03810_));
 sky130_fd_sc_hd__o211a_1 _07882_ (.A1(net940),
    .A2(net283),
    .B1(_03810_),
    .C1(net489),
    .X(_00564_));
 sky130_fd_sc_hd__or2_1 _07883_ (.A(\tms1x00.ins_pla_ors[0][18] ),
    .B(net288),
    .X(_03811_));
 sky130_fd_sc_hd__o211a_1 _07884_ (.A1(net939),
    .A2(net285),
    .B1(_03811_),
    .C1(net487),
    .X(_00565_));
 sky130_fd_sc_hd__or2_1 _07885_ (.A(\tms1x00.ins_pla_ors[0][19] ),
    .B(net287),
    .X(_03812_));
 sky130_fd_sc_hd__o211a_1 _07886_ (.A1(net935),
    .A2(net283),
    .B1(_03812_),
    .C1(net483),
    .X(_00566_));
 sky130_fd_sc_hd__or2_1 _07887_ (.A(\tms1x00.ins_pla_ors[0][20] ),
    .B(net287),
    .X(_03813_));
 sky130_fd_sc_hd__o211a_1 _07888_ (.A1(net1079),
    .A2(net286),
    .B1(_03813_),
    .C1(net483),
    .X(_00567_));
 sky130_fd_sc_hd__or2_1 _07889_ (.A(\tms1x00.ins_pla_ors[0][21] ),
    .B(net287),
    .X(_03814_));
 sky130_fd_sc_hd__o211a_1 _07890_ (.A1(net101),
    .A2(net286),
    .B1(_03814_),
    .C1(net484),
    .X(_00568_));
 sky130_fd_sc_hd__or2_1 _07891_ (.A(\tms1x00.ins_pla_ors[0][22] ),
    .B(net287),
    .X(_03815_));
 sky130_fd_sc_hd__o211a_1 _07892_ (.A1(net1076),
    .A2(net283),
    .B1(_03815_),
    .C1(net482),
    .X(_00569_));
 sky130_fd_sc_hd__or2_1 _07893_ (.A(\tms1x00.ins_pla_ors[0][24] ),
    .B(net289),
    .X(_03816_));
 sky130_fd_sc_hd__o211a_1 _07894_ (.A1(net1073),
    .A2(net285),
    .B1(_03816_),
    .C1(net486),
    .X(_00570_));
 sky130_fd_sc_hd__or2_1 _07895_ (.A(\tms1x00.ins_pla_ors[0][26] ),
    .B(net287),
    .X(_03817_));
 sky130_fd_sc_hd__o211a_1 _07896_ (.A1(net106),
    .A2(net283),
    .B1(_03817_),
    .C1(net482),
    .X(_00571_));
 sky130_fd_sc_hd__or2_1 _07897_ (.A(\tms1x00.ins_pla_ors[0][27] ),
    .B(net287),
    .X(_03818_));
 sky130_fd_sc_hd__o211a_1 _07898_ (.A1(net107),
    .A2(net283),
    .B1(_03818_),
    .C1(net482),
    .X(_00572_));
 sky130_fd_sc_hd__or2_1 _07899_ (.A(\tms1x00.ins_pla_ors[0][28] ),
    .B(net287),
    .X(_03819_));
 sky130_fd_sc_hd__o211a_1 _07900_ (.A1(net108),
    .A2(net283),
    .B1(_03819_),
    .C1(net482),
    .X(_00573_));
 sky130_fd_sc_hd__or2_1 _07901_ (.A(\tms1x00.ins_pla_ors[0][29] ),
    .B(net287),
    .X(_03820_));
 sky130_fd_sc_hd__o211a_1 _07902_ (.A1(net109),
    .A2(net283),
    .B1(_03820_),
    .C1(net482),
    .X(_00574_));
 sky130_fd_sc_hd__nor2_4 _07903_ (.A(net889),
    .B(net345),
    .Y(_03821_));
 sky130_fd_sc_hd__or2_1 _07904_ (.A(net889),
    .B(net345),
    .X(_03822_));
 sky130_fd_sc_hd__mux2_1 _07905_ (.A0(net1070),
    .A1(\tms1x00.ins_pla_ors[5][2] ),
    .S(net281),
    .X(_03823_));
 sky130_fd_sc_hd__or2_1 _07906_ (.A(net549),
    .B(_03823_),
    .X(_00575_));
 sky130_fd_sc_hd__mux2_1 _07907_ (.A0(net1044),
    .A1(\tms1x00.ins_pla_ors[5][5] ),
    .S(net280),
    .X(_03824_));
 sky130_fd_sc_hd__or2_1 _07908_ (.A(net542),
    .B(_03824_),
    .X(_00576_));
 sky130_fd_sc_hd__mux2_1 _07909_ (.A0(net1037),
    .A1(\tms1x00.ins_pla_ors[5][6] ),
    .S(net282),
    .X(_03825_));
 sky130_fd_sc_hd__or2_1 _07910_ (.A(net541),
    .B(_03825_),
    .X(_00577_));
 sky130_fd_sc_hd__mux2_1 _07911_ (.A0(net1013),
    .A1(\tms1x00.ins_pla_ors[5][9] ),
    .S(net282),
    .X(_03826_));
 sky130_fd_sc_hd__or2_1 _07912_ (.A(net550),
    .B(_03826_),
    .X(_00578_));
 sky130_fd_sc_hd__mux2_1 _07913_ (.A0(net975),
    .A1(\tms1x00.ins_pla_ors[5][10] ),
    .S(net280),
    .X(_03827_));
 sky130_fd_sc_hd__or2_1 _07914_ (.A(net541),
    .B(_03827_),
    .X(_00579_));
 sky130_fd_sc_hd__mux2_1 _07915_ (.A0(net971),
    .A1(\tms1x00.ins_pla_ors[5][11] ),
    .S(net281),
    .X(_03828_));
 sky130_fd_sc_hd__or2_1 _07916_ (.A(net549),
    .B(_03828_),
    .X(_00580_));
 sky130_fd_sc_hd__mux2_1 _07917_ (.A0(net966),
    .A1(\tms1x00.ins_pla_ors[5][12] ),
    .S(net281),
    .X(_03829_));
 sky130_fd_sc_hd__or2_1 _07918_ (.A(net545),
    .B(_03829_),
    .X(_00581_));
 sky130_fd_sc_hd__mux2_1 _07919_ (.A0(net962),
    .A1(\tms1x00.ins_pla_ors[5][13] ),
    .S(net280),
    .X(_03830_));
 sky130_fd_sc_hd__or2_1 _07920_ (.A(net542),
    .B(_03830_),
    .X(_00582_));
 sky130_fd_sc_hd__mux2_1 _07921_ (.A0(net955),
    .A1(\tms1x00.ins_pla_ors[5][14] ),
    .S(net281),
    .X(_03831_));
 sky130_fd_sc_hd__or2_1 _07922_ (.A(net547),
    .B(_03831_),
    .X(_00583_));
 sky130_fd_sc_hd__mux2_1 _07923_ (.A0(net950),
    .A1(\tms1x00.ins_pla_ors[5][15] ),
    .S(net281),
    .X(_03832_));
 sky130_fd_sc_hd__or2_1 _07924_ (.A(net544),
    .B(_03832_),
    .X(_00584_));
 sky130_fd_sc_hd__mux2_1 _07925_ (.A0(net940),
    .A1(\tms1x00.ins_pla_ors[5][17] ),
    .S(net281),
    .X(_03833_));
 sky130_fd_sc_hd__or2_1 _07926_ (.A(net550),
    .B(_03833_),
    .X(_00585_));
 sky130_fd_sc_hd__mux2_1 _07927_ (.A0(net938),
    .A1(\tms1x00.ins_pla_ors[5][18] ),
    .S(net280),
    .X(_03834_));
 sky130_fd_sc_hd__or2_1 _07928_ (.A(net541),
    .B(_03834_),
    .X(_00586_));
 sky130_fd_sc_hd__mux2_1 _07929_ (.A0(net935),
    .A1(\tms1x00.ins_pla_ors[5][19] ),
    .S(net281),
    .X(_03835_));
 sky130_fd_sc_hd__or2_1 _07930_ (.A(net546),
    .B(_03835_),
    .X(_00587_));
 sky130_fd_sc_hd__or2_1 _07931_ (.A(\tms1x00.ins_pla_ors[5][20] ),
    .B(_03821_),
    .X(_03836_));
 sky130_fd_sc_hd__o211a_1 _07932_ (.A1(net1079),
    .A2(net281),
    .B1(_03836_),
    .C1(net483),
    .X(_00588_));
 sky130_fd_sc_hd__mux2_1 _07933_ (.A0(net1076),
    .A1(\tms1x00.ins_pla_ors[5][22] ),
    .S(net280),
    .X(_03837_));
 sky130_fd_sc_hd__or2_1 _07934_ (.A(net544),
    .B(_03837_),
    .X(_00589_));
 sky130_fd_sc_hd__mux2_1 _07935_ (.A0(net103),
    .A1(\tms1x00.ins_pla_ors[5][23] ),
    .S(net282),
    .X(_03838_));
 sky130_fd_sc_hd__or2_1 _07936_ (.A(net551),
    .B(_03838_),
    .X(_00590_));
 sky130_fd_sc_hd__mux2_1 _07937_ (.A0(net105),
    .A1(\tms1x00.ins_pla_ors[5][25] ),
    .S(net280),
    .X(_03839_));
 sky130_fd_sc_hd__or2_1 _07938_ (.A(net539),
    .B(_03839_),
    .X(_00591_));
 sky130_fd_sc_hd__and3_4 _07939_ (.A(net874),
    .B(net352),
    .C(net708),
    .X(_03840_));
 sky130_fd_sc_hd__or3_4 _07940_ (.A(net868),
    .B(_03470_),
    .C(net706),
    .X(_03841_));
 sky130_fd_sc_hd__nor2_2 _07941_ (.A(net377),
    .B(_03840_),
    .Y(_03842_));
 sky130_fd_sc_hd__nand2_1 _07942_ (.A(net370),
    .B(_03841_),
    .Y(_03843_));
 sky130_fd_sc_hd__nor2_1 _07943_ (.A(net392),
    .B(_03840_),
    .Y(_03844_));
 sky130_fd_sc_hd__nand2_2 _07944_ (.A(net384),
    .B(_03841_),
    .Y(_03845_));
 sky130_fd_sc_hd__a22o_1 _07945_ (.A1(\tms1x00.ins_pla_ands[3][1] ),
    .A2(_03842_),
    .B1(_03845_),
    .B2(net354),
    .X(_00592_));
 sky130_fd_sc_hd__a22o_1 _07946_ (.A1(\tms1x00.ins_pla_ands[3][3] ),
    .A2(_03842_),
    .B1(_03845_),
    .B2(_03534_),
    .X(_00593_));
 sky130_fd_sc_hd__a22o_1 _07947_ (.A1(\tms1x00.ins_pla_ands[3][5] ),
    .A2(_03842_),
    .B1(_03845_),
    .B2(_03712_),
    .X(_00594_));
 sky130_fd_sc_hd__a22o_1 _07948_ (.A1(\tms1x00.ins_pla_ands[3][6] ),
    .A2(_03842_),
    .B1(_03845_),
    .B2(_03435_),
    .X(_00595_));
 sky130_fd_sc_hd__a22o_1 _07949_ (.A1(\tms1x00.ins_pla_ands[3][8] ),
    .A2(_03842_),
    .B1(_03845_),
    .B2(net353),
    .X(_00596_));
 sky130_fd_sc_hd__o22a_1 _07950_ (.A1(\tms1x00.ins_pla_ands[3][9] ),
    .A2(_03843_),
    .B1(_03844_),
    .B2(_03578_),
    .X(_00597_));
 sky130_fd_sc_hd__a22o_1 _07951_ (.A1(\tms1x00.ins_pla_ands[3][12] ),
    .A2(_03842_),
    .B1(_03845_),
    .B2(_03588_),
    .X(_00598_));
 sky130_fd_sc_hd__o22a_1 _07952_ (.A1(\tms1x00.ins_pla_ands[3][13] ),
    .A2(_03843_),
    .B1(_03844_),
    .B2(_03589_),
    .X(_00599_));
 sky130_fd_sc_hd__mux2_1 _07953_ (.A0(net354),
    .A1(\tms1x00.ins_pla_ors[10][1] ),
    .S(net213),
    .X(_00600_));
 sky130_fd_sc_hd__mux2_1 _07954_ (.A0(_03433_),
    .A1(\tms1x00.ins_pla_ors[10][3] ),
    .S(net214),
    .X(_00601_));
 sky130_fd_sc_hd__mux2_1 _07955_ (.A0(_03577_),
    .A1(\tms1x00.ins_pla_ors[10][5] ),
    .S(net213),
    .X(_00602_));
 sky130_fd_sc_hd__mux2_1 _07956_ (.A0(_03437_),
    .A1(\tms1x00.ins_pla_ors[10][7] ),
    .S(net213),
    .X(_00603_));
 sky130_fd_sc_hd__mux2_1 _07957_ (.A0(_03443_),
    .A1(\tms1x00.ins_pla_ors[10][17] ),
    .S(net214),
    .X(_00604_));
 sky130_fd_sc_hd__a221o_1 _07958_ (.A1(net937),
    .A2(net291),
    .B1(net212),
    .B2(\tms1x00.ins_pla_ors[10][19] ),
    .C1(net389),
    .X(_00605_));
 sky130_fd_sc_hd__mux2_1 _07959_ (.A0(_03520_),
    .A1(\tms1x00.ins_pla_ors[10][24] ),
    .S(net215),
    .X(_00606_));
 sky130_fd_sc_hd__mux2_1 _07960_ (.A0(_03448_),
    .A1(\tms1x00.ins_pla_ors[10][26] ),
    .S(net214),
    .X(_00607_));
 sky130_fd_sc_hd__mux2_1 _07961_ (.A0(_03450_),
    .A1(\tms1x00.ins_pla_ors[10][28] ),
    .S(net214),
    .X(_00608_));
 sky130_fd_sc_hd__a31o_1 _07962_ (.A1(\tms1x00.ins_pla_ors[0][5] ),
    .A2(net372),
    .A3(net284),
    .B1(net394),
    .X(_03846_));
 sky130_fd_sc_hd__a21o_1 _07963_ (.A1(_03457_),
    .A2(net288),
    .B1(_03846_),
    .X(_00609_));
 sky130_fd_sc_hd__a31o_1 _07964_ (.A1(\tms1x00.ins_pla_ors[0][6] ),
    .A2(net373),
    .A3(net284),
    .B1(net396),
    .X(_03847_));
 sky130_fd_sc_hd__a21o_1 _07965_ (.A1(_03434_),
    .A2(net288),
    .B1(_03847_),
    .X(_00610_));
 sky130_fd_sc_hd__mux2_1 _07966_ (.A0(net975),
    .A1(\tms1x00.ins_pla_ors[0][10] ),
    .S(net283),
    .X(_03848_));
 sky130_fd_sc_hd__o21a_1 _07967_ (.A1(net379),
    .A2(_03848_),
    .B1(net387),
    .X(_00611_));
 sky130_fd_sc_hd__a21o_1 _07968_ (.A1(net386),
    .A2(net283),
    .B1(_03485_),
    .X(_03849_));
 sky130_fd_sc_hd__o31a_1 _07969_ (.A1(\tms1x00.ins_pla_ors[0][12] ),
    .A2(net379),
    .A3(net287),
    .B1(_03849_),
    .X(_00612_));
 sky130_fd_sc_hd__mux2_1 _07970_ (.A0(net103),
    .A1(\tms1x00.ins_pla_ors[0][23] ),
    .S(net285),
    .X(_03850_));
 sky130_fd_sc_hd__o21a_1 _07971_ (.A1(net379),
    .A2(_03850_),
    .B1(net387),
    .X(_00613_));
 sky130_fd_sc_hd__a31o_1 _07972_ (.A1(\tms1x00.ins_pla_ors[0][25] ),
    .A2(net372),
    .A3(net283),
    .B1(net395),
    .X(_03851_));
 sky130_fd_sc_hd__a21o_1 _07973_ (.A1(_03498_),
    .A2(net287),
    .B1(_03851_),
    .X(_00614_));
 sky130_fd_sc_hd__o22a_1 _07974_ (.A1(\tms1x00.ins_pla_ands[23][2] ),
    .A2(net317),
    .B1(_03596_),
    .B2(_03428_),
    .X(_00615_));
 sky130_fd_sc_hd__mux2_1 _07975_ (.A0(\tms1x00.ins_pla_ands[23][3] ),
    .A1(net1058),
    .S(net317),
    .X(_03852_));
 sky130_fd_sc_hd__or2_1 _07976_ (.A(net524),
    .B(_03852_),
    .X(_00616_));
 sky130_fd_sc_hd__mux2_1 _07977_ (.A0(\tms1x00.ins_pla_ands[23][4] ),
    .A1(net1049),
    .S(_03595_),
    .X(_03853_));
 sky130_fd_sc_hd__or2_1 _07978_ (.A(net524),
    .B(_03853_),
    .X(_00617_));
 sky130_fd_sc_hd__o22a_1 _07979_ (.A1(\tms1x00.ins_pla_ands[23][5] ),
    .A2(_03595_),
    .B1(_03596_),
    .B2(net366),
    .X(_00618_));
 sky130_fd_sc_hd__mux2_1 _07980_ (.A0(\tms1x00.ins_pla_ands[23][6] ),
    .A1(net1033),
    .S(net317),
    .X(_03854_));
 sky130_fd_sc_hd__or2_1 _07981_ (.A(net524),
    .B(_03854_),
    .X(_00619_));
 sky130_fd_sc_hd__o22a_1 _07982_ (.A1(\tms1x00.ins_pla_ands[23][7] ),
    .A2(_03595_),
    .B1(_03596_),
    .B2(net367),
    .X(_00620_));
 sky130_fd_sc_hd__mux2_1 _07983_ (.A0(\tms1x00.ins_pla_ands[23][8] ),
    .A1(net1014),
    .S(net317),
    .X(_03855_));
 sky130_fd_sc_hd__or2_1 _07984_ (.A(net514),
    .B(_03855_),
    .X(_00621_));
 sky130_fd_sc_hd__o22a_1 _07985_ (.A1(\tms1x00.ins_pla_ands[23][9] ),
    .A2(net317),
    .B1(_03596_),
    .B2(net364),
    .X(_00622_));
 sky130_fd_sc_hd__mux2_1 _07986_ (.A0(\tms1x00.ins_pla_ands[23][12] ),
    .A1(net963),
    .S(net317),
    .X(_03856_));
 sky130_fd_sc_hd__or2_1 _07987_ (.A(net514),
    .B(_03856_),
    .X(_00623_));
 sky130_fd_sc_hd__o22a_1 _07988_ (.A1(\tms1x00.ins_pla_ands[23][13] ),
    .A2(net317),
    .B1(_03596_),
    .B2(net363),
    .X(_00624_));
 sky130_fd_sc_hd__mux2_1 _07989_ (.A0(\tms1x00.ins_pla_ands[23][14] ),
    .A1(net951),
    .S(net317),
    .X(_03857_));
 sky130_fd_sc_hd__or2_1 _07990_ (.A(net513),
    .B(_03857_),
    .X(_00625_));
 sky130_fd_sc_hd__mux2_1 _07991_ (.A0(\tms1x00.ins_pla_ands[23][15] ),
    .A1(net944),
    .S(net317),
    .X(_03858_));
 sky130_fd_sc_hd__and2_1 _07992_ (.A(net459),
    .B(_03858_),
    .X(_00626_));
 sky130_fd_sc_hd__and3_4 _07993_ (.A(net628),
    .B(net351),
    .C(net596),
    .X(_03859_));
 sky130_fd_sc_hd__or3_4 _07994_ (.A(net608),
    .B(net349),
    .C(net594),
    .X(_03860_));
 sky130_fd_sc_hd__or2_1 _07995_ (.A(\tms1x00.ins_pla_ands[14][2] ),
    .B(_03859_),
    .X(_03861_));
 sky130_fd_sc_hd__o211a_1 _07996_ (.A1(net1066),
    .A2(net278),
    .B1(_03861_),
    .C1(net466),
    .X(_00627_));
 sky130_fd_sc_hd__mux2_1 _07997_ (.A0(net1055),
    .A1(\tms1x00.ins_pla_ands[14][3] ),
    .S(net278),
    .X(_03862_));
 sky130_fd_sc_hd__or2_1 _07998_ (.A(net528),
    .B(_03862_),
    .X(_00628_));
 sky130_fd_sc_hd__mux2_1 _07999_ (.A0(net1047),
    .A1(\tms1x00.ins_pla_ands[14][4] ),
    .S(net279),
    .X(_03863_));
 sky130_fd_sc_hd__or2_1 _08000_ (.A(net528),
    .B(_03863_),
    .X(_00629_));
 sky130_fd_sc_hd__or2_1 _08001_ (.A(\tms1x00.ins_pla_ands[14][5] ),
    .B(_03859_),
    .X(_03864_));
 sky130_fd_sc_hd__o211a_1 _08002_ (.A1(net1039),
    .A2(net279),
    .B1(_03864_),
    .C1(net466),
    .X(_00630_));
 sky130_fd_sc_hd__mux2_1 _08003_ (.A0(net1015),
    .A1(\tms1x00.ins_pla_ands[14][8] ),
    .S(net278),
    .X(_03865_));
 sky130_fd_sc_hd__or2_1 _08004_ (.A(net526),
    .B(_03865_),
    .X(_00631_));
 sky130_fd_sc_hd__or2_1 _08005_ (.A(\tms1x00.ins_pla_ands[14][9] ),
    .B(_03859_),
    .X(_03866_));
 sky130_fd_sc_hd__o211a_1 _08006_ (.A1(net1008),
    .A2(net278),
    .B1(_03866_),
    .C1(net464),
    .X(_00632_));
 sky130_fd_sc_hd__or2_1 _08007_ (.A(\tms1x00.ins_pla_ands[14][10] ),
    .B(_03859_),
    .X(_03867_));
 sky130_fd_sc_hd__o211a_1 _08008_ (.A1(net972),
    .A2(net279),
    .B1(_03867_),
    .C1(net466),
    .X(_00633_));
 sky130_fd_sc_hd__mux2_1 _08009_ (.A0(net968),
    .A1(\tms1x00.ins_pla_ands[14][11] ),
    .S(net278),
    .X(_03868_));
 sky130_fd_sc_hd__or2_1 _08010_ (.A(net528),
    .B(_03868_),
    .X(_00634_));
 sky130_fd_sc_hd__mux2_1 _08011_ (.A0(net963),
    .A1(\tms1x00.ins_pla_ands[14][12] ),
    .S(net278),
    .X(_03869_));
 sky130_fd_sc_hd__or2_1 _08012_ (.A(net527),
    .B(_03869_),
    .X(_00635_));
 sky130_fd_sc_hd__or2_1 _08013_ (.A(\tms1x00.ins_pla_ands[14][13] ),
    .B(_03859_),
    .X(_03870_));
 sky130_fd_sc_hd__o211a_1 _08014_ (.A1(net959),
    .A2(net278),
    .B1(_03870_),
    .C1(net463),
    .X(_00636_));
 sky130_fd_sc_hd__mux2_1 _08015_ (.A0(net951),
    .A1(\tms1x00.ins_pla_ands[14][14] ),
    .S(net279),
    .X(_03871_));
 sky130_fd_sc_hd__or2_1 _08016_ (.A(net528),
    .B(_03871_),
    .X(_00637_));
 sky130_fd_sc_hd__or2_1 _08017_ (.A(\tms1x00.ins_pla_ands[14][15] ),
    .B(_03859_),
    .X(_03872_));
 sky130_fd_sc_hd__o211a_1 _08018_ (.A1(net946),
    .A2(net278),
    .B1(_03872_),
    .C1(net463),
    .X(_00638_));
 sky130_fd_sc_hd__or2_1 _08019_ (.A(\tms1x00.ins_pla_ands[4][1] ),
    .B(_03708_),
    .X(_03873_));
 sky130_fd_sc_hd__o211a_1 _08020_ (.A1(net933),
    .A2(net301),
    .B1(_03873_),
    .C1(net490),
    .X(_00639_));
 sky130_fd_sc_hd__or2_1 _08021_ (.A(\tms1x00.ins_pla_ands[4][2] ),
    .B(_03708_),
    .X(_03874_));
 sky130_fd_sc_hd__o211a_1 _08022_ (.A1(net1067),
    .A2(net301),
    .B1(_03874_),
    .C1(net490),
    .X(_00640_));
 sky130_fd_sc_hd__or2_1 _08023_ (.A(\tms1x00.ins_pla_ands[4][4] ),
    .B(_03708_),
    .X(_03875_));
 sky130_fd_sc_hd__o211a_1 _08024_ (.A1(net1050),
    .A2(net301),
    .B1(_03875_),
    .C1(net492),
    .X(_00641_));
 sky130_fd_sc_hd__or2_1 _08025_ (.A(\tms1x00.ins_pla_ands[4][7] ),
    .B(_03708_),
    .X(_03876_));
 sky130_fd_sc_hd__o211a_1 _08026_ (.A1(net1028),
    .A2(net301),
    .B1(_03876_),
    .C1(net490),
    .X(_00642_));
 sky130_fd_sc_hd__mux2_1 _08027_ (.A0(net1019),
    .A1(\tms1x00.ins_pla_ands[4][8] ),
    .S(_03709_),
    .X(_03877_));
 sky130_fd_sc_hd__or2_1 _08028_ (.A(net557),
    .B(_03877_),
    .X(_00643_));
 sky130_fd_sc_hd__or2_1 _08029_ (.A(\tms1x00.ins_pla_ands[4][9] ),
    .B(_03708_),
    .X(_03878_));
 sky130_fd_sc_hd__o211a_1 _08030_ (.A1(net1012),
    .A2(_03709_),
    .B1(_03878_),
    .C1(net490),
    .X(_00644_));
 sky130_fd_sc_hd__mux2_1 _08031_ (.A0(net974),
    .A1(\tms1x00.ins_pla_ands[4][10] ),
    .S(net301),
    .X(_03879_));
 sky130_fd_sc_hd__or2_1 _08032_ (.A(net557),
    .B(_03879_),
    .X(_00645_));
 sky130_fd_sc_hd__or2_1 _08033_ (.A(\tms1x00.ins_pla_ands[4][11] ),
    .B(_03708_),
    .X(_03880_));
 sky130_fd_sc_hd__o211a_1 _08034_ (.A1(net970),
    .A2(net301),
    .B1(_03880_),
    .C1(net490),
    .X(_00646_));
 sky130_fd_sc_hd__mux2_1 _08035_ (.A0(net957),
    .A1(\tms1x00.ins_pla_ands[4][14] ),
    .S(net301),
    .X(_03881_));
 sky130_fd_sc_hd__or2_1 _08036_ (.A(net558),
    .B(_03881_),
    .X(_00647_));
 sky130_fd_sc_hd__or2_1 _08037_ (.A(\tms1x00.ins_pla_ands[4][15] ),
    .B(_03708_),
    .X(_03882_));
 sky130_fd_sc_hd__o211a_1 _08038_ (.A1(net949),
    .A2(net301),
    .B1(_03882_),
    .C1(net493),
    .X(_00648_));
 sky130_fd_sc_hd__mux2_1 _08039_ (.A0(\tms1x00.ins_pla_ands[22][6] ),
    .A1(net1033),
    .S(net316),
    .X(_03883_));
 sky130_fd_sc_hd__or2_1 _08040_ (.A(net524),
    .B(_03883_),
    .X(_00649_));
 sky130_fd_sc_hd__o22a_1 _08041_ (.A1(\tms1x00.ins_pla_ands[22][7] ),
    .A2(net316),
    .B1(_03598_),
    .B2(net368),
    .X(_00650_));
 sky130_fd_sc_hd__mux2_1 _08042_ (.A0(\tms1x00.ins_pla_ands[22][8] ),
    .A1(net1014),
    .S(net316),
    .X(_03884_));
 sky130_fd_sc_hd__or2_1 _08043_ (.A(net514),
    .B(_03884_),
    .X(_00651_));
 sky130_fd_sc_hd__o22a_1 _08044_ (.A1(\tms1x00.ins_pla_ands[22][9] ),
    .A2(net316),
    .B1(_03598_),
    .B2(net364),
    .X(_00652_));
 sky130_fd_sc_hd__o22a_1 _08045_ (.A1(\tms1x00.ins_pla_ands[22][10] ),
    .A2(_03597_),
    .B1(_03598_),
    .B2(_03459_),
    .X(_00653_));
 sky130_fd_sc_hd__mux2_1 _08046_ (.A0(\tms1x00.ins_pla_ands[22][12] ),
    .A1(net963),
    .S(net316),
    .X(_03885_));
 sky130_fd_sc_hd__or2_1 _08047_ (.A(net515),
    .B(_03885_),
    .X(_00654_));
 sky130_fd_sc_hd__o22a_1 _08048_ (.A1(\tms1x00.ins_pla_ands[22][13] ),
    .A2(net316),
    .B1(_03598_),
    .B2(net363),
    .X(_00655_));
 sky130_fd_sc_hd__mux2_1 _08049_ (.A0(\tms1x00.ins_pla_ands[22][14] ),
    .A1(net951),
    .S(net316),
    .X(_03886_));
 sky130_fd_sc_hd__or2_1 _08050_ (.A(net517),
    .B(_03886_),
    .X(_00656_));
 sky130_fd_sc_hd__mux2_1 _08051_ (.A0(\tms1x00.ins_pla_ands[22][15] ),
    .A1(net944),
    .S(net316),
    .X(_03887_));
 sky130_fd_sc_hd__and2_1 _08052_ (.A(net459),
    .B(_03887_),
    .X(_00657_));
 sky130_fd_sc_hd__and3_4 _08053_ (.A(net902),
    .B(net351),
    .C(net596),
    .X(_03888_));
 sky130_fd_sc_hd__or3_4 _08054_ (.A(net882),
    .B(net348),
    .C(net594),
    .X(_03889_));
 sky130_fd_sc_hd__mux2_1 _08055_ (.A0(net1015),
    .A1(\tms1x00.ins_pla_ands[13][8] ),
    .S(_03889_),
    .X(_03890_));
 sky130_fd_sc_hd__or2_1 _08056_ (.A(net527),
    .B(_03890_),
    .X(_00658_));
 sky130_fd_sc_hd__or2_1 _08057_ (.A(\tms1x00.ins_pla_ands[13][9] ),
    .B(_03888_),
    .X(_03891_));
 sky130_fd_sc_hd__o211a_1 _08058_ (.A1(net1008),
    .A2(_03889_),
    .B1(_03891_),
    .C1(net465),
    .X(_00659_));
 sky130_fd_sc_hd__or2_1 _08059_ (.A(\tms1x00.ins_pla_ands[13][10] ),
    .B(_03888_),
    .X(_03892_));
 sky130_fd_sc_hd__o211a_1 _08060_ (.A1(net972),
    .A2(_03889_),
    .B1(_03892_),
    .C1(net466),
    .X(_00660_));
 sky130_fd_sc_hd__mux2_1 _08061_ (.A0(net968),
    .A1(\tms1x00.ins_pla_ands[13][11] ),
    .S(_03889_),
    .X(_03893_));
 sky130_fd_sc_hd__or2_1 _08062_ (.A(net529),
    .B(_03893_),
    .X(_00661_));
 sky130_fd_sc_hd__mux2_1 _08063_ (.A0(net964),
    .A1(\tms1x00.ins_pla_ands[13][12] ),
    .S(_03889_),
    .X(_03894_));
 sky130_fd_sc_hd__or2_1 _08064_ (.A(net527),
    .B(_03894_),
    .X(_00662_));
 sky130_fd_sc_hd__or2_1 _08065_ (.A(\tms1x00.ins_pla_ands[13][13] ),
    .B(_03888_),
    .X(_03895_));
 sky130_fd_sc_hd__o211a_1 _08066_ (.A1(net959),
    .A2(_03889_),
    .B1(_03895_),
    .C1(net464),
    .X(_00663_));
 sky130_fd_sc_hd__mux2_1 _08067_ (.A0(net952),
    .A1(\tms1x00.ins_pla_ands[13][14] ),
    .S(_03889_),
    .X(_03896_));
 sky130_fd_sc_hd__or2_1 _08068_ (.A(net528),
    .B(_03896_),
    .X(_00664_));
 sky130_fd_sc_hd__or2_1 _08069_ (.A(\tms1x00.ins_pla_ands[13][15] ),
    .B(_03888_),
    .X(_03897_));
 sky130_fd_sc_hd__o211a_1 _08070_ (.A1(net946),
    .A2(_03889_),
    .B1(_03897_),
    .C1(net464),
    .X(_00665_));
 sky130_fd_sc_hd__or2_1 _08071_ (.A(\tms1x00.ins_pla_ands[3][0] ),
    .B(_03840_),
    .X(_03898_));
 sky130_fd_sc_hd__o211a_1 _08072_ (.A1(net977),
    .A2(_03841_),
    .B1(_03898_),
    .C1(net470),
    .X(_00666_));
 sky130_fd_sc_hd__or2_1 _08073_ (.A(\tms1x00.ins_pla_ands[3][2] ),
    .B(_03840_),
    .X(_03899_));
 sky130_fd_sc_hd__o211a_1 _08074_ (.A1(net1070),
    .A2(_03841_),
    .B1(_03899_),
    .C1(net469),
    .X(_00667_));
 sky130_fd_sc_hd__or2_1 _08075_ (.A(\tms1x00.ins_pla_ands[3][4] ),
    .B(_03840_),
    .X(_03900_));
 sky130_fd_sc_hd__o211a_1 _08076_ (.A1(net1050),
    .A2(_03841_),
    .B1(_03900_),
    .C1(net469),
    .X(_00668_));
 sky130_fd_sc_hd__or2_1 _08077_ (.A(\tms1x00.ins_pla_ands[3][7] ),
    .B(_03840_),
    .X(_03901_));
 sky130_fd_sc_hd__o211a_1 _08078_ (.A1(net1025),
    .A2(_03841_),
    .B1(_03901_),
    .C1(net469),
    .X(_00669_));
 sky130_fd_sc_hd__mux2_1 _08079_ (.A0(net972),
    .A1(\tms1x00.ins_pla_ands[3][10] ),
    .S(_03841_),
    .X(_03902_));
 sky130_fd_sc_hd__or2_1 _08080_ (.A(net531),
    .B(_03902_),
    .X(_00670_));
 sky130_fd_sc_hd__or2_1 _08081_ (.A(\tms1x00.ins_pla_ands[3][11] ),
    .B(_03840_),
    .X(_03903_));
 sky130_fd_sc_hd__o211a_1 _08082_ (.A1(net968),
    .A2(_03841_),
    .B1(_03903_),
    .C1(net469),
    .X(_00671_));
 sky130_fd_sc_hd__mux2_1 _08083_ (.A0(net953),
    .A1(\tms1x00.ins_pla_ands[3][14] ),
    .S(_03841_),
    .X(_03904_));
 sky130_fd_sc_hd__or2_1 _08084_ (.A(net531),
    .B(_03904_),
    .X(_00672_));
 sky130_fd_sc_hd__or2_1 _08085_ (.A(\tms1x00.ins_pla_ands[3][15] ),
    .B(_03840_),
    .X(_03905_));
 sky130_fd_sc_hd__o211a_1 _08086_ (.A1(net949),
    .A2(_03841_),
    .B1(_03905_),
    .C1(net475),
    .X(_00673_));
 sky130_fd_sc_hd__or3_1 _08087_ (.A(\tms1x00.ins_pla_ands[14][0] ),
    .B(net376),
    .C(_03859_),
    .X(_03906_));
 sky130_fd_sc_hd__o211a_1 _08088_ (.A1(_03574_),
    .A2(net279),
    .B1(_03906_),
    .C1(net383),
    .X(_00674_));
 sky130_fd_sc_hd__a31o_1 _08089_ (.A1(\tms1x00.ins_pla_ands[14][1] ),
    .A2(net369),
    .A3(net278),
    .B1(net391),
    .X(_03907_));
 sky130_fd_sc_hd__a21o_1 _08090_ (.A1(net397),
    .A2(_03859_),
    .B1(_03907_),
    .X(_00675_));
 sky130_fd_sc_hd__or3_1 _08091_ (.A(\tms1x00.ins_pla_ands[14][6] ),
    .B(net376),
    .C(_03859_),
    .X(_03908_));
 sky130_fd_sc_hd__or2_4 _08092_ (.A(net1032),
    .B(net376),
    .X(_03909_));
 sky130_fd_sc_hd__o211a_1 _08093_ (.A1(net279),
    .A2(_03909_),
    .B1(_03908_),
    .C1(net383),
    .X(_00676_));
 sky130_fd_sc_hd__a31o_1 _08094_ (.A1(\tms1x00.ins_pla_ands[14][7] ),
    .A2(net369),
    .A3(net278),
    .B1(net391),
    .X(_03910_));
 sky130_fd_sc_hd__a21o_1 _08095_ (.A1(net368),
    .A2(_03859_),
    .B1(_03910_),
    .X(_00677_));
 sky130_fd_sc_hd__and3_4 _08096_ (.A(net741),
    .B(net351),
    .C(net596),
    .X(_03911_));
 sky130_fd_sc_hd__or3_2 _08097_ (.A(net723),
    .B(net348),
    .C(net594),
    .X(_03912_));
 sky130_fd_sc_hd__or3_1 _08098_ (.A(\tms1x00.ins_pla_ands[10][6] ),
    .B(net377),
    .C(_03911_),
    .X(_03913_));
 sky130_fd_sc_hd__o211a_1 _08099_ (.A1(_03909_),
    .A2(net277),
    .B1(_03913_),
    .C1(net383),
    .X(_00678_));
 sky130_fd_sc_hd__a31o_1 _08100_ (.A1(\tms1x00.ins_pla_ands[10][7] ),
    .A2(net369),
    .A3(net277),
    .B1(net391),
    .X(_03914_));
 sky130_fd_sc_hd__a21o_1 _08101_ (.A1(net368),
    .A2(_03911_),
    .B1(_03914_),
    .X(_00679_));
 sky130_fd_sc_hd__mux2_1 _08102_ (.A0(\tms1x00.ins_pla_ands[21][2] ),
    .A1(net1066),
    .S(net298),
    .X(_03915_));
 sky130_fd_sc_hd__or2_1 _08103_ (.A(net512),
    .B(_03915_),
    .X(_00680_));
 sky130_fd_sc_hd__o22a_1 _08104_ (.A1(\tms1x00.ins_pla_ands[21][3] ),
    .A2(net298),
    .B1(_03720_),
    .B2(_03430_),
    .X(_00681_));
 sky130_fd_sc_hd__o22a_1 _08105_ (.A1(\tms1x00.ins_pla_ands[21][4] ),
    .A2(net297),
    .B1(_03720_),
    .B2(_03478_),
    .X(_00682_));
 sky130_fd_sc_hd__mux2_1 _08106_ (.A0(\tms1x00.ins_pla_ands[21][5] ),
    .A1(net1041),
    .S(net297),
    .X(_03916_));
 sky130_fd_sc_hd__or2_1 _08107_ (.A(net512),
    .B(_03916_),
    .X(_00683_));
 sky130_fd_sc_hd__mux2_1 _08108_ (.A0(\tms1x00.ins_pla_ands[21][6] ),
    .A1(net1033),
    .S(net297),
    .X(_03917_));
 sky130_fd_sc_hd__or2_1 _08109_ (.A(net513),
    .B(_03917_),
    .X(_00684_));
 sky130_fd_sc_hd__o22a_1 _08110_ (.A1(\tms1x00.ins_pla_ands[21][7] ),
    .A2(net297),
    .B1(_03720_),
    .B2(net367),
    .X(_00685_));
 sky130_fd_sc_hd__mux2_1 _08111_ (.A0(\tms1x00.ins_pla_ands[21][8] ),
    .A1(net1014),
    .S(net297),
    .X(_03918_));
 sky130_fd_sc_hd__or2_1 _08112_ (.A(net513),
    .B(_03918_),
    .X(_00686_));
 sky130_fd_sc_hd__o22a_1 _08113_ (.A1(\tms1x00.ins_pla_ands[21][9] ),
    .A2(net297),
    .B1(_03720_),
    .B2(net364),
    .X(_00687_));
 sky130_fd_sc_hd__o22a_1 _08114_ (.A1(\tms1x00.ins_pla_ands[21][10] ),
    .A2(net298),
    .B1(_03720_),
    .B2(_03459_),
    .X(_00688_));
 sky130_fd_sc_hd__mux2_1 _08115_ (.A0(\tms1x00.ins_pla_ands[21][12] ),
    .A1(net963),
    .S(net297),
    .X(_03919_));
 sky130_fd_sc_hd__or2_1 _08116_ (.A(net513),
    .B(_03919_),
    .X(_00689_));
 sky130_fd_sc_hd__o22a_1 _08117_ (.A1(\tms1x00.ins_pla_ands[21][13] ),
    .A2(net297),
    .B1(_03720_),
    .B2(net363),
    .X(_00690_));
 sky130_fd_sc_hd__mux2_1 _08118_ (.A0(\tms1x00.ins_pla_ands[21][14] ),
    .A1(net951),
    .S(net297),
    .X(_03920_));
 sky130_fd_sc_hd__or2_1 _08119_ (.A(net513),
    .B(_03920_),
    .X(_00691_));
 sky130_fd_sc_hd__mux2_1 _08120_ (.A0(\tms1x00.ins_pla_ands[21][15] ),
    .A1(net944),
    .S(net297),
    .X(_03921_));
 sky130_fd_sc_hd__and2_1 _08121_ (.A(net459),
    .B(_03921_),
    .X(_00692_));
 sky130_fd_sc_hd__and3_4 _08122_ (.A(net820),
    .B(net351),
    .C(net596),
    .X(_03922_));
 sky130_fd_sc_hd__or3_1 _08123_ (.A(net801),
    .B(net348),
    .C(net594),
    .X(_03923_));
 sky130_fd_sc_hd__or2_1 _08124_ (.A(\tms1x00.ins_pla_ands[12][0] ),
    .B(_03922_),
    .X(_03924_));
 sky130_fd_sc_hd__o211a_1 _08125_ (.A1(net976),
    .A2(net274),
    .B1(_03924_),
    .C1(net463),
    .X(_00693_));
 sky130_fd_sc_hd__mux2_1 _08126_ (.A0(net1065),
    .A1(\tms1x00.ins_pla_ands[12][2] ),
    .S(net274),
    .X(_03925_));
 sky130_fd_sc_hd__or2_1 _08127_ (.A(net529),
    .B(_03925_),
    .X(_00694_));
 sky130_fd_sc_hd__or2_1 _08128_ (.A(\tms1x00.ins_pla_ands[12][3] ),
    .B(_03922_),
    .X(_03926_));
 sky130_fd_sc_hd__o211a_1 _08129_ (.A1(net1055),
    .A2(net274),
    .B1(_03926_),
    .C1(net463),
    .X(_00695_));
 sky130_fd_sc_hd__or2_1 _08130_ (.A(\tms1x00.ins_pla_ands[12][4] ),
    .B(_03922_),
    .X(_03927_));
 sky130_fd_sc_hd__o211a_1 _08131_ (.A1(net1047),
    .A2(net274),
    .B1(_03927_),
    .C1(net465),
    .X(_00696_));
 sky130_fd_sc_hd__mux2_1 _08132_ (.A0(net1039),
    .A1(\tms1x00.ins_pla_ands[12][5] ),
    .S(net275),
    .X(_03928_));
 sky130_fd_sc_hd__or2_1 _08133_ (.A(net527),
    .B(_03928_),
    .X(_00697_));
 sky130_fd_sc_hd__mux2_1 _08134_ (.A0(net1015),
    .A1(\tms1x00.ins_pla_ands[12][8] ),
    .S(net275),
    .X(_03929_));
 sky130_fd_sc_hd__or2_1 _08135_ (.A(net526),
    .B(_03929_),
    .X(_00698_));
 sky130_fd_sc_hd__or2_1 _08136_ (.A(\tms1x00.ins_pla_ands[12][9] ),
    .B(_03922_),
    .X(_03930_));
 sky130_fd_sc_hd__o211a_1 _08137_ (.A1(net1008),
    .A2(net274),
    .B1(_03930_),
    .C1(net463),
    .X(_00699_));
 sky130_fd_sc_hd__or2_1 _08138_ (.A(\tms1x00.ins_pla_ands[12][10] ),
    .B(_03922_),
    .X(_03931_));
 sky130_fd_sc_hd__o211a_1 _08139_ (.A1(net973),
    .A2(net274),
    .B1(_03931_),
    .C1(net463),
    .X(_00700_));
 sky130_fd_sc_hd__mux2_1 _08140_ (.A0(net969),
    .A1(\tms1x00.ins_pla_ands[12][11] ),
    .S(net274),
    .X(_03932_));
 sky130_fd_sc_hd__or2_1 _08141_ (.A(net527),
    .B(_03932_),
    .X(_00701_));
 sky130_fd_sc_hd__mux2_1 _08142_ (.A0(net964),
    .A1(\tms1x00.ins_pla_ands[12][12] ),
    .S(net275),
    .X(_03933_));
 sky130_fd_sc_hd__or2_1 _08143_ (.A(net527),
    .B(_03933_),
    .X(_00702_));
 sky130_fd_sc_hd__or2_1 _08144_ (.A(\tms1x00.ins_pla_ands[12][13] ),
    .B(_03922_),
    .X(_03934_));
 sky130_fd_sc_hd__o211a_1 _08145_ (.A1(net959),
    .A2(net274),
    .B1(_03934_),
    .C1(net463),
    .X(_00703_));
 sky130_fd_sc_hd__mux2_1 _08146_ (.A0(net952),
    .A1(\tms1x00.ins_pla_ands[12][14] ),
    .S(net275),
    .X(_03935_));
 sky130_fd_sc_hd__or2_1 _08147_ (.A(net526),
    .B(_03935_),
    .X(_00704_));
 sky130_fd_sc_hd__or2_1 _08148_ (.A(\tms1x00.ins_pla_ands[12][15] ),
    .B(_03922_),
    .X(_03936_));
 sky130_fd_sc_hd__o211a_1 _08149_ (.A1(net946),
    .A2(net274),
    .B1(_03936_),
    .C1(net465),
    .X(_00705_));
 sky130_fd_sc_hd__or2_1 _08150_ (.A(\tms1x00.ins_pla_ands[2][1] ),
    .B(_03581_),
    .X(_03937_));
 sky130_fd_sc_hd__o211a_1 _08151_ (.A1(net929),
    .A2(_03582_),
    .B1(_03937_),
    .C1(net469),
    .X(_00706_));
 sky130_fd_sc_hd__or2_1 _08152_ (.A(\tms1x00.ins_pla_ands[2][3] ),
    .B(_03581_),
    .X(_03938_));
 sky130_fd_sc_hd__o211a_1 _08153_ (.A1(net1059),
    .A2(_03582_),
    .B1(_03938_),
    .C1(net490),
    .X(_00707_));
 sky130_fd_sc_hd__or2_1 _08154_ (.A(\tms1x00.ins_pla_ands[2][5] ),
    .B(_03581_),
    .X(_03939_));
 sky130_fd_sc_hd__o211a_1 _08155_ (.A1(net1043),
    .A2(_03582_),
    .B1(_03939_),
    .C1(net493),
    .X(_00708_));
 sky130_fd_sc_hd__or2_1 _08156_ (.A(\tms1x00.ins_pla_ands[2][6] ),
    .B(_03581_),
    .X(_03940_));
 sky130_fd_sc_hd__o211a_1 _08157_ (.A1(net1036),
    .A2(_03582_),
    .B1(_03940_),
    .C1(net490),
    .X(_00709_));
 sky130_fd_sc_hd__mux2_1 _08158_ (.A0(net1019),
    .A1(\tms1x00.ins_pla_ands[2][8] ),
    .S(_03582_),
    .X(_03941_));
 sky130_fd_sc_hd__or2_1 _08159_ (.A(net535),
    .B(_03941_),
    .X(_00710_));
 sky130_fd_sc_hd__or2_1 _08160_ (.A(\tms1x00.ins_pla_ands[2][9] ),
    .B(_03581_),
    .X(_03942_));
 sky130_fd_sc_hd__o211a_1 _08161_ (.A1(net1009),
    .A2(_03582_),
    .B1(_03942_),
    .C1(net493),
    .X(_00711_));
 sky130_fd_sc_hd__mux2_1 _08162_ (.A0(net954),
    .A1(\tms1x00.ins_pla_ands[2][14] ),
    .S(_03582_),
    .X(_03943_));
 sky130_fd_sc_hd__or2_1 _08163_ (.A(net531),
    .B(_03943_),
    .X(_00712_));
 sky130_fd_sc_hd__or2_1 _08164_ (.A(\tms1x00.ins_pla_ands[2][15] ),
    .B(_03581_),
    .X(_03944_));
 sky130_fd_sc_hd__o211a_1 _08165_ (.A1(net949),
    .A2(_03582_),
    .B1(_03944_),
    .C1(net496),
    .X(_00713_));
 sky130_fd_sc_hd__or3_4 _08166_ (.A(net603),
    .B(net348),
    .C(net710),
    .X(_03945_));
 sky130_fd_sc_hd__mux2_1 _08167_ (.A0(net979),
    .A1(\tms1x00.ins_pla_ands[30][0] ),
    .S(net273),
    .X(_00714_));
 sky130_fd_sc_hd__mux2_1 _08168_ (.A0(net930),
    .A1(\tms1x00.ins_pla_ands[30][1] ),
    .S(net273),
    .X(_00715_));
 sky130_fd_sc_hd__mux2_1 _08169_ (.A0(net1066),
    .A1(\tms1x00.ins_pla_ands[30][2] ),
    .S(net273),
    .X(_00716_));
 sky130_fd_sc_hd__mux2_1 _08170_ (.A0(net1058),
    .A1(\tms1x00.ins_pla_ands[30][3] ),
    .S(net272),
    .X(_00717_));
 sky130_fd_sc_hd__mux2_1 _08171_ (.A0(net1049),
    .A1(\tms1x00.ins_pla_ands[30][4] ),
    .S(net272),
    .X(_00718_));
 sky130_fd_sc_hd__mux2_1 _08172_ (.A0(net1041),
    .A1(\tms1x00.ins_pla_ands[30][5] ),
    .S(net273),
    .X(_00719_));
 sky130_fd_sc_hd__mux2_1 _08173_ (.A0(net1033),
    .A1(\tms1x00.ins_pla_ands[30][6] ),
    .S(net272),
    .X(_00720_));
 sky130_fd_sc_hd__mux2_1 _08174_ (.A0(net1026),
    .A1(\tms1x00.ins_pla_ands[30][7] ),
    .S(net273),
    .X(_00721_));
 sky130_fd_sc_hd__mux2_1 _08175_ (.A0(net1014),
    .A1(\tms1x00.ins_pla_ands[30][8] ),
    .S(net272),
    .X(_00722_));
 sky130_fd_sc_hd__mux2_1 _08176_ (.A0(net1010),
    .A1(\tms1x00.ins_pla_ands[30][9] ),
    .S(net272),
    .X(_00723_));
 sky130_fd_sc_hd__mux2_1 _08177_ (.A0(net972),
    .A1(\tms1x00.ins_pla_ands[30][10] ),
    .S(net272),
    .X(_00724_));
 sky130_fd_sc_hd__mux2_1 _08178_ (.A0(net968),
    .A1(\tms1x00.ins_pla_ands[30][11] ),
    .S(net272),
    .X(_00725_));
 sky130_fd_sc_hd__mux2_1 _08179_ (.A0(net963),
    .A1(\tms1x00.ins_pla_ands[30][12] ),
    .S(net272),
    .X(_00726_));
 sky130_fd_sc_hd__mux2_1 _08180_ (.A0(net960),
    .A1(\tms1x00.ins_pla_ands[30][13] ),
    .S(net272),
    .X(_00727_));
 sky130_fd_sc_hd__mux2_1 _08181_ (.A0(net951),
    .A1(\tms1x00.ins_pla_ands[30][14] ),
    .S(net272),
    .X(_00728_));
 sky130_fd_sc_hd__mux2_1 _08182_ (.A0(net945),
    .A1(\tms1x00.ins_pla_ands[30][15] ),
    .S(net273),
    .X(_00729_));
 sky130_fd_sc_hd__o22a_1 _08183_ (.A1(\tms1x00.ins_pla_ands[20][4] ),
    .A2(_03721_),
    .B1(_03722_),
    .B2(_03478_),
    .X(_00730_));
 sky130_fd_sc_hd__mux2_1 _08184_ (.A0(\tms1x00.ins_pla_ands[20][5] ),
    .A1(net1041),
    .S(net296),
    .X(_03946_));
 sky130_fd_sc_hd__or2_1 _08185_ (.A(net511),
    .B(_03946_),
    .X(_00731_));
 sky130_fd_sc_hd__mux2_1 _08186_ (.A0(\tms1x00.ins_pla_ands[20][6] ),
    .A1(net1033),
    .S(net296),
    .X(_03947_));
 sky130_fd_sc_hd__or2_1 _08187_ (.A(net513),
    .B(_03947_),
    .X(_00732_));
 sky130_fd_sc_hd__o22a_1 _08188_ (.A1(\tms1x00.ins_pla_ands[20][7] ),
    .A2(net296),
    .B1(_03722_),
    .B2(net367),
    .X(_00733_));
 sky130_fd_sc_hd__mux2_1 _08189_ (.A0(\tms1x00.ins_pla_ands[20][8] ),
    .A1(net1014),
    .S(net296),
    .X(_03948_));
 sky130_fd_sc_hd__or2_1 _08190_ (.A(net513),
    .B(_03948_),
    .X(_00734_));
 sky130_fd_sc_hd__o22a_1 _08191_ (.A1(\tms1x00.ins_pla_ands[20][9] ),
    .A2(net296),
    .B1(_03722_),
    .B2(net364),
    .X(_00735_));
 sky130_fd_sc_hd__mux2_1 _08192_ (.A0(\tms1x00.ins_pla_ands[20][12] ),
    .A1(net963),
    .S(net296),
    .X(_03949_));
 sky130_fd_sc_hd__or2_1 _08193_ (.A(net513),
    .B(_03949_),
    .X(_00736_));
 sky130_fd_sc_hd__o22a_1 _08194_ (.A1(\tms1x00.ins_pla_ands[20][13] ),
    .A2(net296),
    .B1(_03722_),
    .B2(net363),
    .X(_00737_));
 sky130_fd_sc_hd__mux2_1 _08195_ (.A0(\tms1x00.ins_pla_ands[20][14] ),
    .A1(net951),
    .S(net296),
    .X(_03950_));
 sky130_fd_sc_hd__or2_1 _08196_ (.A(net514),
    .B(_03950_),
    .X(_00738_));
 sky130_fd_sc_hd__mux2_1 _08197_ (.A0(\tms1x00.ins_pla_ands[20][15] ),
    .A1(net944),
    .S(net296),
    .X(_03951_));
 sky130_fd_sc_hd__and2_1 _08198_ (.A(net459),
    .B(_03951_),
    .X(_00739_));
 sky130_fd_sc_hd__and3_4 _08199_ (.A(net876),
    .B(net351),
    .C(net596),
    .X(_03952_));
 sky130_fd_sc_hd__or3_2 _08200_ (.A(net856),
    .B(net348),
    .C(net594),
    .X(_03953_));
 sky130_fd_sc_hd__mux2_1 _08201_ (.A0(net976),
    .A1(\tms1x00.ins_pla_ands[11][0] ),
    .S(net270),
    .X(_03954_));
 sky130_fd_sc_hd__or2_1 _08202_ (.A(net526),
    .B(_03954_),
    .X(_00740_));
 sky130_fd_sc_hd__or2_1 _08203_ (.A(\tms1x00.ins_pla_ands[11][1] ),
    .B(_03952_),
    .X(_03955_));
 sky130_fd_sc_hd__o211a_1 _08204_ (.A1(net928),
    .A2(net270),
    .B1(_03955_),
    .C1(net464),
    .X(_00741_));
 sky130_fd_sc_hd__or2_1 _08205_ (.A(\tms1x00.ins_pla_ands[11][2] ),
    .B(_03952_),
    .X(_03956_));
 sky130_fd_sc_hd__o211a_1 _08206_ (.A1(net1065),
    .A2(net270),
    .B1(_03956_),
    .C1(net468),
    .X(_00742_));
 sky130_fd_sc_hd__mux2_1 _08207_ (.A0(net1054),
    .A1(\tms1x00.ins_pla_ands[11][3] ),
    .S(net270),
    .X(_03957_));
 sky130_fd_sc_hd__or2_1 _08208_ (.A(net530),
    .B(_03957_),
    .X(_00743_));
 sky130_fd_sc_hd__or2_1 _08209_ (.A(\tms1x00.ins_pla_ands[11][4] ),
    .B(_03952_),
    .X(_03958_));
 sky130_fd_sc_hd__o211a_1 _08210_ (.A1(net1047),
    .A2(net271),
    .B1(_03958_),
    .C1(net464),
    .X(_00744_));
 sky130_fd_sc_hd__mux2_1 _08211_ (.A0(net1038),
    .A1(\tms1x00.ins_pla_ands[11][5] ),
    .S(net271),
    .X(_03959_));
 sky130_fd_sc_hd__or2_1 _08212_ (.A(net530),
    .B(_03959_),
    .X(_00745_));
 sky130_fd_sc_hd__mux2_1 _08213_ (.A0(net1015),
    .A1(\tms1x00.ins_pla_ands[11][8] ),
    .S(net270),
    .X(_03960_));
 sky130_fd_sc_hd__or2_1 _08214_ (.A(net526),
    .B(_03960_),
    .X(_00746_));
 sky130_fd_sc_hd__or2_1 _08215_ (.A(\tms1x00.ins_pla_ands[11][9] ),
    .B(_03952_),
    .X(_03961_));
 sky130_fd_sc_hd__o211a_1 _08216_ (.A1(net1008),
    .A2(net270),
    .B1(_03961_),
    .C1(net464),
    .X(_00747_));
 sky130_fd_sc_hd__or2_1 _08217_ (.A(\tms1x00.ins_pla_ands[11][10] ),
    .B(_03952_),
    .X(_03962_));
 sky130_fd_sc_hd__o211a_1 _08218_ (.A1(net973),
    .A2(net271),
    .B1(_03962_),
    .C1(net466),
    .X(_00748_));
 sky130_fd_sc_hd__mux2_1 _08219_ (.A0(net969),
    .A1(\tms1x00.ins_pla_ands[11][11] ),
    .S(net271),
    .X(_03963_));
 sky130_fd_sc_hd__or2_1 _08220_ (.A(net530),
    .B(_03963_),
    .X(_00749_));
 sky130_fd_sc_hd__mux2_1 _08221_ (.A0(net964),
    .A1(\tms1x00.ins_pla_ands[11][12] ),
    .S(net270),
    .X(_03964_));
 sky130_fd_sc_hd__or2_1 _08222_ (.A(net526),
    .B(_03964_),
    .X(_00750_));
 sky130_fd_sc_hd__or2_1 _08223_ (.A(\tms1x00.ins_pla_ands[11][13] ),
    .B(_03952_),
    .X(_03965_));
 sky130_fd_sc_hd__o211a_1 _08224_ (.A1(net959),
    .A2(net270),
    .B1(_03965_),
    .C1(net464),
    .X(_00751_));
 sky130_fd_sc_hd__mux2_1 _08225_ (.A0(net952),
    .A1(\tms1x00.ins_pla_ands[11][14] ),
    .S(net270),
    .X(_03966_));
 sky130_fd_sc_hd__or2_1 _08226_ (.A(net526),
    .B(_03966_),
    .X(_00752_));
 sky130_fd_sc_hd__or2_1 _08227_ (.A(\tms1x00.ins_pla_ands[11][15] ),
    .B(_03952_),
    .X(_03967_));
 sky130_fd_sc_hd__o211a_1 _08228_ (.A1(net946),
    .A2(net270),
    .B1(_03967_),
    .C1(net464),
    .X(_00753_));
 sky130_fd_sc_hd__and3_4 _08229_ (.A(net766),
    .B(net352),
    .C(net708),
    .X(_03968_));
 sky130_fd_sc_hd__or3_4 _08230_ (.A(net752),
    .B(_03470_),
    .C(net707),
    .X(_03969_));
 sky130_fd_sc_hd__or2_1 _08231_ (.A(\tms1x00.ins_pla_ands[1][0] ),
    .B(_03968_),
    .X(_03970_));
 sky130_fd_sc_hd__o211a_1 _08232_ (.A1(net977),
    .A2(_03969_),
    .B1(_03970_),
    .C1(net469),
    .X(_00754_));
 sky130_fd_sc_hd__or2_1 _08233_ (.A(\tms1x00.ins_pla_ands[1][3] ),
    .B(_03968_),
    .X(_03971_));
 sky130_fd_sc_hd__o211a_1 _08234_ (.A1(net1056),
    .A2(_03969_),
    .B1(_03971_),
    .C1(net469),
    .X(_00755_));
 sky130_fd_sc_hd__or2_1 _08235_ (.A(\tms1x00.ins_pla_ands[1][5] ),
    .B(_03968_),
    .X(_03972_));
 sky130_fd_sc_hd__o211a_1 _08236_ (.A1(net1040),
    .A2(_03969_),
    .B1(_03972_),
    .C1(net469),
    .X(_00756_));
 sky130_fd_sc_hd__or2_1 _08237_ (.A(\tms1x00.ins_pla_ands[1][6] ),
    .B(_03968_),
    .X(_03973_));
 sky130_fd_sc_hd__o211a_1 _08238_ (.A1(net1031),
    .A2(_03969_),
    .B1(_03973_),
    .C1(net469),
    .X(_00757_));
 sky130_fd_sc_hd__mux2_1 _08239_ (.A0(net954),
    .A1(\tms1x00.ins_pla_ands[1][14] ),
    .S(_03969_),
    .X(_03974_));
 sky130_fd_sc_hd__or2_1 _08240_ (.A(net531),
    .B(_03974_),
    .X(_00758_));
 sky130_fd_sc_hd__nand2_1 _08241_ (.A(_01632_),
    .B(_03969_),
    .Y(_03975_));
 sky130_fd_sc_hd__o211a_1 _08242_ (.A1(net946),
    .A2(_03969_),
    .B1(_03975_),
    .C1(net475),
    .X(_00759_));
 sky130_fd_sc_hd__or4_4 _08243_ (.A(net905),
    .B(_01637_),
    .C(_03348_),
    .D(_03350_),
    .X(_03976_));
 sky130_fd_sc_hd__nor2_8 _08244_ (.A(net790),
    .B(net342),
    .Y(_03977_));
 sky130_fd_sc_hd__or2_4 _08245_ (.A(net789),
    .B(net342),
    .X(_03978_));
 sky130_fd_sc_hd__or2_1 _08246_ (.A(\tms1x00.O_pla_ors[7][0] ),
    .B(_03977_),
    .X(_03979_));
 sky130_fd_sc_hd__o211a_1 _08247_ (.A1(net980),
    .A2(net268),
    .B1(_03979_),
    .C1(net507),
    .X(_00760_));
 sky130_fd_sc_hd__or2_1 _08248_ (.A(\tms1x00.O_pla_ors[7][1] ),
    .B(_03977_),
    .X(_03980_));
 sky130_fd_sc_hd__o211a_1 _08249_ (.A1(net932),
    .A2(net268),
    .B1(_03980_),
    .C1(net506),
    .X(_00761_));
 sky130_fd_sc_hd__mux2_1 _08250_ (.A0(net1067),
    .A1(\tms1x00.O_pla_ors[7][2] ),
    .S(net269),
    .X(_03981_));
 sky130_fd_sc_hd__or2_1 _08251_ (.A(net561),
    .B(_03981_),
    .X(_00762_));
 sky130_fd_sc_hd__mux2_1 _08252_ (.A0(net1059),
    .A1(\tms1x00.O_pla_ors[7][3] ),
    .S(net269),
    .X(_03982_));
 sky130_fd_sc_hd__or2_1 _08253_ (.A(net557),
    .B(_03982_),
    .X(_00763_));
 sky130_fd_sc_hd__mux2_1 _08254_ (.A0(net1050),
    .A1(\tms1x00.O_pla_ors[7][4] ),
    .S(net269),
    .X(_03983_));
 sky130_fd_sc_hd__or2_1 _08255_ (.A(net558),
    .B(_03983_),
    .X(_00764_));
 sky130_fd_sc_hd__mux2_1 _08256_ (.A0(net1042),
    .A1(\tms1x00.O_pla_ors[7][5] ),
    .S(net268),
    .X(_03984_));
 sky130_fd_sc_hd__or2_1 _08257_ (.A(net576),
    .B(_03984_),
    .X(_00765_));
 sky130_fd_sc_hd__mux2_1 _08258_ (.A0(net1035),
    .A1(\tms1x00.O_pla_ors[7][6] ),
    .S(net268),
    .X(_03985_));
 sky130_fd_sc_hd__or2_1 _08259_ (.A(net570),
    .B(_03985_),
    .X(_00766_));
 sky130_fd_sc_hd__or2_1 _08260_ (.A(\tms1x00.O_pla_ors[7][7] ),
    .B(_03977_),
    .X(_03986_));
 sky130_fd_sc_hd__o211a_1 _08261_ (.A1(net1027),
    .A2(net268),
    .B1(_03986_),
    .C1(net502),
    .X(_00767_));
 sky130_fd_sc_hd__mux2_1 _08262_ (.A0(net1019),
    .A1(\tms1x00.O_pla_ors[7][8] ),
    .S(net269),
    .X(_03987_));
 sky130_fd_sc_hd__or2_1 _08263_ (.A(net556),
    .B(_03987_),
    .X(_00768_));
 sky130_fd_sc_hd__mux2_1 _08264_ (.A0(net1011),
    .A1(\tms1x00.O_pla_ors[7][9] ),
    .S(net269),
    .X(_03988_));
 sky130_fd_sc_hd__or2_1 _08265_ (.A(net572),
    .B(_03988_),
    .X(_00769_));
 sky130_fd_sc_hd__mux2_1 _08266_ (.A0(net974),
    .A1(\tms1x00.O_pla_ors[7][10] ),
    .S(net268),
    .X(_03989_));
 sky130_fd_sc_hd__or2_1 _08267_ (.A(net572),
    .B(_03989_),
    .X(_00770_));
 sky130_fd_sc_hd__mux2_1 _08268_ (.A0(net970),
    .A1(\tms1x00.O_pla_ors[7][11] ),
    .S(net269),
    .X(_03990_));
 sky130_fd_sc_hd__or2_1 _08269_ (.A(net561),
    .B(_03990_),
    .X(_00771_));
 sky130_fd_sc_hd__or2_1 _08270_ (.A(\tms1x00.O_pla_ors[7][12] ),
    .B(_03977_),
    .X(_03991_));
 sky130_fd_sc_hd__o211a_1 _08271_ (.A1(net966),
    .A2(net269),
    .B1(_03991_),
    .C1(net492),
    .X(_00772_));
 sky130_fd_sc_hd__mux2_1 _08272_ (.A0(net962),
    .A1(\tms1x00.O_pla_ors[7][13] ),
    .S(net269),
    .X(_03992_));
 sky130_fd_sc_hd__or2_1 _08273_ (.A(net556),
    .B(_03992_),
    .X(_00773_));
 sky130_fd_sc_hd__mux2_1 _08274_ (.A0(net955),
    .A1(\tms1x00.O_pla_ors[7][14] ),
    .S(net268),
    .X(_03993_));
 sky130_fd_sc_hd__or2_1 _08275_ (.A(net568),
    .B(_03993_),
    .X(_00774_));
 sky130_fd_sc_hd__mux2_1 _08276_ (.A0(net949),
    .A1(\tms1x00.O_pla_ors[7][15] ),
    .S(net268),
    .X(_03994_));
 sky130_fd_sc_hd__or2_1 _08277_ (.A(net567),
    .B(_03994_),
    .X(_00775_));
 sky130_fd_sc_hd__or2_1 _08278_ (.A(\tms1x00.O_pla_ors[7][16] ),
    .B(_03977_),
    .X(_03995_));
 sky130_fd_sc_hd__o211a_1 _08279_ (.A1(net943),
    .A2(net268),
    .B1(_03995_),
    .C1(net502),
    .X(_00776_));
 sky130_fd_sc_hd__or2_1 _08280_ (.A(\tms1x00.O_pla_ors[7][17] ),
    .B(_03977_),
    .X(_03996_));
 sky130_fd_sc_hd__o211a_1 _08281_ (.A1(net941),
    .A2(net269),
    .B1(_03996_),
    .C1(net491),
    .X(_00777_));
 sky130_fd_sc_hd__or2_1 _08282_ (.A(\tms1x00.O_pla_ors[7][18] ),
    .B(_03977_),
    .X(_03997_));
 sky130_fd_sc_hd__o211a_1 _08283_ (.A1(net939),
    .A2(_03978_),
    .B1(_03997_),
    .C1(net506),
    .X(_00778_));
 sky130_fd_sc_hd__or2_1 _08284_ (.A(\tms1x00.O_pla_ors[7][19] ),
    .B(_03977_),
    .X(_03998_));
 sky130_fd_sc_hd__o211a_1 _08285_ (.A1(net935),
    .A2(net268),
    .B1(_03998_),
    .C1(net502),
    .X(_00779_));
 sky130_fd_sc_hd__and3_4 _08286_ (.A(net739),
    .B(net598),
    .C(net351),
    .X(_03999_));
 sky130_fd_sc_hd__nor2_1 _08287_ (.A(net516),
    .B(_03999_),
    .Y(_04000_));
 sky130_fd_sc_hd__or2_4 _08288_ (.A(net516),
    .B(_03999_),
    .X(_04001_));
 sky130_fd_sc_hd__mux2_1 _08289_ (.A0(\tms1x00.ins_pla_ands[18][0] ),
    .A1(_03476_),
    .S(_04001_),
    .X(_00780_));
 sky130_fd_sc_hd__mux2_1 _08290_ (.A0(\tms1x00.ins_pla_ands[18][1] ),
    .A1(net354),
    .S(_04001_),
    .X(_00781_));
 sky130_fd_sc_hd__mux2_1 _08291_ (.A0(\tms1x00.ins_pla_ands[18][2] ),
    .A1(_03477_),
    .S(_04001_),
    .X(_00782_));
 sky130_fd_sc_hd__mux2_1 _08292_ (.A0(\tms1x00.ins_pla_ands[18][3] ),
    .A1(_03534_),
    .S(_04001_),
    .X(_00783_));
 sky130_fd_sc_hd__mux2_1 _08293_ (.A0(\tms1x00.ins_pla_ands[18][4] ),
    .A1(_03479_),
    .S(_04001_),
    .X(_00784_));
 sky130_fd_sc_hd__mux2_1 _08294_ (.A0(\tms1x00.ins_pla_ands[18][5] ),
    .A1(_03712_),
    .S(_04001_),
    .X(_00785_));
 sky130_fd_sc_hd__mux2_1 _08295_ (.A0(\tms1x00.ins_pla_ands[18][6] ),
    .A1(_03435_),
    .S(_04001_),
    .X(_00786_));
 sky130_fd_sc_hd__mux2_1 _08296_ (.A0(\tms1x00.ins_pla_ands[18][7] ),
    .A1(_03536_),
    .S(_04001_),
    .X(_00787_));
 sky130_fd_sc_hd__mux2_1 _08297_ (.A0(\tms1x00.ins_pla_ands[18][10] ),
    .A1(_03482_),
    .S(_04001_),
    .X(_00788_));
 sky130_fd_sc_hd__mux2_1 _08298_ (.A0(\tms1x00.ins_pla_ands[18][11] ),
    .A1(net347),
    .S(_04001_),
    .X(_00789_));
 sky130_fd_sc_hd__and3_4 _08299_ (.A(net795),
    .B(net352),
    .C(net596),
    .X(_04002_));
 sky130_fd_sc_hd__or3_4 _08300_ (.A(net778),
    .B(net349),
    .C(net594),
    .X(_04003_));
 sky130_fd_sc_hd__nor2_1 _08301_ (.A(net376),
    .B(_04002_),
    .Y(_04004_));
 sky130_fd_sc_hd__nand2_1 _08302_ (.A(net369),
    .B(net267),
    .Y(_04005_));
 sky130_fd_sc_hd__nor2_1 _08303_ (.A(net391),
    .B(_04002_),
    .Y(_04006_));
 sky130_fd_sc_hd__nand2_1 _08304_ (.A(net383),
    .B(net267),
    .Y(_04007_));
 sky130_fd_sc_hd__a22o_1 _08305_ (.A1(\tms1x00.ins_pla_ands[15][0] ),
    .A2(_04004_),
    .B1(_04007_),
    .B2(net343),
    .X(_00790_));
 sky130_fd_sc_hd__o22a_1 _08306_ (.A1(\tms1x00.ins_pla_ands[15][1] ),
    .A2(_04005_),
    .B1(_04006_),
    .B2(net344),
    .X(_00791_));
 sky130_fd_sc_hd__o22a_1 _08307_ (.A1(\tms1x00.ins_pla_ands[15][2] ),
    .A2(_04005_),
    .B1(_04006_),
    .B2(_03477_),
    .X(_00792_));
 sky130_fd_sc_hd__a22o_1 _08308_ (.A1(\tms1x00.ins_pla_ands[15][3] ),
    .A2(_04004_),
    .B1(_04007_),
    .B2(_03534_),
    .X(_00793_));
 sky130_fd_sc_hd__o22a_1 _08309_ (.A1(\tms1x00.ins_pla_ands[15][6] ),
    .A2(_04005_),
    .B1(_04006_),
    .B2(_03480_),
    .X(_00794_));
 sky130_fd_sc_hd__a22o_1 _08310_ (.A1(\tms1x00.ins_pla_ands[15][7] ),
    .A2(_04004_),
    .B1(_04007_),
    .B2(_03437_),
    .X(_00795_));
 sky130_fd_sc_hd__or3_4 _08311_ (.A(net777),
    .B(net361),
    .C(net710),
    .X(_04008_));
 sky130_fd_sc_hd__mux2_1 _08312_ (.A0(net976),
    .A1(\tms1x00.O_pla_ands[31][0] ),
    .S(_04008_),
    .X(_00796_));
 sky130_fd_sc_hd__mux2_1 _08313_ (.A0(net927),
    .A1(\tms1x00.O_pla_ands[31][1] ),
    .S(_04008_),
    .X(_00797_));
 sky130_fd_sc_hd__mux2_1 _08314_ (.A0(net1063),
    .A1(\tms1x00.O_pla_ands[31][2] ),
    .S(_04008_),
    .X(_00798_));
 sky130_fd_sc_hd__mux2_1 _08315_ (.A0(net1054),
    .A1(\tms1x00.O_pla_ands[31][3] ),
    .S(_04008_),
    .X(_00799_));
 sky130_fd_sc_hd__mux2_1 _08316_ (.A0(net1046),
    .A1(\tms1x00.O_pla_ands[31][4] ),
    .S(_04008_),
    .X(_00800_));
 sky130_fd_sc_hd__mux2_1 _08317_ (.A0(net1038),
    .A1(\tms1x00.O_pla_ands[31][5] ),
    .S(_04008_),
    .X(_00801_));
 sky130_fd_sc_hd__mux2_1 _08318_ (.A0(net1030),
    .A1(\tms1x00.O_pla_ands[31][6] ),
    .S(_04008_),
    .X(_00802_));
 sky130_fd_sc_hd__mux2_1 _08319_ (.A0(net1024),
    .A1(\tms1x00.O_pla_ands[31][7] ),
    .S(_04008_),
    .X(_00803_));
 sky130_fd_sc_hd__mux2_1 _08320_ (.A0(net1015),
    .A1(\tms1x00.O_pla_ands[31][8] ),
    .S(_04008_),
    .X(_00804_));
 sky130_fd_sc_hd__mux2_1 _08321_ (.A0(net1007),
    .A1(\tms1x00.O_pla_ands[31][9] ),
    .S(_04008_),
    .X(_00805_));
 sky130_fd_sc_hd__nor2_4 _08322_ (.A(net378),
    .B(_03968_),
    .Y(_04009_));
 sky130_fd_sc_hd__nand2_1 _08323_ (.A(net370),
    .B(_03969_),
    .Y(_04010_));
 sky130_fd_sc_hd__nor2_1 _08324_ (.A(net392),
    .B(_03968_),
    .Y(_04011_));
 sky130_fd_sc_hd__nand2_4 _08325_ (.A(net384),
    .B(_03969_),
    .Y(_04012_));
 sky130_fd_sc_hd__a22o_1 _08326_ (.A1(\tms1x00.ins_pla_ands[1][1] ),
    .A2(_04009_),
    .B1(_04012_),
    .B2(net354),
    .X(_00806_));
 sky130_fd_sc_hd__a22o_1 _08327_ (.A1(\tms1x00.ins_pla_ands[1][2] ),
    .A2(_04009_),
    .B1(_04012_),
    .B2(_03429_),
    .X(_00807_));
 sky130_fd_sc_hd__a22o_1 _08328_ (.A1(\tms1x00.ins_pla_ands[1][4] ),
    .A2(_04009_),
    .B1(_04012_),
    .B2(_03535_),
    .X(_00808_));
 sky130_fd_sc_hd__a22o_1 _08329_ (.A1(\tms1x00.ins_pla_ands[1][7] ),
    .A2(_04009_),
    .B1(_04012_),
    .B2(_03437_),
    .X(_00809_));
 sky130_fd_sc_hd__a22o_1 _08330_ (.A1(\tms1x00.ins_pla_ands[1][8] ),
    .A2(_04009_),
    .B1(_04012_),
    .B2(net353),
    .X(_00810_));
 sky130_fd_sc_hd__o22a_1 _08331_ (.A1(\tms1x00.ins_pla_ands[1][9] ),
    .A2(_04010_),
    .B1(_04011_),
    .B2(_03578_),
    .X(_00811_));
 sky130_fd_sc_hd__a22o_1 _08332_ (.A1(\tms1x00.ins_pla_ands[1][10] ),
    .A2(_04009_),
    .B1(_04012_),
    .B2(_03579_),
    .X(_00812_));
 sky130_fd_sc_hd__o22a_1 _08333_ (.A1(\tms1x00.ins_pla_ands[1][11] ),
    .A2(_04010_),
    .B1(_04011_),
    .B2(_03580_),
    .X(_00813_));
 sky130_fd_sc_hd__a22o_1 _08334_ (.A1(\tms1x00.ins_pla_ands[1][12] ),
    .A2(_04009_),
    .B1(_04012_),
    .B2(_03588_),
    .X(_00814_));
 sky130_fd_sc_hd__o22a_1 _08335_ (.A1(\tms1x00.ins_pla_ands[1][13] ),
    .A2(_04010_),
    .B1(_04011_),
    .B2(_03589_),
    .X(_00815_));
 sky130_fd_sc_hd__or2_1 _08336_ (.A(\tms1x00.ins_pla_ands[10][0] ),
    .B(_03911_),
    .X(_04013_));
 sky130_fd_sc_hd__o211a_1 _08337_ (.A1(net976),
    .A2(net276),
    .B1(_04013_),
    .C1(net464),
    .X(_00816_));
 sky130_fd_sc_hd__mux2_1 _08338_ (.A0(net928),
    .A1(\tms1x00.ins_pla_ands[10][1] ),
    .S(net276),
    .X(_04014_));
 sky130_fd_sc_hd__or2_1 _08339_ (.A(net530),
    .B(_04014_),
    .X(_00817_));
 sky130_fd_sc_hd__or2_1 _08340_ (.A(\tms1x00.ins_pla_ands[10][2] ),
    .B(_03911_),
    .X(_04015_));
 sky130_fd_sc_hd__o211a_1 _08341_ (.A1(net1065),
    .A2(net276),
    .B1(_04015_),
    .C1(net468),
    .X(_00818_));
 sky130_fd_sc_hd__mux2_1 _08342_ (.A0(net1054),
    .A1(\tms1x00.ins_pla_ands[10][3] ),
    .S(net276),
    .X(_04016_));
 sky130_fd_sc_hd__or2_1 _08343_ (.A(net530),
    .B(_04016_),
    .X(_00819_));
 sky130_fd_sc_hd__or2_1 _08344_ (.A(\tms1x00.ins_pla_ands[10][4] ),
    .B(_03911_),
    .X(_04017_));
 sky130_fd_sc_hd__o211a_1 _08345_ (.A1(net1047),
    .A2(net276),
    .B1(_04017_),
    .C1(net465),
    .X(_00820_));
 sky130_fd_sc_hd__mux2_1 _08346_ (.A0(net1038),
    .A1(\tms1x00.ins_pla_ands[10][5] ),
    .S(net277),
    .X(_04018_));
 sky130_fd_sc_hd__or2_1 _08347_ (.A(net530),
    .B(_04018_),
    .X(_00821_));
 sky130_fd_sc_hd__mux2_1 _08348_ (.A0(net1015),
    .A1(\tms1x00.ins_pla_ands[10][8] ),
    .S(net277),
    .X(_04019_));
 sky130_fd_sc_hd__or2_1 _08349_ (.A(net527),
    .B(_04019_),
    .X(_00822_));
 sky130_fd_sc_hd__or2_1 _08350_ (.A(\tms1x00.ins_pla_ands[10][9] ),
    .B(_03911_),
    .X(_04020_));
 sky130_fd_sc_hd__o211a_1 _08351_ (.A1(net1008),
    .A2(net276),
    .B1(_04020_),
    .C1(net464),
    .X(_00823_));
 sky130_fd_sc_hd__or2_1 _08352_ (.A(\tms1x00.ins_pla_ands[10][10] ),
    .B(_03911_),
    .X(_04021_));
 sky130_fd_sc_hd__o211a_1 _08353_ (.A1(net973),
    .A2(net277),
    .B1(_04021_),
    .C1(net466),
    .X(_00824_));
 sky130_fd_sc_hd__mux2_1 _08354_ (.A0(net969),
    .A1(\tms1x00.ins_pla_ands[10][11] ),
    .S(net277),
    .X(_04022_));
 sky130_fd_sc_hd__or2_1 _08355_ (.A(net530),
    .B(_04022_),
    .X(_00825_));
 sky130_fd_sc_hd__mux2_1 _08356_ (.A0(net964),
    .A1(\tms1x00.ins_pla_ands[10][12] ),
    .S(net276),
    .X(_04023_));
 sky130_fd_sc_hd__or2_1 _08357_ (.A(net526),
    .B(_04023_),
    .X(_00826_));
 sky130_fd_sc_hd__or2_1 _08358_ (.A(\tms1x00.ins_pla_ands[10][13] ),
    .B(_03911_),
    .X(_04024_));
 sky130_fd_sc_hd__o211a_1 _08359_ (.A1(net959),
    .A2(net276),
    .B1(_04024_),
    .C1(net468),
    .X(_00827_));
 sky130_fd_sc_hd__mux2_1 _08360_ (.A0(net952),
    .A1(\tms1x00.ins_pla_ands[10][14] ),
    .S(net276),
    .X(_04025_));
 sky130_fd_sc_hd__or2_1 _08361_ (.A(net527),
    .B(_04025_),
    .X(_00828_));
 sky130_fd_sc_hd__or2_1 _08362_ (.A(\tms1x00.ins_pla_ands[10][15] ),
    .B(_03911_),
    .X(_04026_));
 sky130_fd_sc_hd__o211a_1 _08363_ (.A1(net946),
    .A2(net276),
    .B1(_04026_),
    .C1(net468),
    .X(_00829_));
 sky130_fd_sc_hd__and3_2 _08364_ (.A(net847),
    .B(net351),
    .C(net708),
    .X(_04027_));
 sky130_fd_sc_hd__or3_2 _08365_ (.A(net835),
    .B(net349),
    .C(net707),
    .X(_04028_));
 sky130_fd_sc_hd__or2_1 _08366_ (.A(\tms1x00.ins_pla_ands[0][2] ),
    .B(_04027_),
    .X(_04029_));
 sky130_fd_sc_hd__o211a_1 _08367_ (.A1(net1071),
    .A2(net266),
    .B1(_04029_),
    .C1(net470),
    .X(_00830_));
 sky130_fd_sc_hd__mux2_1 _08368_ (.A0(net1056),
    .A1(\tms1x00.ins_pla_ands[0][3] ),
    .S(net266),
    .X(_04030_));
 sky130_fd_sc_hd__or2_1 _08369_ (.A(net535),
    .B(_04030_),
    .X(_00831_));
 sky130_fd_sc_hd__or2_1 _08370_ (.A(\tms1x00.ins_pla_ands[0][4] ),
    .B(_04027_),
    .X(_04031_));
 sky130_fd_sc_hd__o211a_1 _08371_ (.A1(net1048),
    .A2(net266),
    .B1(_04031_),
    .C1(net470),
    .X(_00832_));
 sky130_fd_sc_hd__mux2_1 _08372_ (.A0(net1040),
    .A1(\tms1x00.ins_pla_ands[0][5] ),
    .S(net266),
    .X(_04032_));
 sky130_fd_sc_hd__or2_1 _08373_ (.A(net535),
    .B(_04032_),
    .X(_00833_));
 sky130_fd_sc_hd__or2_1 _08374_ (.A(\tms1x00.ins_pla_ands[0][6] ),
    .B(_04027_),
    .X(_04033_));
 sky130_fd_sc_hd__o211a_1 _08375_ (.A1(net1031),
    .A2(net266),
    .B1(_04033_),
    .C1(net470),
    .X(_00834_));
 sky130_fd_sc_hd__mux2_1 _08376_ (.A0(net1025),
    .A1(\tms1x00.ins_pla_ands[0][7] ),
    .S(net266),
    .X(_04034_));
 sky130_fd_sc_hd__or2_1 _08377_ (.A(net535),
    .B(_04034_),
    .X(_00835_));
 sky130_fd_sc_hd__mux2_1 _08378_ (.A0(net954),
    .A1(\tms1x00.ins_pla_ands[0][14] ),
    .S(net266),
    .X(_04035_));
 sky130_fd_sc_hd__or2_1 _08379_ (.A(net534),
    .B(_04035_),
    .X(_00836_));
 sky130_fd_sc_hd__nand2_1 _08380_ (.A(_01631_),
    .B(net266),
    .Y(_04036_));
 sky130_fd_sc_hd__o211a_1 _08381_ (.A1(net947),
    .A2(_04028_),
    .B1(_04036_),
    .C1(net472),
    .X(_00837_));
 sky130_fd_sc_hd__nor2_8 _08382_ (.A(net624),
    .B(net341),
    .Y(_04037_));
 sky130_fd_sc_hd__or2_4 _08383_ (.A(net623),
    .B(net342),
    .X(_04038_));
 sky130_fd_sc_hd__mux2_1 _08384_ (.A0(net983),
    .A1(\tms1x00.O_pla_ors[6][0] ),
    .S(net265),
    .X(_04039_));
 sky130_fd_sc_hd__or2_1 _08385_ (.A(net569),
    .B(_04039_),
    .X(_00838_));
 sky130_fd_sc_hd__or2_1 _08386_ (.A(\tms1x00.O_pla_ors[6][1] ),
    .B(_04037_),
    .X(_04040_));
 sky130_fd_sc_hd__o211a_1 _08387_ (.A1(net932),
    .A2(net265),
    .B1(_04040_),
    .C1(net506),
    .X(_00839_));
 sky130_fd_sc_hd__or2_1 _08388_ (.A(\tms1x00.O_pla_ors[6][2] ),
    .B(_04037_),
    .X(_04041_));
 sky130_fd_sc_hd__o211a_1 _08389_ (.A1(net1067),
    .A2(net264),
    .B1(_04041_),
    .C1(net498),
    .X(_00840_));
 sky130_fd_sc_hd__or2_1 _08390_ (.A(\tms1x00.O_pla_ors[6][3] ),
    .B(_04037_),
    .X(_04042_));
 sky130_fd_sc_hd__o211a_1 _08391_ (.A1(net1059),
    .A2(net264),
    .B1(_04042_),
    .C1(net492),
    .X(_00841_));
 sky130_fd_sc_hd__mux2_1 _08392_ (.A0(net1050),
    .A1(\tms1x00.O_pla_ors[6][4] ),
    .S(net264),
    .X(_04043_));
 sky130_fd_sc_hd__or2_1 _08393_ (.A(net561),
    .B(_04043_),
    .X(_00842_));
 sky130_fd_sc_hd__mux2_1 _08394_ (.A0(net1042),
    .A1(\tms1x00.O_pla_ors[6][5] ),
    .S(net265),
    .X(_04044_));
 sky130_fd_sc_hd__or2_1 _08395_ (.A(net576),
    .B(_04044_),
    .X(_00843_));
 sky130_fd_sc_hd__mux2_1 _08396_ (.A0(net1034),
    .A1(\tms1x00.O_pla_ors[6][6] ),
    .S(net265),
    .X(_04045_));
 sky130_fd_sc_hd__or2_1 _08397_ (.A(net570),
    .B(_04045_),
    .X(_00844_));
 sky130_fd_sc_hd__or2_1 _08398_ (.A(\tms1x00.O_pla_ors[6][7] ),
    .B(_04037_),
    .X(_04046_));
 sky130_fd_sc_hd__o211a_1 _08399_ (.A1(net1027),
    .A2(net265),
    .B1(_04046_),
    .C1(net499),
    .X(_00845_));
 sky130_fd_sc_hd__mux2_1 _08400_ (.A0(net1019),
    .A1(\tms1x00.O_pla_ors[6][8] ),
    .S(net264),
    .X(_04047_));
 sky130_fd_sc_hd__or2_1 _08401_ (.A(net557),
    .B(_04047_),
    .X(_00846_));
 sky130_fd_sc_hd__mux2_1 _08402_ (.A0(net1011),
    .A1(\tms1x00.O_pla_ors[6][9] ),
    .S(net265),
    .X(_04048_));
 sky130_fd_sc_hd__or2_1 _08403_ (.A(net570),
    .B(_04048_),
    .X(_00847_));
 sky130_fd_sc_hd__mux2_1 _08404_ (.A0(net974),
    .A1(\tms1x00.O_pla_ors[6][10] ),
    .S(net265),
    .X(_04049_));
 sky130_fd_sc_hd__or2_1 _08405_ (.A(net572),
    .B(_04049_),
    .X(_00848_));
 sky130_fd_sc_hd__mux2_1 _08406_ (.A0(net970),
    .A1(\tms1x00.O_pla_ors[6][11] ),
    .S(net264),
    .X(_04050_));
 sky130_fd_sc_hd__or2_1 _08407_ (.A(net558),
    .B(_04050_),
    .X(_00849_));
 sky130_fd_sc_hd__mux2_1 _08408_ (.A0(net966),
    .A1(\tms1x00.O_pla_ors[6][12] ),
    .S(net264),
    .X(_04051_));
 sky130_fd_sc_hd__or2_1 _08409_ (.A(net556),
    .B(_04051_),
    .X(_00850_));
 sky130_fd_sc_hd__or2_1 _08410_ (.A(\tms1x00.O_pla_ors[6][13] ),
    .B(_04037_),
    .X(_04052_));
 sky130_fd_sc_hd__o211a_1 _08411_ (.A1(net962),
    .A2(net264),
    .B1(_04052_),
    .C1(net491),
    .X(_00851_));
 sky130_fd_sc_hd__mux2_1 _08412_ (.A0(net955),
    .A1(\tms1x00.O_pla_ors[6][14] ),
    .S(net264),
    .X(_04053_));
 sky130_fd_sc_hd__or2_1 _08413_ (.A(net567),
    .B(_04053_),
    .X(_00852_));
 sky130_fd_sc_hd__mux2_1 _08414_ (.A0(net949),
    .A1(\tms1x00.O_pla_ors[6][15] ),
    .S(net264),
    .X(_04054_));
 sky130_fd_sc_hd__or2_1 _08415_ (.A(net567),
    .B(_04054_),
    .X(_00853_));
 sky130_fd_sc_hd__or2_1 _08416_ (.A(\tms1x00.O_pla_ors[6][16] ),
    .B(_04037_),
    .X(_04055_));
 sky130_fd_sc_hd__o211a_1 _08417_ (.A1(net943),
    .A2(net265),
    .B1(_04055_),
    .C1(net502),
    .X(_00854_));
 sky130_fd_sc_hd__or2_1 _08418_ (.A(\tms1x00.O_pla_ors[6][17] ),
    .B(_04037_),
    .X(_04056_));
 sky130_fd_sc_hd__o211a_1 _08419_ (.A1(net941),
    .A2(net264),
    .B1(_04056_),
    .C1(net491),
    .X(_00855_));
 sky130_fd_sc_hd__or2_1 _08420_ (.A(\tms1x00.O_pla_ors[6][18] ),
    .B(_04037_),
    .X(_04057_));
 sky130_fd_sc_hd__o211a_1 _08421_ (.A1(net939),
    .A2(net265),
    .B1(_04057_),
    .C1(net507),
    .X(_00856_));
 sky130_fd_sc_hd__or2_1 _08422_ (.A(\tms1x00.O_pla_ors[6][19] ),
    .B(_04037_),
    .X(_04058_));
 sky130_fd_sc_hd__o211a_1 _08423_ (.A1(net935),
    .A2(_04038_),
    .B1(_04058_),
    .C1(net501),
    .X(_00857_));
 sky130_fd_sc_hd__nor2_2 _08424_ (.A(net377),
    .B(_03888_),
    .Y(_04059_));
 sky130_fd_sc_hd__nand2_2 _08425_ (.A(net369),
    .B(_03889_),
    .Y(_04060_));
 sky130_fd_sc_hd__nor2_2 _08426_ (.A(net392),
    .B(_03888_),
    .Y(_04061_));
 sky130_fd_sc_hd__nand2_2 _08427_ (.A(net383),
    .B(_03889_),
    .Y(_04062_));
 sky130_fd_sc_hd__a22o_1 _08428_ (.A1(\tms1x00.ins_pla_ands[13][0] ),
    .A2(_04059_),
    .B1(_04062_),
    .B2(net343),
    .X(_00858_));
 sky130_fd_sc_hd__o22a_1 _08429_ (.A1(\tms1x00.ins_pla_ands[13][1] ),
    .A2(_04060_),
    .B1(_04061_),
    .B2(net344),
    .X(_00859_));
 sky130_fd_sc_hd__a22o_1 _08430_ (.A1(\tms1x00.ins_pla_ands[13][2] ),
    .A2(_04059_),
    .B1(_04062_),
    .B2(_03429_),
    .X(_00860_));
 sky130_fd_sc_hd__o22a_1 _08431_ (.A1(\tms1x00.ins_pla_ands[13][3] ),
    .A2(_04060_),
    .B1(_04061_),
    .B2(_03433_),
    .X(_00861_));
 sky130_fd_sc_hd__o22a_1 _08432_ (.A1(\tms1x00.ins_pla_ands[13][4] ),
    .A2(_04060_),
    .B1(_04061_),
    .B2(_03479_),
    .X(_00862_));
 sky130_fd_sc_hd__a22o_1 _08433_ (.A1(\tms1x00.ins_pla_ands[13][5] ),
    .A2(_04059_),
    .B1(_04062_),
    .B2(_03712_),
    .X(_00863_));
 sky130_fd_sc_hd__o22a_1 _08434_ (.A1(\tms1x00.ins_pla_ands[13][6] ),
    .A2(_04060_),
    .B1(_04061_),
    .B2(_03480_),
    .X(_00864_));
 sky130_fd_sc_hd__a22o_1 _08435_ (.A1(\tms1x00.ins_pla_ands[13][7] ),
    .A2(_04059_),
    .B1(_04062_),
    .B2(_03437_),
    .X(_00865_));
 sky130_fd_sc_hd__nor2_2 _08436_ (.A(net377),
    .B(_04027_),
    .Y(_04063_));
 sky130_fd_sc_hd__nand2_2 _08437_ (.A(net369),
    .B(net266),
    .Y(_04064_));
 sky130_fd_sc_hd__nor2_2 _08438_ (.A(net392),
    .B(_04027_),
    .Y(_04065_));
 sky130_fd_sc_hd__nand2_2 _08439_ (.A(net384),
    .B(net266),
    .Y(_04066_));
 sky130_fd_sc_hd__a22o_1 _08440_ (.A1(\tms1x00.ins_pla_ands[0][0] ),
    .A2(_04063_),
    .B1(_04066_),
    .B2(net343),
    .X(_00866_));
 sky130_fd_sc_hd__o22a_1 _08441_ (.A1(\tms1x00.ins_pla_ands[0][1] ),
    .A2(_04064_),
    .B1(_04065_),
    .B2(net344),
    .X(_00867_));
 sky130_fd_sc_hd__a22o_1 _08442_ (.A1(\tms1x00.ins_pla_ands[0][8] ),
    .A2(_04063_),
    .B1(_04066_),
    .B2(net353),
    .X(_00868_));
 sky130_fd_sc_hd__o22a_1 _08443_ (.A1(\tms1x00.ins_pla_ands[0][9] ),
    .A2(_04064_),
    .B1(_04065_),
    .B2(_03578_),
    .X(_00869_));
 sky130_fd_sc_hd__a22o_1 _08444_ (.A1(\tms1x00.ins_pla_ands[0][10] ),
    .A2(_04063_),
    .B1(_04066_),
    .B2(_03579_),
    .X(_00870_));
 sky130_fd_sc_hd__o22a_1 _08445_ (.A1(\tms1x00.ins_pla_ands[0][11] ),
    .A2(_04064_),
    .B1(_04065_),
    .B2(_03580_),
    .X(_00871_));
 sky130_fd_sc_hd__a22o_1 _08446_ (.A1(\tms1x00.ins_pla_ands[0][12] ),
    .A2(_04063_),
    .B1(_04066_),
    .B2(_03588_),
    .X(_00872_));
 sky130_fd_sc_hd__o22a_1 _08447_ (.A1(\tms1x00.ins_pla_ands[0][13] ),
    .A2(_04064_),
    .B1(_04065_),
    .B2(_03589_),
    .X(_00873_));
 sky130_fd_sc_hd__o22a_1 _08448_ (.A1(\tms1x00.ins_pla_ands[28][0] ),
    .A2(net300),
    .B1(net217),
    .B2(_03456_),
    .X(_00874_));
 sky130_fd_sc_hd__o22a_1 _08449_ (.A1(\tms1x00.ins_pla_ands[28][1] ),
    .A2(_03714_),
    .B1(net217),
    .B2(net397),
    .X(_00875_));
 sky130_fd_sc_hd__o22a_1 _08450_ (.A1(\tms1x00.ins_pla_ands[28][2] ),
    .A2(_03714_),
    .B1(net216),
    .B2(_03428_),
    .X(_00876_));
 sky130_fd_sc_hd__o22a_1 _08451_ (.A1(\tms1x00.ins_pla_ands[28][3] ),
    .A2(net300),
    .B1(net216),
    .B2(_03430_),
    .X(_00877_));
 sky130_fd_sc_hd__o22a_1 _08452_ (.A1(\tms1x00.ins_pla_ands[28][4] ),
    .A2(net300),
    .B1(net216),
    .B2(_03478_),
    .X(_00878_));
 sky130_fd_sc_hd__o22a_1 _08453_ (.A1(\tms1x00.ins_pla_ands[28][5] ),
    .A2(net300),
    .B1(net217),
    .B2(net366),
    .X(_00879_));
 sky130_fd_sc_hd__o22a_1 _08454_ (.A1(\tms1x00.ins_pla_ands[28][6] ),
    .A2(net300),
    .B1(net216),
    .B2(_03434_),
    .X(_00880_));
 sky130_fd_sc_hd__o22a_1 _08455_ (.A1(\tms1x00.ins_pla_ands[28][7] ),
    .A2(net300),
    .B1(net216),
    .B2(net367),
    .X(_00881_));
 sky130_fd_sc_hd__o22a_1 _08456_ (.A1(\tms1x00.ins_pla_ands[28][8] ),
    .A2(net300),
    .B1(net216),
    .B2(_03438_),
    .X(_00882_));
 sky130_fd_sc_hd__o22a_1 _08457_ (.A1(\tms1x00.ins_pla_ands[28][11] ),
    .A2(_03714_),
    .B1(net217),
    .B2(_03460_),
    .X(_00883_));
 sky130_fd_sc_hd__o22a_1 _08458_ (.A1(\tms1x00.ins_pla_ands[28][12] ),
    .A2(net300),
    .B1(net216),
    .B2(_03484_),
    .X(_00884_));
 sky130_fd_sc_hd__mux2_1 _08459_ (.A0(\tms1x00.ins_pla_ands[28][15] ),
    .A1(net944),
    .S(net300),
    .X(_04067_));
 sky130_fd_sc_hd__and2_1 _08460_ (.A(net460),
    .B(_04067_),
    .X(_00885_));
 sky130_fd_sc_hd__mux2_1 _08461_ (.A0(\tms1x00.ins_pla_ands[18][8] ),
    .A1(net1014),
    .S(_03999_),
    .X(_04068_));
 sky130_fd_sc_hd__or2_1 _08462_ (.A(net515),
    .B(_04068_),
    .X(_00886_));
 sky130_fd_sc_hd__o22a_1 _08463_ (.A1(\tms1x00.ins_pla_ands[18][9] ),
    .A2(_03999_),
    .B1(_04000_),
    .B2(net364),
    .X(_00887_));
 sky130_fd_sc_hd__mux2_1 _08464_ (.A0(\tms1x00.ins_pla_ands[18][12] ),
    .A1(net964),
    .S(_03999_),
    .X(_04069_));
 sky130_fd_sc_hd__or2_1 _08465_ (.A(net515),
    .B(_04069_),
    .X(_00888_));
 sky130_fd_sc_hd__o22a_1 _08466_ (.A1(\tms1x00.ins_pla_ands[18][13] ),
    .A2(_03999_),
    .B1(_04000_),
    .B2(net363),
    .X(_00889_));
 sky130_fd_sc_hd__mux2_1 _08467_ (.A0(\tms1x00.ins_pla_ands[18][14] ),
    .A1(net952),
    .S(_03999_),
    .X(_04070_));
 sky130_fd_sc_hd__or2_1 _08468_ (.A(net515),
    .B(_04070_),
    .X(_00890_));
 sky130_fd_sc_hd__or4_2 _08469_ (.A(net946),
    .B(net715),
    .C(_03353_),
    .D(net348),
    .X(_04071_));
 sky130_fd_sc_hd__o211a_1 _08470_ (.A1(\tms1x00.ins_pla_ands[18][15] ),
    .A2(_03999_),
    .B1(_04071_),
    .C1(net459),
    .X(_00891_));
 sky130_fd_sc_hd__and3_4 _08471_ (.A(net766),
    .B(net352),
    .C(net596),
    .X(_04072_));
 sky130_fd_sc_hd__or3_2 _08472_ (.A(net749),
    .B(net349),
    .C(net594),
    .X(_04073_));
 sky130_fd_sc_hd__or2_1 _08473_ (.A(\tms1x00.ins_pla_ands[9][0] ),
    .B(_04072_),
    .X(_04074_));
 sky130_fd_sc_hd__o211a_1 _08474_ (.A1(net977),
    .A2(net262),
    .B1(_04074_),
    .C1(net468),
    .X(_00892_));
 sky130_fd_sc_hd__or2_1 _08475_ (.A(\tms1x00.ins_pla_ands[9][1] ),
    .B(_04072_),
    .X(_04075_));
 sky130_fd_sc_hd__o211a_1 _08476_ (.A1(net928),
    .A2(net262),
    .B1(_04075_),
    .C1(net468),
    .X(_00893_));
 sky130_fd_sc_hd__or2_1 _08477_ (.A(\tms1x00.ins_pla_ands[9][2] ),
    .B(_04072_),
    .X(_04076_));
 sky130_fd_sc_hd__o211a_1 _08478_ (.A1(net1065),
    .A2(net263),
    .B1(_04076_),
    .C1(net471),
    .X(_00894_));
 sky130_fd_sc_hd__or2_1 _08479_ (.A(\tms1x00.ins_pla_ands[9][3] ),
    .B(_04072_),
    .X(_04077_));
 sky130_fd_sc_hd__o211a_1 _08480_ (.A1(net1056),
    .A2(net263),
    .B1(_04077_),
    .C1(net471),
    .X(_00895_));
 sky130_fd_sc_hd__mux2_1 _08481_ (.A0(net1046),
    .A1(\tms1x00.ins_pla_ands[9][4] ),
    .S(net262),
    .X(_04078_));
 sky130_fd_sc_hd__or2_1 _08482_ (.A(net530),
    .B(_04078_),
    .X(_00896_));
 sky130_fd_sc_hd__or2_1 _08483_ (.A(\tms1x00.ins_pla_ands[9][5] ),
    .B(_04072_),
    .X(_04079_));
 sky130_fd_sc_hd__o211a_1 _08484_ (.A1(net1039),
    .A2(net262),
    .B1(_04079_),
    .C1(net466),
    .X(_00897_));
 sky130_fd_sc_hd__or2_1 _08485_ (.A(\tms1x00.ins_pla_ands[9][6] ),
    .B(_04072_),
    .X(_04080_));
 sky130_fd_sc_hd__o211a_1 _08486_ (.A1(net1030),
    .A2(net262),
    .B1(_04080_),
    .C1(net468),
    .X(_00898_));
 sky130_fd_sc_hd__mux2_1 _08487_ (.A0(net1024),
    .A1(\tms1x00.ins_pla_ands[9][7] ),
    .S(net262),
    .X(_04081_));
 sky130_fd_sc_hd__or2_1 _08488_ (.A(net528),
    .B(_04081_),
    .X(_00899_));
 sky130_fd_sc_hd__or2_1 _08489_ (.A(\tms1x00.ins_pla_ands[9][8] ),
    .B(_04072_),
    .X(_04082_));
 sky130_fd_sc_hd__o211a_1 _08490_ (.A1(net1015),
    .A2(net262),
    .B1(_04082_),
    .C1(net468),
    .X(_00900_));
 sky130_fd_sc_hd__mux2_1 _08491_ (.A0(net1007),
    .A1(\tms1x00.ins_pla_ands[9][9] ),
    .S(net262),
    .X(_04083_));
 sky130_fd_sc_hd__or2_1 _08492_ (.A(net530),
    .B(_04083_),
    .X(_00901_));
 sky130_fd_sc_hd__or2_1 _08493_ (.A(\tms1x00.ins_pla_ands[9][10] ),
    .B(_04072_),
    .X(_04084_));
 sky130_fd_sc_hd__o211a_1 _08494_ (.A1(net973),
    .A2(net263),
    .B1(_04084_),
    .C1(net470),
    .X(_00902_));
 sky130_fd_sc_hd__mux2_1 _08495_ (.A0(net969),
    .A1(\tms1x00.ins_pla_ands[9][11] ),
    .S(net263),
    .X(_04085_));
 sky130_fd_sc_hd__or2_1 _08496_ (.A(net534),
    .B(_04085_),
    .X(_00903_));
 sky130_fd_sc_hd__mux2_1 _08497_ (.A0(net965),
    .A1(\tms1x00.ins_pla_ands[9][12] ),
    .S(net262),
    .X(_04086_));
 sky130_fd_sc_hd__or2_1 _08498_ (.A(net528),
    .B(_04086_),
    .X(_00904_));
 sky130_fd_sc_hd__or2_1 _08499_ (.A(\tms1x00.ins_pla_ands[9][13] ),
    .B(_04072_),
    .X(_04087_));
 sky130_fd_sc_hd__o211a_1 _08500_ (.A1(net959),
    .A2(net262),
    .B1(_04087_),
    .C1(net467),
    .X(_00905_));
 sky130_fd_sc_hd__mux2_1 _08501_ (.A0(net954),
    .A1(\tms1x00.ins_pla_ands[9][14] ),
    .S(net263),
    .X(_04088_));
 sky130_fd_sc_hd__or2_1 _08502_ (.A(net535),
    .B(_04088_),
    .X(_00906_));
 sky130_fd_sc_hd__or2_1 _08503_ (.A(\tms1x00.ins_pla_ands[9][15] ),
    .B(_04072_),
    .X(_04089_));
 sky130_fd_sc_hd__o211a_1 _08504_ (.A1(net947),
    .A2(net263),
    .B1(_04089_),
    .C1(net470),
    .X(_00907_));
 sky130_fd_sc_hd__nor2_8 _08505_ (.A(net898),
    .B(net341),
    .Y(_04090_));
 sky130_fd_sc_hd__or2_4 _08506_ (.A(net898),
    .B(net341),
    .X(_04091_));
 sky130_fd_sc_hd__mux2_1 _08507_ (.A0(net980),
    .A1(\tms1x00.O_pla_ors[5][0] ),
    .S(net261),
    .X(_04092_));
 sky130_fd_sc_hd__or2_1 _08508_ (.A(net576),
    .B(_04092_),
    .X(_00908_));
 sky130_fd_sc_hd__or2_1 _08509_ (.A(\tms1x00.O_pla_ors[5][1] ),
    .B(_04090_),
    .X(_04093_));
 sky130_fd_sc_hd__o211a_1 _08510_ (.A1(net931),
    .A2(net261),
    .B1(_04093_),
    .C1(net506),
    .X(_00909_));
 sky130_fd_sc_hd__mux2_1 _08511_ (.A0(net1068),
    .A1(\tms1x00.O_pla_ors[5][2] ),
    .S(net260),
    .X(_04094_));
 sky130_fd_sc_hd__or2_1 _08512_ (.A(net562),
    .B(_04094_),
    .X(_00910_));
 sky130_fd_sc_hd__or2_1 _08513_ (.A(\tms1x00.O_pla_ors[5][3] ),
    .B(_04090_),
    .X(_04095_));
 sky130_fd_sc_hd__o211a_1 _08514_ (.A1(net1060),
    .A2(net260),
    .B1(_04095_),
    .C1(net498),
    .X(_00911_));
 sky130_fd_sc_hd__or2_1 _08515_ (.A(\tms1x00.O_pla_ors[5][4] ),
    .B(_04090_),
    .X(_04096_));
 sky130_fd_sc_hd__o211a_1 _08516_ (.A1(net1052),
    .A2(net260),
    .B1(_04096_),
    .C1(net491),
    .X(_00912_));
 sky130_fd_sc_hd__or2_1 _08517_ (.A(\tms1x00.O_pla_ors[5][5] ),
    .B(_04090_),
    .X(_04097_));
 sky130_fd_sc_hd__o211a_1 _08518_ (.A1(net1042),
    .A2(net261),
    .B1(_04097_),
    .C1(net507),
    .X(_00913_));
 sky130_fd_sc_hd__mux2_1 _08519_ (.A0(net1034),
    .A1(\tms1x00.O_pla_ors[5][6] ),
    .S(net261),
    .X(_04098_));
 sky130_fd_sc_hd__or2_1 _08520_ (.A(net570),
    .B(_04098_),
    .X(_00914_));
 sky130_fd_sc_hd__or2_1 _08521_ (.A(\tms1x00.O_pla_ors[5][7] ),
    .B(_04090_),
    .X(_04099_));
 sky130_fd_sc_hd__o211a_1 _08522_ (.A1(net1027),
    .A2(net260),
    .B1(_04099_),
    .C1(net499),
    .X(_00915_));
 sky130_fd_sc_hd__mux2_1 _08523_ (.A0(net1020),
    .A1(\tms1x00.O_pla_ors[5][8] ),
    .S(net260),
    .X(_04100_));
 sky130_fd_sc_hd__or2_1 _08524_ (.A(net562),
    .B(_04100_),
    .X(_00916_));
 sky130_fd_sc_hd__or2_1 _08525_ (.A(\tms1x00.O_pla_ors[5][9] ),
    .B(_04090_),
    .X(_04101_));
 sky130_fd_sc_hd__o211a_1 _08526_ (.A1(net1011),
    .A2(net261),
    .B1(_04101_),
    .C1(net501),
    .X(_00917_));
 sky130_fd_sc_hd__mux2_1 _08527_ (.A0(net974),
    .A1(\tms1x00.O_pla_ors[5][10] ),
    .S(net261),
    .X(_04102_));
 sky130_fd_sc_hd__or2_1 _08528_ (.A(net571),
    .B(_04102_),
    .X(_00918_));
 sky130_fd_sc_hd__mux2_1 _08529_ (.A0(net970),
    .A1(\tms1x00.O_pla_ors[5][11] ),
    .S(net261),
    .X(_04103_));
 sky130_fd_sc_hd__or2_1 _08530_ (.A(net562),
    .B(_04103_),
    .X(_00919_));
 sky130_fd_sc_hd__mux2_1 _08531_ (.A0(net966),
    .A1(\tms1x00.O_pla_ors[5][12] ),
    .S(net260),
    .X(_04104_));
 sky130_fd_sc_hd__or2_1 _08532_ (.A(net556),
    .B(_04104_),
    .X(_00920_));
 sky130_fd_sc_hd__mux2_1 _08533_ (.A0(net961),
    .A1(\tms1x00.O_pla_ors[5][13] ),
    .S(net260),
    .X(_04105_));
 sky130_fd_sc_hd__or2_1 _08534_ (.A(net556),
    .B(_04105_),
    .X(_00921_));
 sky130_fd_sc_hd__mux2_1 _08535_ (.A0(net955),
    .A1(\tms1x00.O_pla_ors[5][14] ),
    .S(net260),
    .X(_04106_));
 sky130_fd_sc_hd__or2_1 _08536_ (.A(net568),
    .B(_04106_),
    .X(_00922_));
 sky130_fd_sc_hd__mux2_1 _08537_ (.A0(net949),
    .A1(\tms1x00.O_pla_ors[5][15] ),
    .S(net260),
    .X(_04107_));
 sky130_fd_sc_hd__or2_1 _08538_ (.A(net567),
    .B(_04107_),
    .X(_00923_));
 sky130_fd_sc_hd__or2_1 _08539_ (.A(\tms1x00.O_pla_ors[5][16] ),
    .B(_04090_),
    .X(_04108_));
 sky130_fd_sc_hd__o211a_1 _08540_ (.A1(net943),
    .A2(net261),
    .B1(_04108_),
    .C1(net502),
    .X(_00924_));
 sky130_fd_sc_hd__or2_1 _08541_ (.A(\tms1x00.O_pla_ors[5][17] ),
    .B(_04090_),
    .X(_04109_));
 sky130_fd_sc_hd__o211a_1 _08542_ (.A1(net941),
    .A2(net260),
    .B1(_04109_),
    .C1(net491),
    .X(_00925_));
 sky130_fd_sc_hd__or2_1 _08543_ (.A(\tms1x00.O_pla_ors[5][18] ),
    .B(_04090_),
    .X(_04110_));
 sky130_fd_sc_hd__o211a_1 _08544_ (.A1(net939),
    .A2(_04091_),
    .B1(_04110_),
    .C1(net507),
    .X(_00926_));
 sky130_fd_sc_hd__or2_1 _08545_ (.A(\tms1x00.O_pla_ors[5][19] ),
    .B(_04090_),
    .X(_04111_));
 sky130_fd_sc_hd__o211a_1 _08546_ (.A1(net936),
    .A2(net261),
    .B1(_04111_),
    .C1(net502),
    .X(_00927_));
 sky130_fd_sc_hd__o22a_1 _08547_ (.A1(\tms1x00.ins_pla_ands[27][0] ),
    .A2(_03593_),
    .B1(net218),
    .B2(_03456_),
    .X(_00928_));
 sky130_fd_sc_hd__o22a_1 _08548_ (.A1(\tms1x00.ins_pla_ands[27][1] ),
    .A2(net318),
    .B1(net219),
    .B2(net397),
    .X(_00929_));
 sky130_fd_sc_hd__o22a_1 _08549_ (.A1(\tms1x00.ins_pla_ands[27][2] ),
    .A2(net318),
    .B1(net218),
    .B2(_03428_),
    .X(_00930_));
 sky130_fd_sc_hd__o22a_1 _08550_ (.A1(\tms1x00.ins_pla_ands[27][3] ),
    .A2(net318),
    .B1(net218),
    .B2(_03430_),
    .X(_00931_));
 sky130_fd_sc_hd__o22a_1 _08551_ (.A1(\tms1x00.ins_pla_ands[27][4] ),
    .A2(net318),
    .B1(net218),
    .B2(_03478_),
    .X(_00932_));
 sky130_fd_sc_hd__o22a_1 _08552_ (.A1(\tms1x00.ins_pla_ands[27][5] ),
    .A2(net318),
    .B1(net218),
    .B2(net366),
    .X(_00933_));
 sky130_fd_sc_hd__o22a_1 _08553_ (.A1(\tms1x00.ins_pla_ands[27][6] ),
    .A2(net318),
    .B1(net218),
    .B2(_03434_),
    .X(_00934_));
 sky130_fd_sc_hd__o22a_1 _08554_ (.A1(\tms1x00.ins_pla_ands[27][7] ),
    .A2(net318),
    .B1(net218),
    .B2(net367),
    .X(_00935_));
 sky130_fd_sc_hd__o22a_1 _08555_ (.A1(\tms1x00.ins_pla_ands[27][9] ),
    .A2(net318),
    .B1(net219),
    .B2(net365),
    .X(_00936_));
 sky130_fd_sc_hd__o22a_1 _08556_ (.A1(\tms1x00.ins_pla_ands[27][10] ),
    .A2(net318),
    .B1(net218),
    .B2(_03459_),
    .X(_00937_));
 sky130_fd_sc_hd__o22a_1 _08557_ (.A1(\tms1x00.ins_pla_ands[27][12] ),
    .A2(_03593_),
    .B1(net219),
    .B2(_03484_),
    .X(_00938_));
 sky130_fd_sc_hd__mux2_1 _08558_ (.A0(\tms1x00.ins_pla_ands[27][15] ),
    .A1(net944),
    .S(net318),
    .X(_04112_));
 sky130_fd_sc_hd__and2_1 _08559_ (.A(net460),
    .B(_04112_),
    .X(_00939_));
 sky130_fd_sc_hd__and3_2 _08560_ (.A(net766),
    .B(net598),
    .C(net350),
    .X(_04113_));
 sky130_fd_sc_hd__mux2_1 _08561_ (.A0(\tms1x00.ins_pla_ands[17][0] ),
    .A1(net979),
    .S(net259),
    .X(_04114_));
 sky130_fd_sc_hd__or2_1 _08562_ (.A(net524),
    .B(_04114_),
    .X(_00940_));
 sky130_fd_sc_hd__nor2_2 _08563_ (.A(net516),
    .B(net259),
    .Y(_04115_));
 sky130_fd_sc_hd__or2_4 _08564_ (.A(net516),
    .B(net259),
    .X(_04116_));
 sky130_fd_sc_hd__o22a_1 _08565_ (.A1(\tms1x00.ins_pla_ands[17][1] ),
    .A2(net259),
    .B1(_04115_),
    .B2(net397),
    .X(_00941_));
 sky130_fd_sc_hd__o22a_1 _08566_ (.A1(\tms1x00.ins_pla_ands[17][6] ),
    .A2(_04113_),
    .B1(_04115_),
    .B2(_03434_),
    .X(_00942_));
 sky130_fd_sc_hd__mux2_1 _08567_ (.A0(\tms1x00.ins_pla_ands[17][7] ),
    .A1(net1026),
    .S(_04113_),
    .X(_04117_));
 sky130_fd_sc_hd__or2_1 _08568_ (.A(net524),
    .B(_04117_),
    .X(_00943_));
 sky130_fd_sc_hd__mux2_1 _08569_ (.A0(\tms1x00.ins_pla_ands[17][8] ),
    .A1(net1018),
    .S(net259),
    .X(_04118_));
 sky130_fd_sc_hd__or2_1 _08570_ (.A(net515),
    .B(_04118_),
    .X(_00944_));
 sky130_fd_sc_hd__o22a_1 _08571_ (.A1(\tms1x00.ins_pla_ands[17][9] ),
    .A2(net259),
    .B1(_04115_),
    .B2(net364),
    .X(_00945_));
 sky130_fd_sc_hd__mux2_1 _08572_ (.A0(\tms1x00.ins_pla_ands[17][12] ),
    .A1(net964),
    .S(net259),
    .X(_04119_));
 sky130_fd_sc_hd__or2_1 _08573_ (.A(net516),
    .B(_04119_),
    .X(_00946_));
 sky130_fd_sc_hd__o22a_1 _08574_ (.A1(\tms1x00.ins_pla_ands[17][13] ),
    .A2(net259),
    .B1(_04115_),
    .B2(net363),
    .X(_00947_));
 sky130_fd_sc_hd__mux2_1 _08575_ (.A0(\tms1x00.ins_pla_ands[17][14] ),
    .A1(net952),
    .S(net259),
    .X(_04120_));
 sky130_fd_sc_hd__or2_1 _08576_ (.A(net515),
    .B(_04120_),
    .X(_00948_));
 sky130_fd_sc_hd__mux2_1 _08577_ (.A0(\tms1x00.ins_pla_ands[17][15] ),
    .A1(net946),
    .S(net259),
    .X(_04121_));
 sky130_fd_sc_hd__and2_1 _08578_ (.A(net459),
    .B(_04121_),
    .X(_00949_));
 sky130_fd_sc_hd__mux2_1 _08579_ (.A0(net1065),
    .A1(\tms1x00.ins_pla_ands[8][2] ),
    .S(_03735_),
    .X(_04122_));
 sky130_fd_sc_hd__or2_1 _08580_ (.A(net528),
    .B(_04122_),
    .X(_00950_));
 sky130_fd_sc_hd__or2_1 _08581_ (.A(\tms1x00.ins_pla_ands[8][3] ),
    .B(_03734_),
    .X(_04123_));
 sky130_fd_sc_hd__o211a_1 _08582_ (.A1(net1055),
    .A2(_03735_),
    .B1(_04123_),
    .C1(net467),
    .X(_00951_));
 sky130_fd_sc_hd__or2_1 _08583_ (.A(\tms1x00.ins_pla_ands[8][4] ),
    .B(_03734_),
    .X(_04124_));
 sky130_fd_sc_hd__o211a_1 _08584_ (.A1(net1047),
    .A2(_03735_),
    .B1(_04124_),
    .C1(net466),
    .X(_00952_));
 sky130_fd_sc_hd__mux2_1 _08585_ (.A0(net965),
    .A1(\tms1x00.ins_pla_ands[8][12] ),
    .S(_03735_),
    .X(_04125_));
 sky130_fd_sc_hd__or2_1 _08586_ (.A(net535),
    .B(_04125_),
    .X(_00953_));
 sky130_fd_sc_hd__or2_1 _08587_ (.A(\tms1x00.ins_pla_ands[8][13] ),
    .B(_03734_),
    .X(_04126_));
 sky130_fd_sc_hd__o211a_1 _08588_ (.A1(net959),
    .A2(_03735_),
    .B1(_04126_),
    .C1(net467),
    .X(_00954_));
 sky130_fd_sc_hd__mux2_1 _08589_ (.A0(net952),
    .A1(\tms1x00.ins_pla_ands[8][14] ),
    .S(_03735_),
    .X(_04127_));
 sky130_fd_sc_hd__or2_1 _08590_ (.A(net529),
    .B(_04127_),
    .X(_00955_));
 sky130_fd_sc_hd__or2_1 _08591_ (.A(\tms1x00.ins_pla_ands[8][15] ),
    .B(_03734_),
    .X(_04128_));
 sky130_fd_sc_hd__o211a_1 _08592_ (.A1(net947),
    .A2(_03735_),
    .B1(_04128_),
    .C1(net470),
    .X(_00956_));
 sky130_fd_sc_hd__nor2_8 _08593_ (.A(net816),
    .B(net341),
    .Y(_04129_));
 sky130_fd_sc_hd__or2_4 _08594_ (.A(net814),
    .B(net342),
    .X(_04130_));
 sky130_fd_sc_hd__mux2_1 _08595_ (.A0(net980),
    .A1(\tms1x00.O_pla_ors[4][0] ),
    .S(net258),
    .X(_04131_));
 sky130_fd_sc_hd__or2_1 _08596_ (.A(net574),
    .B(_04131_),
    .X(_00957_));
 sky130_fd_sc_hd__or2_1 _08597_ (.A(\tms1x00.O_pla_ors[4][1] ),
    .B(_04129_),
    .X(_04132_));
 sky130_fd_sc_hd__o211a_1 _08598_ (.A1(net932),
    .A2(net258),
    .B1(_04132_),
    .C1(net501),
    .X(_00958_));
 sky130_fd_sc_hd__mux2_1 _08599_ (.A0(net1067),
    .A1(\tms1x00.O_pla_ors[4][2] ),
    .S(net257),
    .X(_04133_));
 sky130_fd_sc_hd__or2_1 _08600_ (.A(net560),
    .B(_04133_),
    .X(_00959_));
 sky130_fd_sc_hd__mux2_1 _08601_ (.A0(net1060),
    .A1(\tms1x00.O_pla_ors[4][3] ),
    .S(net257),
    .X(_04134_));
 sky130_fd_sc_hd__or2_1 _08602_ (.A(net557),
    .B(_04134_),
    .X(_00960_));
 sky130_fd_sc_hd__or2_1 _08603_ (.A(\tms1x00.O_pla_ors[4][4] ),
    .B(_04129_),
    .X(_04135_));
 sky130_fd_sc_hd__o211a_1 _08604_ (.A1(net1050),
    .A2(net257),
    .B1(_04135_),
    .C1(net492),
    .X(_00961_));
 sky130_fd_sc_hd__mux2_1 _08605_ (.A0(net1043),
    .A1(\tms1x00.O_pla_ors[4][5] ),
    .S(net257),
    .X(_04136_));
 sky130_fd_sc_hd__or2_1 _08606_ (.A(net556),
    .B(_04136_),
    .X(_00962_));
 sky130_fd_sc_hd__mux2_1 _08607_ (.A0(net1034),
    .A1(\tms1x00.O_pla_ors[4][6] ),
    .S(net258),
    .X(_04137_));
 sky130_fd_sc_hd__or2_1 _08608_ (.A(net571),
    .B(_04137_),
    .X(_00963_));
 sky130_fd_sc_hd__or2_1 _08609_ (.A(\tms1x00.O_pla_ors[4][7] ),
    .B(_04129_),
    .X(_04138_));
 sky130_fd_sc_hd__o211a_1 _08610_ (.A1(net1027),
    .A2(net258),
    .B1(_04138_),
    .C1(net499),
    .X(_00964_));
 sky130_fd_sc_hd__mux2_1 _08611_ (.A0(net1019),
    .A1(\tms1x00.O_pla_ors[4][8] ),
    .S(net257),
    .X(_04139_));
 sky130_fd_sc_hd__or2_1 _08612_ (.A(net557),
    .B(_04139_),
    .X(_00965_));
 sky130_fd_sc_hd__mux2_1 _08613_ (.A0(net1011),
    .A1(\tms1x00.O_pla_ors[4][9] ),
    .S(net258),
    .X(_04140_));
 sky130_fd_sc_hd__or2_1 _08614_ (.A(net571),
    .B(_04140_),
    .X(_00966_));
 sky130_fd_sc_hd__or2_1 _08615_ (.A(\tms1x00.O_pla_ors[4][10] ),
    .B(_04129_),
    .X(_04141_));
 sky130_fd_sc_hd__o211a_1 _08616_ (.A1(net974),
    .A2(net258),
    .B1(_04141_),
    .C1(net501),
    .X(_00967_));
 sky130_fd_sc_hd__mux2_1 _08617_ (.A0(net970),
    .A1(\tms1x00.O_pla_ors[4][11] ),
    .S(net257),
    .X(_04142_));
 sky130_fd_sc_hd__or2_1 _08618_ (.A(net560),
    .B(_04142_),
    .X(_00968_));
 sky130_fd_sc_hd__mux2_1 _08619_ (.A0(net966),
    .A1(\tms1x00.O_pla_ors[4][12] ),
    .S(net257),
    .X(_04143_));
 sky130_fd_sc_hd__or2_1 _08620_ (.A(net557),
    .B(_04143_),
    .X(_00969_));
 sky130_fd_sc_hd__mux2_1 _08621_ (.A0(net962),
    .A1(\tms1x00.O_pla_ors[4][13] ),
    .S(net257),
    .X(_04144_));
 sky130_fd_sc_hd__or2_1 _08622_ (.A(net556),
    .B(_04144_),
    .X(_00970_));
 sky130_fd_sc_hd__mux2_1 _08623_ (.A0(net956),
    .A1(\tms1x00.O_pla_ors[4][14] ),
    .S(net258),
    .X(_04145_));
 sky130_fd_sc_hd__or2_1 _08624_ (.A(net569),
    .B(_04145_),
    .X(_00971_));
 sky130_fd_sc_hd__or2_1 _08625_ (.A(\tms1x00.O_pla_ors[4][15] ),
    .B(_04129_),
    .X(_04146_));
 sky130_fd_sc_hd__o211a_1 _08626_ (.A1(net949),
    .A2(net258),
    .B1(_04146_),
    .C1(net499),
    .X(_00972_));
 sky130_fd_sc_hd__or2_1 _08627_ (.A(\tms1x00.O_pla_ors[4][16] ),
    .B(_04129_),
    .X(_04147_));
 sky130_fd_sc_hd__o211a_1 _08628_ (.A1(net943),
    .A2(net258),
    .B1(_04147_),
    .C1(net502),
    .X(_00973_));
 sky130_fd_sc_hd__or2_1 _08629_ (.A(\tms1x00.O_pla_ors[4][17] ),
    .B(_04129_),
    .X(_04148_));
 sky130_fd_sc_hd__o211a_1 _08630_ (.A1(net941),
    .A2(net257),
    .B1(_04148_),
    .C1(net491),
    .X(_00974_));
 sky130_fd_sc_hd__or2_1 _08631_ (.A(\tms1x00.O_pla_ors[4][18] ),
    .B(_04129_),
    .X(_04149_));
 sky130_fd_sc_hd__o211a_1 _08632_ (.A1(net939),
    .A2(net258),
    .B1(_04149_),
    .C1(net503),
    .X(_00975_));
 sky130_fd_sc_hd__or2_1 _08633_ (.A(\tms1x00.O_pla_ors[4][19] ),
    .B(_04129_),
    .X(_04150_));
 sky130_fd_sc_hd__o211a_1 _08634_ (.A1(net937),
    .A2(net257),
    .B1(_04150_),
    .C1(net491),
    .X(_00976_));
 sky130_fd_sc_hd__a31o_1 _08635_ (.A1(\tms1x00.ins_pla_ands[12][1] ),
    .A2(net369),
    .A3(net274),
    .B1(net392),
    .X(_04151_));
 sky130_fd_sc_hd__a21o_1 _08636_ (.A1(net397),
    .A2(_03922_),
    .B1(_04151_),
    .X(_00977_));
 sky130_fd_sc_hd__or3_1 _08637_ (.A(\tms1x00.ins_pla_ands[12][6] ),
    .B(net377),
    .C(_03922_),
    .X(_04152_));
 sky130_fd_sc_hd__o211a_1 _08638_ (.A1(_03909_),
    .A2(net275),
    .B1(_04152_),
    .C1(net383),
    .X(_00978_));
 sky130_fd_sc_hd__a31o_1 _08639_ (.A1(\tms1x00.ins_pla_ands[12][7] ),
    .A2(net369),
    .A3(net275),
    .B1(net392),
    .X(_04153_));
 sky130_fd_sc_hd__a21o_1 _08640_ (.A1(net368),
    .A2(_03922_),
    .B1(_04153_),
    .X(_00979_));
 sky130_fd_sc_hd__o22a_1 _08641_ (.A1(\tms1x00.ins_pla_ands[26][1] ),
    .A2(_03473_),
    .B1(_03474_),
    .B2(net397),
    .X(_00980_));
 sky130_fd_sc_hd__o22a_1 _08642_ (.A1(\tms1x00.ins_pla_ands[26][3] ),
    .A2(_03473_),
    .B1(_03474_),
    .B2(_03430_),
    .X(_00981_));
 sky130_fd_sc_hd__o22a_1 _08643_ (.A1(\tms1x00.ins_pla_ands[26][5] ),
    .A2(_03473_),
    .B1(_03474_),
    .B2(net366),
    .X(_00982_));
 sky130_fd_sc_hd__o22a_1 _08644_ (.A1(\tms1x00.ins_pla_ands[26][7] ),
    .A2(_03473_),
    .B1(_03474_),
    .B2(net367),
    .X(_00983_));
 sky130_fd_sc_hd__mux2_1 _08645_ (.A0(\tms1x00.ins_pla_ands[26][14] ),
    .A1(net951),
    .S(_03473_),
    .X(_04154_));
 sky130_fd_sc_hd__or2_1 _08646_ (.A(net518),
    .B(_04154_),
    .X(_00984_));
 sky130_fd_sc_hd__or4_2 _08647_ (.A(net945),
    .B(net714),
    .C(net348),
    .D(net710),
    .X(_04155_));
 sky130_fd_sc_hd__o211a_1 _08648_ (.A1(\tms1x00.ins_pla_ands[26][15] ),
    .A2(_03473_),
    .B1(_04155_),
    .C1(net460),
    .X(_00985_));
 sky130_fd_sc_hd__and3_4 _08649_ (.A(net847),
    .B(net598),
    .C(net351),
    .X(_04156_));
 sky130_fd_sc_hd__or3_2 _08650_ (.A(net825),
    .B(_03353_),
    .C(net348),
    .X(_04157_));
 sky130_fd_sc_hd__or3_1 _08651_ (.A(\tms1x00.ins_pla_ands[16][0] ),
    .B(net376),
    .C(_04156_),
    .X(_04158_));
 sky130_fd_sc_hd__o211a_1 _08652_ (.A1(_03574_),
    .A2(net255),
    .B1(_04158_),
    .C1(net383),
    .X(_00986_));
 sky130_fd_sc_hd__a31o_1 _08653_ (.A1(\tms1x00.ins_pla_ands[16][1] ),
    .A2(net369),
    .A3(net255),
    .B1(net391),
    .X(_04159_));
 sky130_fd_sc_hd__a21o_1 _08654_ (.A1(net397),
    .A2(_04156_),
    .B1(_04159_),
    .X(_00987_));
 sky130_fd_sc_hd__or3_1 _08655_ (.A(\tms1x00.ins_pla_ands[16][6] ),
    .B(net376),
    .C(_04156_),
    .X(_04160_));
 sky130_fd_sc_hd__o211a_1 _08656_ (.A1(_03909_),
    .A2(net256),
    .B1(_04160_),
    .C1(net383),
    .X(_00988_));
 sky130_fd_sc_hd__a31o_1 _08657_ (.A1(\tms1x00.ins_pla_ands[16][7] ),
    .A2(net369),
    .A3(net256),
    .B1(net391),
    .X(_04161_));
 sky130_fd_sc_hd__a21o_1 _08658_ (.A1(net368),
    .A2(_04156_),
    .B1(_04161_),
    .X(_00989_));
 sky130_fd_sc_hd__mux2_1 _08659_ (.A0(\tms1x00.ins_pla_ands[7][12] ),
    .A1(net965),
    .S(_03727_),
    .X(_04162_));
 sky130_fd_sc_hd__or2_1 _08660_ (.A(net535),
    .B(_04162_),
    .X(_00990_));
 sky130_fd_sc_hd__or4_1 _08661_ (.A(net960),
    .B(net781),
    .C(net348),
    .D(net707),
    .X(_04163_));
 sky130_fd_sc_hd__o211a_1 _08662_ (.A1(\tms1x00.ins_pla_ands[7][13] ),
    .A2(_03727_),
    .B1(_04163_),
    .C1(net470),
    .X(_00991_));
 sky130_fd_sc_hd__mux2_1 _08663_ (.A0(\tms1x00.ins_pla_ands[7][14] ),
    .A1(net954),
    .S(_03727_),
    .X(_04164_));
 sky130_fd_sc_hd__or2_1 _08664_ (.A(net534),
    .B(_04164_),
    .X(_00992_));
 sky130_fd_sc_hd__or4_1 _08665_ (.A(net947),
    .B(net781),
    .C(net349),
    .D(net707),
    .X(_04165_));
 sky130_fd_sc_hd__o211a_1 _08666_ (.A1(\tms1x00.ins_pla_ands[7][15] ),
    .A2(_03727_),
    .B1(_04165_),
    .C1(net471),
    .X(_00993_));
 sky130_fd_sc_hd__nor2_4 _08667_ (.A(net871),
    .B(net341),
    .Y(_04166_));
 sky130_fd_sc_hd__or2_4 _08668_ (.A(net871),
    .B(net342),
    .X(_04167_));
 sky130_fd_sc_hd__mux2_1 _08669_ (.A0(net983),
    .A1(\tms1x00.O_pla_ors[3][0] ),
    .S(net254),
    .X(_04168_));
 sky130_fd_sc_hd__or2_1 _08670_ (.A(net573),
    .B(_04168_),
    .X(_00994_));
 sky130_fd_sc_hd__mux2_1 _08671_ (.A0(net932),
    .A1(\tms1x00.O_pla_ors[3][1] ),
    .S(net254),
    .X(_04169_));
 sky130_fd_sc_hd__or2_1 _08672_ (.A(net574),
    .B(_04169_),
    .X(_00995_));
 sky130_fd_sc_hd__or2_1 _08673_ (.A(\tms1x00.O_pla_ors[3][2] ),
    .B(_04166_),
    .X(_04170_));
 sky130_fd_sc_hd__o211a_1 _08674_ (.A1(net1068),
    .A2(net253),
    .B1(_04170_),
    .C1(net498),
    .X(_00996_));
 sky130_fd_sc_hd__mux2_1 _08675_ (.A0(net1059),
    .A1(\tms1x00.O_pla_ors[3][3] ),
    .S(net253),
    .X(_04171_));
 sky130_fd_sc_hd__or2_1 _08676_ (.A(net556),
    .B(_04171_),
    .X(_00997_));
 sky130_fd_sc_hd__mux2_1 _08677_ (.A0(net1050),
    .A1(\tms1x00.O_pla_ors[3][4] ),
    .S(net253),
    .X(_04172_));
 sky130_fd_sc_hd__or2_1 _08678_ (.A(net561),
    .B(_04172_),
    .X(_00998_));
 sky130_fd_sc_hd__mux2_1 _08679_ (.A0(net1044),
    .A1(\tms1x00.O_pla_ors[3][5] ),
    .S(net253),
    .X(_04173_));
 sky130_fd_sc_hd__or2_1 _08680_ (.A(net569),
    .B(_04173_),
    .X(_00999_));
 sky130_fd_sc_hd__mux2_1 _08681_ (.A0(net1035),
    .A1(\tms1x00.O_pla_ors[3][6] ),
    .S(net254),
    .X(_04174_));
 sky130_fd_sc_hd__or2_1 _08682_ (.A(net571),
    .B(_04174_),
    .X(_01000_));
 sky130_fd_sc_hd__mux2_1 _08683_ (.A0(net1027),
    .A1(\tms1x00.O_pla_ors[3][7] ),
    .S(_04167_),
    .X(_04175_));
 sky130_fd_sc_hd__or2_1 _08684_ (.A(net567),
    .B(_04175_),
    .X(_01001_));
 sky130_fd_sc_hd__mux2_1 _08685_ (.A0(net1020),
    .A1(\tms1x00.O_pla_ors[3][8] ),
    .S(net253),
    .X(_04176_));
 sky130_fd_sc_hd__or2_1 _08686_ (.A(net561),
    .B(_04176_),
    .X(_01002_));
 sky130_fd_sc_hd__mux2_1 _08687_ (.A0(net1011),
    .A1(\tms1x00.O_pla_ors[3][9] ),
    .S(net254),
    .X(_04177_));
 sky130_fd_sc_hd__or2_1 _08688_ (.A(net570),
    .B(_04177_),
    .X(_01003_));
 sky130_fd_sc_hd__mux2_1 _08689_ (.A0(net974),
    .A1(\tms1x00.O_pla_ors[3][10] ),
    .S(net254),
    .X(_04178_));
 sky130_fd_sc_hd__or2_1 _08690_ (.A(net570),
    .B(_04178_),
    .X(_01004_));
 sky130_fd_sc_hd__mux2_1 _08691_ (.A0(net970),
    .A1(\tms1x00.O_pla_ors[3][11] ),
    .S(net253),
    .X(_04179_));
 sky130_fd_sc_hd__or2_1 _08692_ (.A(net561),
    .B(_04179_),
    .X(_01005_));
 sky130_fd_sc_hd__or2_1 _08693_ (.A(\tms1x00.O_pla_ors[3][12] ),
    .B(_04166_),
    .X(_04180_));
 sky130_fd_sc_hd__o211a_1 _08694_ (.A1(net967),
    .A2(net253),
    .B1(_04180_),
    .C1(net492),
    .X(_01006_));
 sky130_fd_sc_hd__mux2_1 _08695_ (.A0(net961),
    .A1(\tms1x00.O_pla_ors[3][13] ),
    .S(net253),
    .X(_04181_));
 sky130_fd_sc_hd__or2_1 _08696_ (.A(net566),
    .B(_04181_),
    .X(_01007_));
 sky130_fd_sc_hd__or2_1 _08697_ (.A(\tms1x00.O_pla_ors[3][14] ),
    .B(_04166_),
    .X(_04182_));
 sky130_fd_sc_hd__o211a_1 _08698_ (.A1(net956),
    .A2(net254),
    .B1(_04182_),
    .C1(net499),
    .X(_01008_));
 sky130_fd_sc_hd__or2_1 _08699_ (.A(\tms1x00.O_pla_ors[3][15] ),
    .B(_04166_),
    .X(_04183_));
 sky130_fd_sc_hd__o211a_1 _08700_ (.A1(net949),
    .A2(net253),
    .B1(_04183_),
    .C1(net499),
    .X(_01009_));
 sky130_fd_sc_hd__or2_1 _08701_ (.A(\tms1x00.O_pla_ors[3][16] ),
    .B(_04166_),
    .X(_04184_));
 sky130_fd_sc_hd__o211a_1 _08702_ (.A1(net943),
    .A2(net254),
    .B1(_04184_),
    .C1(net499),
    .X(_01010_));
 sky130_fd_sc_hd__or2_1 _08703_ (.A(\tms1x00.O_pla_ors[3][17] ),
    .B(_04166_),
    .X(_04185_));
 sky130_fd_sc_hd__o211a_1 _08704_ (.A1(net941),
    .A2(net253),
    .B1(_04185_),
    .C1(net491),
    .X(_01011_));
 sky130_fd_sc_hd__or2_1 _08705_ (.A(\tms1x00.O_pla_ors[3][18] ),
    .B(_04166_),
    .X(_04186_));
 sky130_fd_sc_hd__o211a_1 _08706_ (.A1(net939),
    .A2(net254),
    .B1(_04186_),
    .C1(net503),
    .X(_01012_));
 sky130_fd_sc_hd__mux2_1 _08707_ (.A0(net936),
    .A1(\tms1x00.O_pla_ors[3][19] ),
    .S(net254),
    .X(_04187_));
 sky130_fd_sc_hd__or2_1 _08708_ (.A(net570),
    .B(_04187_),
    .X(_01013_));
 sky130_fd_sc_hd__mux2_1 _08709_ (.A0(\tms1x00.ins_pla_ands[25][2] ),
    .A1(net1066),
    .S(net290),
    .X(_04188_));
 sky130_fd_sc_hd__or2_1 _08710_ (.A(net511),
    .B(_04188_),
    .X(_01014_));
 sky130_fd_sc_hd__o22a_1 _08711_ (.A1(\tms1x00.ins_pla_ands[25][3] ),
    .A2(_03793_),
    .B1(_03794_),
    .B2(_03430_),
    .X(_01015_));
 sky130_fd_sc_hd__mux2_1 _08712_ (.A0(\tms1x00.ins_pla_ands[25][4] ),
    .A1(net1049),
    .S(net290),
    .X(_04189_));
 sky130_fd_sc_hd__or2_1 _08713_ (.A(net512),
    .B(_04189_),
    .X(_01016_));
 sky130_fd_sc_hd__o22a_1 _08714_ (.A1(\tms1x00.ins_pla_ands[25][5] ),
    .A2(_03793_),
    .B1(_03794_),
    .B2(net366),
    .X(_01017_));
 sky130_fd_sc_hd__mux2_1 _08715_ (.A0(\tms1x00.ins_pla_ands[25][6] ),
    .A1(net1033),
    .S(net290),
    .X(_04190_));
 sky130_fd_sc_hd__or2_1 _08716_ (.A(net511),
    .B(_04190_),
    .X(_01018_));
 sky130_fd_sc_hd__o22a_1 _08717_ (.A1(\tms1x00.ins_pla_ands[25][7] ),
    .A2(net290),
    .B1(_03794_),
    .B2(net367),
    .X(_01019_));
 sky130_fd_sc_hd__mux2_1 _08718_ (.A0(\tms1x00.ins_pla_ands[25][8] ),
    .A1(net1014),
    .S(_03793_),
    .X(_04191_));
 sky130_fd_sc_hd__or2_1 _08719_ (.A(net511),
    .B(_04191_),
    .X(_01020_));
 sky130_fd_sc_hd__o22a_1 _08720_ (.A1(\tms1x00.ins_pla_ands[25][9] ),
    .A2(net290),
    .B1(_03794_),
    .B2(net364),
    .X(_01021_));
 sky130_fd_sc_hd__mux2_1 _08721_ (.A0(\tms1x00.ins_pla_ands[25][12] ),
    .A1(net963),
    .S(net290),
    .X(_04192_));
 sky130_fd_sc_hd__or2_1 _08722_ (.A(net511),
    .B(_04192_),
    .X(_01022_));
 sky130_fd_sc_hd__o22a_1 _08723_ (.A1(\tms1x00.ins_pla_ands[25][13] ),
    .A2(net290),
    .B1(_03794_),
    .B2(net363),
    .X(_01023_));
 sky130_fd_sc_hd__mux2_1 _08724_ (.A0(\tms1x00.ins_pla_ands[25][14] ),
    .A1(net951),
    .S(net290),
    .X(_04193_));
 sky130_fd_sc_hd__or2_1 _08725_ (.A(net511),
    .B(_04193_),
    .X(_01024_));
 sky130_fd_sc_hd__mux2_1 _08726_ (.A0(\tms1x00.ins_pla_ands[25][15] ),
    .A1(net944),
    .S(net290),
    .X(_04194_));
 sky130_fd_sc_hd__and2_1 _08727_ (.A(net460),
    .B(_04194_),
    .X(_01025_));
 sky130_fd_sc_hd__mux2_1 _08728_ (.A0(net1066),
    .A1(\tms1x00.ins_pla_ands[16][2] ),
    .S(net256),
    .X(_04195_));
 sky130_fd_sc_hd__or2_1 _08729_ (.A(net516),
    .B(_04195_),
    .X(_01026_));
 sky130_fd_sc_hd__or2_1 _08730_ (.A(\tms1x00.ins_pla_ands[16][3] ),
    .B(_04156_),
    .X(_04196_));
 sky130_fd_sc_hd__o211a_1 _08731_ (.A1(net1058),
    .A2(net255),
    .B1(_04196_),
    .C1(net460),
    .X(_01027_));
 sky130_fd_sc_hd__mux2_1 _08732_ (.A0(net1049),
    .A1(\tms1x00.ins_pla_ands[16][4] ),
    .S(net256),
    .X(_04197_));
 sky130_fd_sc_hd__or2_1 _08733_ (.A(net524),
    .B(_04197_),
    .X(_01028_));
 sky130_fd_sc_hd__or2_1 _08734_ (.A(\tms1x00.ins_pla_ands[16][5] ),
    .B(_04156_),
    .X(_04198_));
 sky130_fd_sc_hd__o211a_1 _08735_ (.A1(net1041),
    .A2(net256),
    .B1(_04198_),
    .C1(net462),
    .X(_01029_));
 sky130_fd_sc_hd__mux2_1 _08736_ (.A0(net1018),
    .A1(\tms1x00.ins_pla_ands[16][8] ),
    .S(net255),
    .X(_04199_));
 sky130_fd_sc_hd__or2_1 _08737_ (.A(net515),
    .B(_04199_),
    .X(_01030_));
 sky130_fd_sc_hd__or2_1 _08738_ (.A(\tms1x00.ins_pla_ands[16][9] ),
    .B(_04156_),
    .X(_04200_));
 sky130_fd_sc_hd__o211a_1 _08739_ (.A1(net1010),
    .A2(net255),
    .B1(_04200_),
    .C1(net459),
    .X(_01031_));
 sky130_fd_sc_hd__or2_1 _08740_ (.A(\tms1x00.ins_pla_ands[16][10] ),
    .B(_04156_),
    .X(_04201_));
 sky130_fd_sc_hd__o211a_1 _08741_ (.A1(net973),
    .A2(net255),
    .B1(_04201_),
    .C1(net460),
    .X(_01032_));
 sky130_fd_sc_hd__mux2_1 _08742_ (.A0(net969),
    .A1(\tms1x00.ins_pla_ands[16][11] ),
    .S(net256),
    .X(_04202_));
 sky130_fd_sc_hd__or2_1 _08743_ (.A(net516),
    .B(_04202_),
    .X(_01033_));
 sky130_fd_sc_hd__mux2_1 _08744_ (.A0(net964),
    .A1(\tms1x00.ins_pla_ands[16][12] ),
    .S(net255),
    .X(_04203_));
 sky130_fd_sc_hd__or2_1 _08745_ (.A(net516),
    .B(_04203_),
    .X(_01034_));
 sky130_fd_sc_hd__or2_1 _08746_ (.A(\tms1x00.ins_pla_ands[16][13] ),
    .B(_04156_),
    .X(_04204_));
 sky130_fd_sc_hd__o211a_1 _08747_ (.A1(net959),
    .A2(net255),
    .B1(_04204_),
    .C1(net459),
    .X(_01035_));
 sky130_fd_sc_hd__mux2_1 _08748_ (.A0(net952),
    .A1(\tms1x00.ins_pla_ands[16][14] ),
    .S(net255),
    .X(_04205_));
 sky130_fd_sc_hd__or2_1 _08749_ (.A(net515),
    .B(_04205_),
    .X(_01036_));
 sky130_fd_sc_hd__or2_1 _08750_ (.A(\tms1x00.ins_pla_ands[16][15] ),
    .B(_04156_),
    .X(_04206_));
 sky130_fd_sc_hd__o211a_1 _08751_ (.A1(net946),
    .A2(net255),
    .B1(_04206_),
    .C1(net459),
    .X(_01037_));
 sky130_fd_sc_hd__or2_1 _08752_ (.A(\tms1x00.ins_pla_ands[6][2] ),
    .B(_03570_),
    .X(_04207_));
 sky130_fd_sc_hd__o211a_1 _08753_ (.A1(net1066),
    .A2(_03571_),
    .B1(_04207_),
    .C1(net469),
    .X(_01038_));
 sky130_fd_sc_hd__mux2_1 _08754_ (.A0(net1056),
    .A1(\tms1x00.ins_pla_ands[6][3] ),
    .S(_03571_),
    .X(_04208_));
 sky130_fd_sc_hd__or2_1 _08755_ (.A(net535),
    .B(_04208_),
    .X(_01039_));
 sky130_fd_sc_hd__mux2_1 _08756_ (.A0(net965),
    .A1(\tms1x00.ins_pla_ands[6][12] ),
    .S(_03571_),
    .X(_04209_));
 sky130_fd_sc_hd__or2_1 _08757_ (.A(net535),
    .B(_04209_),
    .X(_01040_));
 sky130_fd_sc_hd__or2_1 _08758_ (.A(\tms1x00.ins_pla_ands[6][13] ),
    .B(_03570_),
    .X(_04210_));
 sky130_fd_sc_hd__o211a_1 _08759_ (.A1(net960),
    .A2(_03571_),
    .B1(_04210_),
    .C1(net475),
    .X(_01041_));
 sky130_fd_sc_hd__mux2_1 _08760_ (.A0(net954),
    .A1(\tms1x00.ins_pla_ands[6][14] ),
    .S(_03571_),
    .X(_04211_));
 sky130_fd_sc_hd__or2_1 _08761_ (.A(net531),
    .B(_04211_),
    .X(_01042_));
 sky130_fd_sc_hd__or2_1 _08762_ (.A(\tms1x00.ins_pla_ands[6][15] ),
    .B(_03570_),
    .X(_04212_));
 sky130_fd_sc_hd__o211a_1 _08763_ (.A1(net947),
    .A2(_03571_),
    .B1(_04212_),
    .C1(net475),
    .X(_01043_));
 sky130_fd_sc_hd__nor2_8 _08764_ (.A(net737),
    .B(net341),
    .Y(_04213_));
 sky130_fd_sc_hd__or2_4 _08765_ (.A(net737),
    .B(net341),
    .X(_04214_));
 sky130_fd_sc_hd__mux2_1 _08766_ (.A0(net980),
    .A1(\tms1x00.O_pla_ors[2][0] ),
    .S(net252),
    .X(_04215_));
 sky130_fd_sc_hd__or2_1 _08767_ (.A(net576),
    .B(_04215_),
    .X(_01044_));
 sky130_fd_sc_hd__mux2_1 _08768_ (.A0(net931),
    .A1(\tms1x00.O_pla_ors[2][1] ),
    .S(net252),
    .X(_04216_));
 sky130_fd_sc_hd__or2_1 _08769_ (.A(net576),
    .B(_04216_),
    .X(_01045_));
 sky130_fd_sc_hd__mux2_1 _08770_ (.A0(net1067),
    .A1(\tms1x00.O_pla_ors[2][2] ),
    .S(net251),
    .X(_04217_));
 sky130_fd_sc_hd__or2_1 _08771_ (.A(net561),
    .B(_04217_),
    .X(_01046_));
 sky130_fd_sc_hd__mux2_1 _08772_ (.A0(net1060),
    .A1(\tms1x00.O_pla_ors[2][3] ),
    .S(net251),
    .X(_04218_));
 sky130_fd_sc_hd__or2_1 _08773_ (.A(net566),
    .B(_04218_),
    .X(_01047_));
 sky130_fd_sc_hd__mux2_1 _08774_ (.A0(net1050),
    .A1(\tms1x00.O_pla_ors[2][4] ),
    .S(net251),
    .X(_04219_));
 sky130_fd_sc_hd__or2_1 _08775_ (.A(net556),
    .B(_04219_),
    .X(_01048_));
 sky130_fd_sc_hd__or2_1 _08776_ (.A(\tms1x00.O_pla_ors[2][5] ),
    .B(_04213_),
    .X(_04220_));
 sky130_fd_sc_hd__o211a_1 _08777_ (.A1(net1042),
    .A2(net252),
    .B1(_04220_),
    .C1(net507),
    .X(_01049_));
 sky130_fd_sc_hd__or2_1 _08778_ (.A(\tms1x00.O_pla_ors[2][6] ),
    .B(_04213_),
    .X(_04221_));
 sky130_fd_sc_hd__o211a_1 _08779_ (.A1(net1035),
    .A2(net252),
    .B1(_04221_),
    .C1(net501),
    .X(_01050_));
 sky130_fd_sc_hd__mux2_1 _08780_ (.A0(net1027),
    .A1(\tms1x00.O_pla_ors[2][7] ),
    .S(net252),
    .X(_04222_));
 sky130_fd_sc_hd__or2_1 _08781_ (.A(net572),
    .B(_04222_),
    .X(_01051_));
 sky130_fd_sc_hd__mux2_1 _08782_ (.A0(net1020),
    .A1(\tms1x00.O_pla_ors[2][8] ),
    .S(net251),
    .X(_04223_));
 sky130_fd_sc_hd__or2_1 _08783_ (.A(net562),
    .B(_04223_),
    .X(_01052_));
 sky130_fd_sc_hd__mux2_1 _08784_ (.A0(net1011),
    .A1(\tms1x00.O_pla_ors[2][9] ),
    .S(net252),
    .X(_04224_));
 sky130_fd_sc_hd__or2_1 _08785_ (.A(net570),
    .B(_04224_),
    .X(_01053_));
 sky130_fd_sc_hd__mux2_1 _08786_ (.A0(net974),
    .A1(\tms1x00.O_pla_ors[2][10] ),
    .S(net252),
    .X(_04225_));
 sky130_fd_sc_hd__or2_1 _08787_ (.A(net570),
    .B(_04225_),
    .X(_01054_));
 sky130_fd_sc_hd__or2_1 _08788_ (.A(\tms1x00.O_pla_ors[2][11] ),
    .B(_04213_),
    .X(_04226_));
 sky130_fd_sc_hd__o211a_1 _08789_ (.A1(net970),
    .A2(net251),
    .B1(_04226_),
    .C1(net498),
    .X(_01055_));
 sky130_fd_sc_hd__or2_1 _08790_ (.A(\tms1x00.O_pla_ors[2][12] ),
    .B(_04213_),
    .X(_04227_));
 sky130_fd_sc_hd__o211a_1 _08791_ (.A1(net967),
    .A2(net251),
    .B1(_04227_),
    .C1(net492),
    .X(_01056_));
 sky130_fd_sc_hd__mux2_1 _08792_ (.A0(net961),
    .A1(\tms1x00.O_pla_ors[2][13] ),
    .S(net251),
    .X(_04228_));
 sky130_fd_sc_hd__or2_1 _08793_ (.A(net556),
    .B(_04228_),
    .X(_01057_));
 sky130_fd_sc_hd__or2_1 _08794_ (.A(\tms1x00.O_pla_ors[2][14] ),
    .B(_04213_),
    .X(_04229_));
 sky130_fd_sc_hd__o211a_1 _08795_ (.A1(net956),
    .A2(net251),
    .B1(_04229_),
    .C1(net499),
    .X(_01058_));
 sky130_fd_sc_hd__or2_1 _08796_ (.A(\tms1x00.O_pla_ors[2][15] ),
    .B(_04213_),
    .X(_04230_));
 sky130_fd_sc_hd__o211a_1 _08797_ (.A1(net949),
    .A2(net251),
    .B1(_04230_),
    .C1(net499),
    .X(_01059_));
 sky130_fd_sc_hd__or2_1 _08798_ (.A(\tms1x00.O_pla_ors[2][16] ),
    .B(_04213_),
    .X(_04231_));
 sky130_fd_sc_hd__o211a_1 _08799_ (.A1(net943),
    .A2(net252),
    .B1(_04231_),
    .C1(net502),
    .X(_01060_));
 sky130_fd_sc_hd__or2_1 _08800_ (.A(\tms1x00.O_pla_ors[2][17] ),
    .B(_04213_),
    .X(_04232_));
 sky130_fd_sc_hd__o211a_1 _08801_ (.A1(net941),
    .A2(net251),
    .B1(_04232_),
    .C1(net491),
    .X(_01061_));
 sky130_fd_sc_hd__mux2_1 _08802_ (.A0(net939),
    .A1(\tms1x00.O_pla_ors[2][18] ),
    .S(net252),
    .X(_04233_));
 sky130_fd_sc_hd__or2_1 _08803_ (.A(net576),
    .B(_04233_),
    .X(_01062_));
 sky130_fd_sc_hd__or2_1 _08804_ (.A(\tms1x00.O_pla_ors[2][19] ),
    .B(_04213_),
    .X(_04234_));
 sky130_fd_sc_hd__o211a_1 _08805_ (.A1(net936),
    .A2(net252),
    .B1(_04234_),
    .C1(net501),
    .X(_01063_));
 sky130_fd_sc_hd__mux2_1 _08806_ (.A0(\tms1x00.ins_pla_ands[24][4] ),
    .A1(net1049),
    .S(net299),
    .X(_04235_));
 sky130_fd_sc_hd__or2_1 _08807_ (.A(net512),
    .B(_04235_),
    .X(_01064_));
 sky130_fd_sc_hd__o22a_1 _08808_ (.A1(\tms1x00.ins_pla_ands[24][5] ),
    .A2(net299),
    .B1(_03717_),
    .B2(net366),
    .X(_01065_));
 sky130_fd_sc_hd__mux2_1 _08809_ (.A0(\tms1x00.ins_pla_ands[24][6] ),
    .A1(net1033),
    .S(net299),
    .X(_04236_));
 sky130_fd_sc_hd__or2_1 _08810_ (.A(net511),
    .B(_04236_),
    .X(_01066_));
 sky130_fd_sc_hd__o22a_1 _08811_ (.A1(\tms1x00.ins_pla_ands[24][7] ),
    .A2(_03716_),
    .B1(_03717_),
    .B2(net367),
    .X(_01067_));
 sky130_fd_sc_hd__mux2_1 _08812_ (.A0(\tms1x00.ins_pla_ands[24][8] ),
    .A1(net1014),
    .S(net299),
    .X(_04237_));
 sky130_fd_sc_hd__or2_1 _08813_ (.A(net512),
    .B(_04237_),
    .X(_01068_));
 sky130_fd_sc_hd__o22a_1 _08814_ (.A1(\tms1x00.ins_pla_ands[24][9] ),
    .A2(net299),
    .B1(_03717_),
    .B2(net364),
    .X(_01069_));
 sky130_fd_sc_hd__mux2_1 _08815_ (.A0(\tms1x00.ins_pla_ands[24][12] ),
    .A1(net963),
    .S(net299),
    .X(_04238_));
 sky130_fd_sc_hd__or2_1 _08816_ (.A(net518),
    .B(_04238_),
    .X(_01070_));
 sky130_fd_sc_hd__o22a_1 _08817_ (.A1(\tms1x00.ins_pla_ands[24][13] ),
    .A2(net299),
    .B1(_03717_),
    .B2(net363),
    .X(_01071_));
 sky130_fd_sc_hd__mux2_1 _08818_ (.A0(\tms1x00.ins_pla_ands[24][14] ),
    .A1(net951),
    .S(net299),
    .X(_04239_));
 sky130_fd_sc_hd__or2_1 _08819_ (.A(net512),
    .B(_04239_),
    .X(_01072_));
 sky130_fd_sc_hd__mux2_1 _08820_ (.A0(\tms1x00.ins_pla_ands[24][15] ),
    .A1(net944),
    .S(net299),
    .X(_04240_));
 sky130_fd_sc_hd__and2_1 _08821_ (.A(net460),
    .B(_04240_),
    .X(_01073_));
 sky130_fd_sc_hd__mux2_1 _08822_ (.A0(net1047),
    .A1(\tms1x00.ins_pla_ands[15][4] ),
    .S(net267),
    .X(_04241_));
 sky130_fd_sc_hd__or2_1 _08823_ (.A(net528),
    .B(_04241_),
    .X(_01074_));
 sky130_fd_sc_hd__or2_1 _08824_ (.A(\tms1x00.ins_pla_ands[15][5] ),
    .B(_04002_),
    .X(_04242_));
 sky130_fd_sc_hd__o211a_1 _08825_ (.A1(net1039),
    .A2(net267),
    .B1(_04242_),
    .C1(net466),
    .X(_01075_));
 sky130_fd_sc_hd__mux2_1 _08826_ (.A0(net1015),
    .A1(\tms1x00.ins_pla_ands[15][8] ),
    .S(net267),
    .X(_04243_));
 sky130_fd_sc_hd__or2_1 _08827_ (.A(net526),
    .B(_04243_),
    .X(_01076_));
 sky130_fd_sc_hd__or2_1 _08828_ (.A(\tms1x00.ins_pla_ands[15][9] ),
    .B(_04002_),
    .X(_04244_));
 sky130_fd_sc_hd__o211a_1 _08829_ (.A1(net1008),
    .A2(net267),
    .B1(_04244_),
    .C1(net463),
    .X(_01077_));
 sky130_fd_sc_hd__or2_1 _08830_ (.A(\tms1x00.ins_pla_ands[15][10] ),
    .B(_04002_),
    .X(_04245_));
 sky130_fd_sc_hd__o211a_1 _08831_ (.A1(net973),
    .A2(_04003_),
    .B1(_04245_),
    .C1(net466),
    .X(_01078_));
 sky130_fd_sc_hd__mux2_1 _08832_ (.A0(net969),
    .A1(\tms1x00.ins_pla_ands[15][11] ),
    .S(_04003_),
    .X(_04246_));
 sky130_fd_sc_hd__or2_1 _08833_ (.A(net528),
    .B(_04246_),
    .X(_01079_));
 sky130_fd_sc_hd__mux2_1 _08834_ (.A0(net964),
    .A1(\tms1x00.ins_pla_ands[15][12] ),
    .S(net267),
    .X(_04247_));
 sky130_fd_sc_hd__or2_1 _08835_ (.A(net527),
    .B(_04247_),
    .X(_01080_));
 sky130_fd_sc_hd__or2_1 _08836_ (.A(\tms1x00.ins_pla_ands[15][13] ),
    .B(_04002_),
    .X(_04248_));
 sky130_fd_sc_hd__o211a_1 _08837_ (.A1(net959),
    .A2(net267),
    .B1(_04248_),
    .C1(net463),
    .X(_01081_));
 sky130_fd_sc_hd__mux2_1 _08838_ (.A0(net952),
    .A1(\tms1x00.ins_pla_ands[15][14] ),
    .S(net267),
    .X(_04249_));
 sky130_fd_sc_hd__or2_1 _08839_ (.A(net526),
    .B(_04249_),
    .X(_01082_));
 sky130_fd_sc_hd__or2_1 _08840_ (.A(\tms1x00.ins_pla_ands[15][15] ),
    .B(_04002_),
    .X(_04250_));
 sky130_fd_sc_hd__o211a_1 _08841_ (.A1(net946),
    .A2(net267),
    .B1(_04250_),
    .C1(net463),
    .X(_01083_));
 sky130_fd_sc_hd__or2_1 _08842_ (.A(\tms1x00.ins_pla_ands[5][4] ),
    .B(_03702_),
    .X(_04251_));
 sky130_fd_sc_hd__o211a_1 _08843_ (.A1(net1050),
    .A2(_03703_),
    .B1(_04251_),
    .C1(net493),
    .X(_01084_));
 sky130_fd_sc_hd__mux2_1 _08844_ (.A0(net1043),
    .A1(\tms1x00.ins_pla_ands[5][5] ),
    .S(_03703_),
    .X(_04252_));
 sky130_fd_sc_hd__or2_1 _08845_ (.A(net557),
    .B(_04252_),
    .X(_01085_));
 sky130_fd_sc_hd__mux2_1 _08846_ (.A0(net966),
    .A1(\tms1x00.ins_pla_ands[5][12] ),
    .S(_03703_),
    .X(_04253_));
 sky130_fd_sc_hd__or2_1 _08847_ (.A(net557),
    .B(_04253_),
    .X(_01086_));
 sky130_fd_sc_hd__or2_1 _08848_ (.A(\tms1x00.ins_pla_ands[5][13] ),
    .B(_03702_),
    .X(_04254_));
 sky130_fd_sc_hd__o211a_1 _08849_ (.A1(net962),
    .A2(_03703_),
    .B1(_04254_),
    .C1(net490),
    .X(_01087_));
 sky130_fd_sc_hd__mux2_1 _08850_ (.A0(net957),
    .A1(\tms1x00.ins_pla_ands[5][14] ),
    .S(_03703_),
    .X(_04255_));
 sky130_fd_sc_hd__or2_1 _08851_ (.A(net558),
    .B(_04255_),
    .X(_01088_));
 sky130_fd_sc_hd__or2_1 _08852_ (.A(\tms1x00.ins_pla_ands[5][15] ),
    .B(_03702_),
    .X(_04256_));
 sky130_fd_sc_hd__o211a_1 _08853_ (.A1(net949),
    .A2(_03703_),
    .B1(_04256_),
    .C1(net490),
    .X(_01089_));
 sky130_fd_sc_hd__nor2_4 _08854_ (.A(net762),
    .B(net341),
    .Y(_04257_));
 sky130_fd_sc_hd__or2_1 _08855_ (.A(net762),
    .B(net341),
    .X(_04258_));
 sky130_fd_sc_hd__mux2_1 _08856_ (.A0(net980),
    .A1(\tms1x00.O_pla_ors[1][0] ),
    .S(net250),
    .X(_04259_));
 sky130_fd_sc_hd__or2_1 _08857_ (.A(net576),
    .B(_04259_),
    .X(_01090_));
 sky130_fd_sc_hd__or2_1 _08858_ (.A(\tms1x00.O_pla_ors[1][1] ),
    .B(_04257_),
    .X(_04260_));
 sky130_fd_sc_hd__o211a_1 _08859_ (.A1(net931),
    .A2(net249),
    .B1(_04260_),
    .C1(net506),
    .X(_01091_));
 sky130_fd_sc_hd__mux2_1 _08860_ (.A0(net1068),
    .A1(\tms1x00.O_pla_ors[1][2] ),
    .S(net248),
    .X(_04261_));
 sky130_fd_sc_hd__or2_1 _08861_ (.A(net574),
    .B(_04261_),
    .X(_01092_));
 sky130_fd_sc_hd__mux2_1 _08862_ (.A0(net1060),
    .A1(\tms1x00.O_pla_ors[1][3] ),
    .S(net248),
    .X(_04262_));
 sky130_fd_sc_hd__or2_1 _08863_ (.A(net574),
    .B(_04262_),
    .X(_01093_));
 sky130_fd_sc_hd__or2_1 _08864_ (.A(\tms1x00.O_pla_ors[1][4] ),
    .B(_04257_),
    .X(_04263_));
 sky130_fd_sc_hd__o211a_1 _08865_ (.A1(net1052),
    .A2(net248),
    .B1(_04263_),
    .C1(net505),
    .X(_01094_));
 sky130_fd_sc_hd__mux2_1 _08866_ (.A0(net1045),
    .A1(\tms1x00.O_pla_ors[1][5] ),
    .S(net250),
    .X(_04264_));
 sky130_fd_sc_hd__or2_1 _08867_ (.A(net576),
    .B(_04264_),
    .X(_01095_));
 sky130_fd_sc_hd__mux2_1 _08868_ (.A0(net1034),
    .A1(\tms1x00.O_pla_ors[1][6] ),
    .S(net250),
    .X(_04265_));
 sky130_fd_sc_hd__or2_1 _08869_ (.A(net576),
    .B(_04265_),
    .X(_01096_));
 sky130_fd_sc_hd__mux2_1 _08870_ (.A0(net1027),
    .A1(\tms1x00.O_pla_ors[1][7] ),
    .S(net249),
    .X(_04266_));
 sky130_fd_sc_hd__or2_1 _08871_ (.A(net569),
    .B(_04266_),
    .X(_01097_));
 sky130_fd_sc_hd__mux2_1 _08872_ (.A0(net1020),
    .A1(\tms1x00.O_pla_ors[1][8] ),
    .S(net248),
    .X(_04267_));
 sky130_fd_sc_hd__or2_1 _08873_ (.A(net574),
    .B(_04267_),
    .X(_01098_));
 sky130_fd_sc_hd__mux2_1 _08874_ (.A0(net1011),
    .A1(\tms1x00.O_pla_ors[1][9] ),
    .S(net250),
    .X(_04268_));
 sky130_fd_sc_hd__or2_1 _08875_ (.A(net570),
    .B(_04268_),
    .X(_01099_));
 sky130_fd_sc_hd__mux2_1 _08876_ (.A0(net974),
    .A1(\tms1x00.O_pla_ors[1][10] ),
    .S(net248),
    .X(_04269_));
 sky130_fd_sc_hd__or2_1 _08877_ (.A(net569),
    .B(_04269_),
    .X(_01100_));
 sky130_fd_sc_hd__or2_1 _08878_ (.A(\tms1x00.O_pla_ors[1][11] ),
    .B(_04257_),
    .X(_04270_));
 sky130_fd_sc_hd__o211a_1 _08879_ (.A1(net971),
    .A2(net248),
    .B1(_04270_),
    .C1(net503),
    .X(_01101_));
 sky130_fd_sc_hd__mux2_1 _08880_ (.A0(net967),
    .A1(\tms1x00.O_pla_ors[1][12] ),
    .S(net248),
    .X(_04271_));
 sky130_fd_sc_hd__or2_1 _08881_ (.A(net569),
    .B(_04271_),
    .X(_01102_));
 sky130_fd_sc_hd__or2_1 _08882_ (.A(\tms1x00.O_pla_ors[1][13] ),
    .B(_04257_),
    .X(_04272_));
 sky130_fd_sc_hd__o211a_1 _08883_ (.A1(net961),
    .A2(net248),
    .B1(_04272_),
    .C1(net500),
    .X(_01103_));
 sky130_fd_sc_hd__mux2_1 _08884_ (.A0(net956),
    .A1(\tms1x00.O_pla_ors[1][14] ),
    .S(net249),
    .X(_04273_));
 sky130_fd_sc_hd__or2_1 _08885_ (.A(net569),
    .B(_04273_),
    .X(_01104_));
 sky130_fd_sc_hd__mux2_1 _08886_ (.A0(net950),
    .A1(\tms1x00.O_pla_ors[1][15] ),
    .S(net248),
    .X(_04274_));
 sky130_fd_sc_hd__or2_1 _08887_ (.A(net569),
    .B(_04274_),
    .X(_01105_));
 sky130_fd_sc_hd__or2_1 _08888_ (.A(\tms1x00.O_pla_ors[1][16] ),
    .B(_04257_),
    .X(_04275_));
 sky130_fd_sc_hd__o211a_1 _08889_ (.A1(net943),
    .A2(net249),
    .B1(_04275_),
    .C1(net500),
    .X(_01106_));
 sky130_fd_sc_hd__mux2_1 _08890_ (.A0(net941),
    .A1(\tms1x00.O_pla_ors[1][17] ),
    .S(net248),
    .X(_04276_));
 sky130_fd_sc_hd__or2_1 _08891_ (.A(net569),
    .B(_04276_),
    .X(_01107_));
 sky130_fd_sc_hd__or2_1 _08892_ (.A(\tms1x00.O_pla_ors[1][18] ),
    .B(_04257_),
    .X(_04277_));
 sky130_fd_sc_hd__o211a_1 _08893_ (.A1(net939),
    .A2(net249),
    .B1(_04277_),
    .C1(net506),
    .X(_01108_));
 sky130_fd_sc_hd__or2_1 _08894_ (.A(\tms1x00.O_pla_ors[1][19] ),
    .B(_04257_),
    .X(_04278_));
 sky130_fd_sc_hd__o211a_1 _08895_ (.A1(net936),
    .A2(net250),
    .B1(_04278_),
    .C1(net501),
    .X(_01109_));
 sky130_fd_sc_hd__mux2_1 _08896_ (.A0(\tms1x00.ins_pla_ands[17][2] ),
    .A1(_03429_),
    .S(_04116_),
    .X(_01110_));
 sky130_fd_sc_hd__mux2_1 _08897_ (.A0(\tms1x00.ins_pla_ands[17][3] ),
    .A1(_03433_),
    .S(_04116_),
    .X(_01111_));
 sky130_fd_sc_hd__mux2_1 _08898_ (.A0(\tms1x00.ins_pla_ands[17][4] ),
    .A1(_03535_),
    .S(_04116_),
    .X(_01112_));
 sky130_fd_sc_hd__mux2_1 _08899_ (.A0(\tms1x00.ins_pla_ands[17][5] ),
    .A1(_03577_),
    .S(_04116_),
    .X(_01113_));
 sky130_fd_sc_hd__mux2_1 _08900_ (.A0(\tms1x00.ins_pla_ands[17][10] ),
    .A1(_03482_),
    .S(_04116_),
    .X(_01114_));
 sky130_fd_sc_hd__mux2_1 _08901_ (.A0(\tms1x00.ins_pla_ands[17][11] ),
    .A1(net347),
    .S(_04116_),
    .X(_01115_));
 sky130_fd_sc_hd__or3_1 _08902_ (.A(\tms1x00.ins_pla_ands[11][6] ),
    .B(net377),
    .C(_03952_),
    .X(_04279_));
 sky130_fd_sc_hd__o211a_1 _08903_ (.A1(_03909_),
    .A2(net271),
    .B1(_04279_),
    .C1(net383),
    .X(_01116_));
 sky130_fd_sc_hd__a31o_1 _08904_ (.A1(\tms1x00.ins_pla_ands[11][7] ),
    .A2(net370),
    .A3(net271),
    .B1(net391),
    .X(_04280_));
 sky130_fd_sc_hd__a21o_1 _08905_ (.A1(net368),
    .A2(_03952_),
    .B1(_04280_),
    .X(_01117_));
 sky130_fd_sc_hd__nor2_1 _08906_ (.A(net842),
    .B(net341),
    .Y(_04281_));
 sky130_fd_sc_hd__or2_2 _08907_ (.A(net842),
    .B(net342),
    .X(_04282_));
 sky130_fd_sc_hd__or2_1 _08908_ (.A(\tms1x00.O_pla_ors[0][0] ),
    .B(net247),
    .X(_04283_));
 sky130_fd_sc_hd__o211a_1 _08909_ (.A1(net980),
    .A2(net245),
    .B1(_04283_),
    .C1(net507),
    .X(_01118_));
 sky130_fd_sc_hd__or2_1 _08910_ (.A(\tms1x00.O_pla_ors[0][1] ),
    .B(net247),
    .X(_04284_));
 sky130_fd_sc_hd__o211a_1 _08911_ (.A1(net931),
    .A2(net245),
    .B1(_04284_),
    .C1(net506),
    .X(_01119_));
 sky130_fd_sc_hd__or2_1 _08912_ (.A(\tms1x00.O_pla_ors[0][2] ),
    .B(net246),
    .X(_04285_));
 sky130_fd_sc_hd__o211a_1 _08913_ (.A1(net1068),
    .A2(net245),
    .B1(_04285_),
    .C1(net503),
    .X(_01120_));
 sky130_fd_sc_hd__or2_1 _08914_ (.A(\tms1x00.O_pla_ors[0][3] ),
    .B(net247),
    .X(_04286_));
 sky130_fd_sc_hd__o211a_1 _08915_ (.A1(net1060),
    .A2(net245),
    .B1(_04286_),
    .C1(net503),
    .X(_01121_));
 sky130_fd_sc_hd__or2_1 _08916_ (.A(\tms1x00.O_pla_ors[0][4] ),
    .B(net246),
    .X(_04287_));
 sky130_fd_sc_hd__o211a_1 _08917_ (.A1(net1052),
    .A2(net244),
    .B1(_04287_),
    .C1(net500),
    .X(_01122_));
 sky130_fd_sc_hd__or2_1 _08918_ (.A(\tms1x00.O_pla_ors[0][5] ),
    .B(net247),
    .X(_04288_));
 sky130_fd_sc_hd__o211a_1 _08919_ (.A1(net1045),
    .A2(net245),
    .B1(_04288_),
    .C1(net507),
    .X(_01123_));
 sky130_fd_sc_hd__or2_1 _08920_ (.A(\tms1x00.O_pla_ors[0][6] ),
    .B(net247),
    .X(_04289_));
 sky130_fd_sc_hd__o211a_1 _08921_ (.A1(net1034),
    .A2(net245),
    .B1(_04289_),
    .C1(net502),
    .X(_01124_));
 sky130_fd_sc_hd__or2_1 _08922_ (.A(\tms1x00.O_pla_ors[0][7] ),
    .B(net246),
    .X(_04290_));
 sky130_fd_sc_hd__o211a_1 _08923_ (.A1(net1027),
    .A2(net244),
    .B1(_04290_),
    .C1(net500),
    .X(_01125_));
 sky130_fd_sc_hd__or2_1 _08924_ (.A(\tms1x00.O_pla_ors[0][8] ),
    .B(net246),
    .X(_04291_));
 sky130_fd_sc_hd__o211a_1 _08925_ (.A1(net1020),
    .A2(net244),
    .B1(_04291_),
    .C1(net505),
    .X(_01126_));
 sky130_fd_sc_hd__or2_1 _08926_ (.A(\tms1x00.O_pla_ors[0][9] ),
    .B(net247),
    .X(_04292_));
 sky130_fd_sc_hd__o211a_1 _08927_ (.A1(net1011),
    .A2(net245),
    .B1(_04292_),
    .C1(net501),
    .X(_01127_));
 sky130_fd_sc_hd__or2_1 _08928_ (.A(\tms1x00.O_pla_ors[0][10] ),
    .B(net247),
    .X(_04293_));
 sky130_fd_sc_hd__o211a_1 _08929_ (.A1(net975),
    .A2(net245),
    .B1(_04293_),
    .C1(net501),
    .X(_01128_));
 sky130_fd_sc_hd__or2_1 _08930_ (.A(\tms1x00.O_pla_ors[0][11] ),
    .B(net246),
    .X(_04294_));
 sky130_fd_sc_hd__o211a_1 _08931_ (.A1(net971),
    .A2(net244),
    .B1(_04294_),
    .C1(net503),
    .X(_01129_));
 sky130_fd_sc_hd__or2_1 _08932_ (.A(\tms1x00.O_pla_ors[0][12] ),
    .B(net246),
    .X(_04295_));
 sky130_fd_sc_hd__o211a_1 _08933_ (.A1(net967),
    .A2(net244),
    .B1(_04295_),
    .C1(net500),
    .X(_01130_));
 sky130_fd_sc_hd__or2_1 _08934_ (.A(\tms1x00.O_pla_ors[0][13] ),
    .B(net246),
    .X(_04296_));
 sky130_fd_sc_hd__o211a_1 _08935_ (.A1(net962),
    .A2(net244),
    .B1(_04296_),
    .C1(net500),
    .X(_01131_));
 sky130_fd_sc_hd__or2_1 _08936_ (.A(\tms1x00.O_pla_ors[0][14] ),
    .B(net246),
    .X(_04297_));
 sky130_fd_sc_hd__o211a_1 _08937_ (.A1(net956),
    .A2(net244),
    .B1(_04297_),
    .C1(net499),
    .X(_01132_));
 sky130_fd_sc_hd__or2_1 _08938_ (.A(\tms1x00.O_pla_ors[0][15] ),
    .B(net246),
    .X(_04298_));
 sky130_fd_sc_hd__o211a_1 _08939_ (.A1(net950),
    .A2(net244),
    .B1(_04298_),
    .C1(net500),
    .X(_01133_));
 sky130_fd_sc_hd__mux2_1 _08940_ (.A0(net95),
    .A1(\tms1x00.O_pla_ors[0][16] ),
    .S(net244),
    .X(_04299_));
 sky130_fd_sc_hd__or2_1 _08941_ (.A(net569),
    .B(_04299_),
    .X(_01134_));
 sky130_fd_sc_hd__or2_1 _08942_ (.A(\tms1x00.O_pla_ors[0][17] ),
    .B(net246),
    .X(_04300_));
 sky130_fd_sc_hd__o211a_1 _08943_ (.A1(net941),
    .A2(net244),
    .B1(_04300_),
    .C1(net500),
    .X(_01135_));
 sky130_fd_sc_hd__or2_1 _08944_ (.A(\tms1x00.O_pla_ors[0][18] ),
    .B(net247),
    .X(_04301_));
 sky130_fd_sc_hd__o211a_1 _08945_ (.A1(net97),
    .A2(net245),
    .B1(_04301_),
    .C1(net505),
    .X(_01136_));
 sky130_fd_sc_hd__or2_1 _08946_ (.A(\tms1x00.O_pla_ors[0][19] ),
    .B(net247),
    .X(_04302_));
 sky130_fd_sc_hd__o211a_1 _08947_ (.A1(net936),
    .A2(_04282_),
    .B1(_04302_),
    .C1(net501),
    .X(_01137_));
 sky130_fd_sc_hd__nand2_2 _08948_ (.A(net688),
    .B(_01628_),
    .Y(_04303_));
 sky130_fd_sc_hd__nor3_2 _08949_ (.A(_03378_),
    .B(_03394_),
    .C(_04303_),
    .Y(_04304_));
 sky130_fd_sc_hd__nand2_4 _08950_ (.A(\tms1x00.cycle[0] ),
    .B(_03373_),
    .Y(_04305_));
 sky130_fd_sc_hd__or3b_4 _08951_ (.A(_04305_),
    .B(\tms1x00.cycle[2] ),
    .C_N(\tms1x00.cycle[1] ),
    .X(_04306_));
 sky130_fd_sc_hd__nand2_1 _08952_ (.A(net705),
    .B(_04304_),
    .Y(_04307_));
 sky130_fd_sc_hd__a21oi_1 _08953_ (.A1(net685),
    .A2(net693),
    .B1(net705),
    .Y(_04308_));
 sky130_fd_sc_hd__a2111o_4 _08954_ (.A1(net684),
    .A2(net705),
    .B1(_02010_),
    .C1(_04308_),
    .D1(_01627_),
    .X(_04309_));
 sky130_fd_sc_hd__or2_1 _08955_ (.A(_03375_),
    .B(_03378_),
    .X(_04310_));
 sky130_fd_sc_hd__or4_1 _08956_ (.A(net688),
    .B(net693),
    .C(net144),
    .D(_04310_),
    .X(_04311_));
 sky130_fd_sc_hd__a31o_1 _08957_ (.A1(_04307_),
    .A2(_04309_),
    .A3(_04311_),
    .B1(net340),
    .X(_04312_));
 sky130_fd_sc_hd__nor2_2 _08958_ (.A(_04304_),
    .B(_04312_),
    .Y(_04313_));
 sky130_fd_sc_hd__mux2_1 _08959_ (.A0(_01628_),
    .A1(_01629_),
    .S(_01638_),
    .X(_04314_));
 sky130_fd_sc_hd__mux2_1 _08960_ (.A0(_04314_),
    .A1(\tms1x00.X[0] ),
    .S(_04309_),
    .X(_04315_));
 sky130_fd_sc_hd__nand2_1 _08961_ (.A(_04313_),
    .B(_04315_),
    .Y(_04316_));
 sky130_fd_sc_hd__o211a_1 _08962_ (.A1(\tms1x00.X[0] ),
    .A2(_04313_),
    .B1(_04316_),
    .C1(net636),
    .X(_01138_));
 sky130_fd_sc_hd__mux2_1 _08963_ (.A0(_01629_),
    .A1(_01630_),
    .S(_01638_),
    .X(_04317_));
 sky130_fd_sc_hd__mux2_1 _08964_ (.A0(_04317_),
    .A1(\tms1x00.X[1] ),
    .S(_04309_),
    .X(_04318_));
 sky130_fd_sc_hd__nand2_1 _08965_ (.A(_04313_),
    .B(_04318_),
    .Y(_04319_));
 sky130_fd_sc_hd__o211a_1 _08966_ (.A1(\tms1x00.X[1] ),
    .A2(_04313_),
    .B1(_04319_),
    .C1(net636),
    .X(_01139_));
 sky130_fd_sc_hd__mux2_1 _08967_ (.A0(\K_override[0] ),
    .A1(net1015),
    .S(net582),
    .X(_01140_));
 sky130_fd_sc_hd__mux2_1 _08968_ (.A0(\K_override[1] ),
    .A1(net1007),
    .S(net582),
    .X(_01141_));
 sky130_fd_sc_hd__mux2_1 _08969_ (.A0(\K_override[2] ),
    .A1(net973),
    .S(net582),
    .X(_01142_));
 sky130_fd_sc_hd__mux2_1 _08970_ (.A0(\K_override[3] ),
    .A1(net969),
    .S(net582),
    .X(_01143_));
 sky130_fd_sc_hd__and3_4 _08971_ (.A(net794),
    .B(net360),
    .C(net596),
    .X(_04320_));
 sky130_fd_sc_hd__or3_4 _08972_ (.A(net790),
    .B(net358),
    .C(net594),
    .X(_04321_));
 sky130_fd_sc_hd__or2_1 _08973_ (.A(\tms1x00.O_pla_ands[15][0] ),
    .B(_04320_),
    .X(_04322_));
 sky130_fd_sc_hd__o211a_1 _08974_ (.A1(net980),
    .A2(_04321_),
    .B1(_04322_),
    .C1(net508),
    .X(_01144_));
 sky130_fd_sc_hd__a21o_1 _08975_ (.A1(net931),
    .A2(_04320_),
    .B1(net575),
    .X(_04323_));
 sky130_fd_sc_hd__a21o_1 _08976_ (.A1(\tms1x00.O_pla_ands[15][1] ),
    .A2(_04321_),
    .B1(_04323_),
    .X(_01145_));
 sky130_fd_sc_hd__or2_1 _08977_ (.A(\tms1x00.O_pla_ands[15][2] ),
    .B(_04320_),
    .X(_04324_));
 sky130_fd_sc_hd__o211a_1 _08978_ (.A1(net1068),
    .A2(_04321_),
    .B1(_04324_),
    .C1(net505),
    .X(_01146_));
 sky130_fd_sc_hd__a21o_1 _08979_ (.A1(net1060),
    .A2(_04320_),
    .B1(net577),
    .X(_04325_));
 sky130_fd_sc_hd__a21o_1 _08980_ (.A1(\tms1x00.O_pla_ands[15][3] ),
    .A2(_04321_),
    .B1(_04325_),
    .X(_01147_));
 sky130_fd_sc_hd__or2_1 _08981_ (.A(\tms1x00.O_pla_ands[15][4] ),
    .B(_04320_),
    .X(_04326_));
 sky130_fd_sc_hd__o211a_1 _08982_ (.A1(net1052),
    .A2(_04321_),
    .B1(_04326_),
    .C1(net508),
    .X(_01148_));
 sky130_fd_sc_hd__a21o_1 _08983_ (.A1(net1042),
    .A2(_04320_),
    .B1(net575),
    .X(_04327_));
 sky130_fd_sc_hd__a21o_1 _08984_ (.A1(\tms1x00.O_pla_ands[15][5] ),
    .A2(_04321_),
    .B1(_04327_),
    .X(_01149_));
 sky130_fd_sc_hd__or2_1 _08985_ (.A(\tms1x00.O_pla_ands[15][6] ),
    .B(_04320_),
    .X(_04328_));
 sky130_fd_sc_hd__o211a_1 _08986_ (.A1(net1034),
    .A2(_04321_),
    .B1(_04328_),
    .C1(net508),
    .X(_01150_));
 sky130_fd_sc_hd__a21o_1 _08987_ (.A1(net1027),
    .A2(_04320_),
    .B1(net577),
    .X(_04329_));
 sky130_fd_sc_hd__a21o_1 _08988_ (.A1(\tms1x00.O_pla_ands[15][7] ),
    .A2(_04321_),
    .B1(_04329_),
    .X(_01151_));
 sky130_fd_sc_hd__or2_1 _08989_ (.A(\tms1x00.O_pla_ands[15][8] ),
    .B(_04320_),
    .X(_04330_));
 sky130_fd_sc_hd__o211a_1 _08990_ (.A1(net1020),
    .A2(_04321_),
    .B1(_04330_),
    .C1(net505),
    .X(_01152_));
 sky130_fd_sc_hd__a21o_1 _08991_ (.A1(net1011),
    .A2(_04320_),
    .B1(net575),
    .X(_04331_));
 sky130_fd_sc_hd__a21o_1 _08992_ (.A1(\tms1x00.O_pla_ands[15][9] ),
    .A2(_04321_),
    .B1(_04331_),
    .X(_01153_));
 sky130_fd_sc_hd__and3_4 _08993_ (.A(net768),
    .B(_03352_),
    .C(net359),
    .X(_04332_));
 sky130_fd_sc_hd__or3_4 _08994_ (.A(net753),
    .B(_03353_),
    .C(net357),
    .X(_04333_));
 sky130_fd_sc_hd__or2_1 _08995_ (.A(\tms1x00.O_pla_ands[17][0] ),
    .B(_04332_),
    .X(_04334_));
 sky130_fd_sc_hd__o211a_1 _08996_ (.A1(net977),
    .A2(_04333_),
    .B1(_04334_),
    .C1(net475),
    .X(_01154_));
 sky130_fd_sc_hd__or2_1 _08997_ (.A(\tms1x00.O_pla_ands[17][1] ),
    .B(_04332_),
    .X(_04335_));
 sky130_fd_sc_hd__o211a_1 _08998_ (.A1(net929),
    .A2(_04333_),
    .B1(_04335_),
    .C1(net472),
    .X(_01155_));
 sky130_fd_sc_hd__or2_1 _08999_ (.A(\tms1x00.O_pla_ands[17][2] ),
    .B(_04332_),
    .X(_04336_));
 sky130_fd_sc_hd__o211a_1 _09000_ (.A1(net1064),
    .A2(_04333_),
    .B1(_04336_),
    .C1(net471),
    .X(_01156_));
 sky130_fd_sc_hd__a21o_1 _09001_ (.A1(net1056),
    .A2(_04332_),
    .B1(net531),
    .X(_04337_));
 sky130_fd_sc_hd__a21o_1 _09002_ (.A1(\tms1x00.O_pla_ands[17][3] ),
    .A2(_04333_),
    .B1(_04337_),
    .X(_01157_));
 sky130_fd_sc_hd__or2_1 _09003_ (.A(\tms1x00.O_pla_ands[17][4] ),
    .B(_04332_),
    .X(_04338_));
 sky130_fd_sc_hd__o211a_1 _09004_ (.A1(net1048),
    .A2(_04333_),
    .B1(_04338_),
    .C1(net471),
    .X(_01158_));
 sky130_fd_sc_hd__or2_1 _09005_ (.A(\tms1x00.O_pla_ands[17][5] ),
    .B(_04332_),
    .X(_04339_));
 sky130_fd_sc_hd__o211a_1 _09006_ (.A1(net1040),
    .A2(_04333_),
    .B1(_04339_),
    .C1(net471),
    .X(_01159_));
 sky130_fd_sc_hd__or2_1 _09007_ (.A(\tms1x00.O_pla_ands[17][6] ),
    .B(_04332_),
    .X(_04340_));
 sky130_fd_sc_hd__o211a_1 _09008_ (.A1(net1031),
    .A2(_04333_),
    .B1(_04340_),
    .C1(net472),
    .X(_01160_));
 sky130_fd_sc_hd__or2_1 _09009_ (.A(\tms1x00.O_pla_ands[17][7] ),
    .B(_04332_),
    .X(_04341_));
 sky130_fd_sc_hd__o211a_1 _09010_ (.A1(net1025),
    .A2(_04333_),
    .B1(_04341_),
    .C1(net472),
    .X(_01161_));
 sky130_fd_sc_hd__a21o_1 _09011_ (.A1(net1017),
    .A2(_04332_),
    .B1(net534),
    .X(_04342_));
 sky130_fd_sc_hd__a21o_1 _09012_ (.A1(\tms1x00.O_pla_ands[17][8] ),
    .A2(_04333_),
    .B1(_04342_),
    .X(_01162_));
 sky130_fd_sc_hd__or2_1 _09013_ (.A(\tms1x00.O_pla_ands[17][9] ),
    .B(_04332_),
    .X(_04343_));
 sky130_fd_sc_hd__o211a_1 _09014_ (.A1(net1009),
    .A2(_04333_),
    .B1(_04343_),
    .C1(net471),
    .X(_01163_));
 sky130_fd_sc_hd__and3_4 _09015_ (.A(net849),
    .B(_03352_),
    .C(net359),
    .X(_04344_));
 sky130_fd_sc_hd__or3_4 _09016_ (.A(net835),
    .B(_03353_),
    .C(net357),
    .X(_04345_));
 sky130_fd_sc_hd__or2_1 _09017_ (.A(\tms1x00.O_pla_ands[16][0] ),
    .B(_04344_),
    .X(_04346_));
 sky130_fd_sc_hd__o211a_1 _09018_ (.A1(net977),
    .A2(_04345_),
    .B1(_04346_),
    .C1(net475),
    .X(_01164_));
 sky130_fd_sc_hd__a21o_1 _09019_ (.A1(net929),
    .A2(_04344_),
    .B1(net534),
    .X(_04347_));
 sky130_fd_sc_hd__a21o_1 _09020_ (.A1(\tms1x00.O_pla_ands[16][1] ),
    .A2(_04345_),
    .B1(_04347_),
    .X(_01165_));
 sky130_fd_sc_hd__or2_1 _09021_ (.A(\tms1x00.O_pla_ands[16][2] ),
    .B(_04344_),
    .X(_04348_));
 sky130_fd_sc_hd__o211a_1 _09022_ (.A1(net1064),
    .A2(_04345_),
    .B1(_04348_),
    .C1(net468),
    .X(_01166_));
 sky130_fd_sc_hd__or2_1 _09023_ (.A(\tms1x00.O_pla_ands[16][3] ),
    .B(_04344_),
    .X(_04349_));
 sky130_fd_sc_hd__o211a_1 _09024_ (.A1(net1056),
    .A2(_04345_),
    .B1(_04349_),
    .C1(net475),
    .X(_01167_));
 sky130_fd_sc_hd__or2_1 _09025_ (.A(\tms1x00.O_pla_ands[16][4] ),
    .B(_04344_),
    .X(_04350_));
 sky130_fd_sc_hd__o211a_1 _09026_ (.A1(net1048),
    .A2(_04345_),
    .B1(_04350_),
    .C1(net472),
    .X(_01168_));
 sky130_fd_sc_hd__or2_1 _09027_ (.A(\tms1x00.O_pla_ands[16][5] ),
    .B(_04344_),
    .X(_04351_));
 sky130_fd_sc_hd__o211a_1 _09028_ (.A1(net1040),
    .A2(_04345_),
    .B1(_04351_),
    .C1(net471),
    .X(_01169_));
 sky130_fd_sc_hd__or2_1 _09029_ (.A(\tms1x00.O_pla_ands[16][6] ),
    .B(_04344_),
    .X(_04352_));
 sky130_fd_sc_hd__o211a_1 _09030_ (.A1(net1031),
    .A2(_04345_),
    .B1(_04352_),
    .C1(net471),
    .X(_01170_));
 sky130_fd_sc_hd__or2_1 _09031_ (.A(\tms1x00.O_pla_ands[16][7] ),
    .B(_04344_),
    .X(_04353_));
 sky130_fd_sc_hd__o211a_1 _09032_ (.A1(net1025),
    .A2(_04345_),
    .B1(_04353_),
    .C1(net472),
    .X(_01171_));
 sky130_fd_sc_hd__a21o_1 _09033_ (.A1(net1017),
    .A2(_04344_),
    .B1(net534),
    .X(_04354_));
 sky130_fd_sc_hd__a21o_1 _09034_ (.A1(\tms1x00.O_pla_ands[16][8] ),
    .A2(_04345_),
    .B1(_04354_),
    .X(_01172_));
 sky130_fd_sc_hd__or2_1 _09035_ (.A(\tms1x00.O_pla_ands[16][9] ),
    .B(_04344_),
    .X(_04355_));
 sky130_fd_sc_hd__o211a_1 _09036_ (.A1(net1009),
    .A2(_04345_),
    .B1(_04355_),
    .C1(net471),
    .X(_01173_));
 sky130_fd_sc_hd__and3_4 _09037_ (.A(net822),
    .B(net360),
    .C(net596),
    .X(_04356_));
 sky130_fd_sc_hd__or3_4 _09038_ (.A(net816),
    .B(net358),
    .C(net594),
    .X(_04357_));
 sky130_fd_sc_hd__a21o_1 _09039_ (.A1(net980),
    .A2(_04356_),
    .B1(net575),
    .X(_04358_));
 sky130_fd_sc_hd__a21o_1 _09040_ (.A1(\tms1x00.O_pla_ands[12][0] ),
    .A2(_04357_),
    .B1(_04358_),
    .X(_01174_));
 sky130_fd_sc_hd__or2_1 _09041_ (.A(\tms1x00.O_pla_ands[12][1] ),
    .B(_04356_),
    .X(_04359_));
 sky130_fd_sc_hd__o211a_1 _09042_ (.A1(net931),
    .A2(_04357_),
    .B1(_04359_),
    .C1(net504),
    .X(_01175_));
 sky130_fd_sc_hd__a21o_1 _09043_ (.A1(net1068),
    .A2(_04356_),
    .B1(net564),
    .X(_04360_));
 sky130_fd_sc_hd__a21o_1 _09044_ (.A1(\tms1x00.O_pla_ands[12][2] ),
    .A2(_04357_),
    .B1(_04360_),
    .X(_01176_));
 sky130_fd_sc_hd__or2_1 _09045_ (.A(\tms1x00.O_pla_ands[12][3] ),
    .B(_04356_),
    .X(_04361_));
 sky130_fd_sc_hd__o211a_1 _09046_ (.A1(net1060),
    .A2(_04357_),
    .B1(_04361_),
    .C1(net504),
    .X(_01177_));
 sky130_fd_sc_hd__or2_1 _09047_ (.A(\tms1x00.O_pla_ands[12][4] ),
    .B(_04356_),
    .X(_04362_));
 sky130_fd_sc_hd__o211a_1 _09048_ (.A1(net1052),
    .A2(_04357_),
    .B1(_04362_),
    .C1(net509),
    .X(_01178_));
 sky130_fd_sc_hd__a21o_1 _09049_ (.A1(net1042),
    .A2(_04356_),
    .B1(net575),
    .X(_04363_));
 sky130_fd_sc_hd__a21o_1 _09050_ (.A1(\tms1x00.O_pla_ands[12][5] ),
    .A2(_04357_),
    .B1(_04363_),
    .X(_01179_));
 sky130_fd_sc_hd__or2_1 _09051_ (.A(\tms1x00.O_pla_ands[12][6] ),
    .B(_04356_),
    .X(_04364_));
 sky130_fd_sc_hd__o211a_1 _09052_ (.A1(net1034),
    .A2(_04357_),
    .B1(_04364_),
    .C1(net504),
    .X(_01180_));
 sky130_fd_sc_hd__a21o_1 _09053_ (.A1(net1029),
    .A2(_04356_),
    .B1(net577),
    .X(_04365_));
 sky130_fd_sc_hd__a21o_1 _09054_ (.A1(\tms1x00.O_pla_ands[12][7] ),
    .A2(_04357_),
    .B1(_04365_),
    .X(_01181_));
 sky130_fd_sc_hd__or2_1 _09055_ (.A(\tms1x00.O_pla_ands[12][8] ),
    .B(_04356_),
    .X(_04366_));
 sky130_fd_sc_hd__o211a_1 _09056_ (.A1(net1020),
    .A2(_04357_),
    .B1(_04366_),
    .C1(net504),
    .X(_01182_));
 sky130_fd_sc_hd__a21o_1 _09057_ (.A1(net1012),
    .A2(_04356_),
    .B1(net564),
    .X(_04367_));
 sky130_fd_sc_hd__a21o_1 _09058_ (.A1(\tms1x00.O_pla_ands[12][9] ),
    .A2(_04357_),
    .B1(_04367_),
    .X(_01183_));
 sky130_fd_sc_hd__and3_4 _09059_ (.A(net627),
    .B(net360),
    .C(net597),
    .X(_04368_));
 sky130_fd_sc_hd__or3_4 _09060_ (.A(net624),
    .B(net358),
    .C(net595),
    .X(_04369_));
 sky130_fd_sc_hd__a21o_1 _09061_ (.A1(net981),
    .A2(_04368_),
    .B1(net561),
    .X(_04370_));
 sky130_fd_sc_hd__a21o_1 _09062_ (.A1(\tms1x00.O_pla_ands[14][0] ),
    .A2(_04369_),
    .B1(_04370_),
    .X(_01184_));
 sky130_fd_sc_hd__or2_1 _09063_ (.A(\tms1x00.O_pla_ands[14][1] ),
    .B(_04368_),
    .X(_04371_));
 sky130_fd_sc_hd__o211a_1 _09064_ (.A1(net931),
    .A2(_04369_),
    .B1(_04371_),
    .C1(net503),
    .X(_01185_));
 sky130_fd_sc_hd__or2_1 _09065_ (.A(\tms1x00.O_pla_ands[14][2] ),
    .B(_04368_),
    .X(_04372_));
 sky130_fd_sc_hd__o211a_1 _09066_ (.A1(net1068),
    .A2(_04369_),
    .B1(_04372_),
    .C1(net503),
    .X(_01186_));
 sky130_fd_sc_hd__a21o_1 _09067_ (.A1(net1060),
    .A2(_04368_),
    .B1(net562),
    .X(_04373_));
 sky130_fd_sc_hd__a21o_1 _09068_ (.A1(\tms1x00.O_pla_ands[14][3] ),
    .A2(_04369_),
    .B1(_04373_),
    .X(_01187_));
 sky130_fd_sc_hd__or2_1 _09069_ (.A(\tms1x00.O_pla_ands[14][4] ),
    .B(_04368_),
    .X(_04374_));
 sky130_fd_sc_hd__o211a_1 _09070_ (.A1(net1050),
    .A2(_04369_),
    .B1(_04374_),
    .C1(net498),
    .X(_01188_));
 sky130_fd_sc_hd__a21o_1 _09071_ (.A1(net1042),
    .A2(_04368_),
    .B1(net562),
    .X(_04375_));
 sky130_fd_sc_hd__a21o_1 _09072_ (.A1(\tms1x00.O_pla_ands[14][5] ),
    .A2(_04369_),
    .B1(_04375_),
    .X(_01189_));
 sky130_fd_sc_hd__or2_1 _09073_ (.A(\tms1x00.O_pla_ands[14][6] ),
    .B(_04368_),
    .X(_04376_));
 sky130_fd_sc_hd__o211a_1 _09074_ (.A1(net1034),
    .A2(_04369_),
    .B1(_04376_),
    .C1(net503),
    .X(_01190_));
 sky130_fd_sc_hd__a21o_1 _09075_ (.A1(net1028),
    .A2(_04368_),
    .B1(net561),
    .X(_04377_));
 sky130_fd_sc_hd__a21o_1 _09076_ (.A1(\tms1x00.O_pla_ands[14][7] ),
    .A2(_04369_),
    .B1(_04377_),
    .X(_01191_));
 sky130_fd_sc_hd__or2_1 _09077_ (.A(\tms1x00.O_pla_ands[14][8] ),
    .B(_04368_),
    .X(_04378_));
 sky130_fd_sc_hd__o211a_1 _09078_ (.A1(net1020),
    .A2(_04369_),
    .B1(_04378_),
    .C1(net503),
    .X(_01192_));
 sky130_fd_sc_hd__a21o_1 _09079_ (.A1(net1012),
    .A2(_04368_),
    .B1(net562),
    .X(_04379_));
 sky130_fd_sc_hd__a21o_1 _09080_ (.A1(\tms1x00.O_pla_ands[14][9] ),
    .A2(_04369_),
    .B1(_04379_),
    .X(_01193_));
 sky130_fd_sc_hd__and3_4 _09081_ (.A(net904),
    .B(net360),
    .C(net597),
    .X(_04380_));
 sky130_fd_sc_hd__or3_4 _09082_ (.A(net898),
    .B(net358),
    .C(net595),
    .X(_04381_));
 sky130_fd_sc_hd__or2_1 _09083_ (.A(\tms1x00.O_pla_ands[13][0] ),
    .B(_04380_),
    .X(_04382_));
 sky130_fd_sc_hd__o211a_1 _09084_ (.A1(net980),
    .A2(_04381_),
    .B1(_04382_),
    .C1(net506),
    .X(_01194_));
 sky130_fd_sc_hd__a21o_1 _09085_ (.A1(net931),
    .A2(_04380_),
    .B1(net574),
    .X(_04383_));
 sky130_fd_sc_hd__a21o_1 _09086_ (.A1(\tms1x00.O_pla_ands[13][1] ),
    .A2(_04381_),
    .B1(_04383_),
    .X(_01195_));
 sky130_fd_sc_hd__a21o_1 _09087_ (.A1(net1068),
    .A2(_04380_),
    .B1(net574),
    .X(_04384_));
 sky130_fd_sc_hd__a21o_1 _09088_ (.A1(\tms1x00.O_pla_ands[13][2] ),
    .A2(_04381_),
    .B1(_04384_),
    .X(_01196_));
 sky130_fd_sc_hd__or2_1 _09089_ (.A(\tms1x00.O_pla_ands[13][3] ),
    .B(_04380_),
    .X(_04385_));
 sky130_fd_sc_hd__o211a_1 _09090_ (.A1(net1060),
    .A2(_04381_),
    .B1(_04385_),
    .C1(net506),
    .X(_01197_));
 sky130_fd_sc_hd__or2_1 _09091_ (.A(\tms1x00.O_pla_ands[13][4] ),
    .B(_04380_),
    .X(_04386_));
 sky130_fd_sc_hd__o211a_1 _09092_ (.A1(net1052),
    .A2(_04381_),
    .B1(_04386_),
    .C1(net506),
    .X(_01198_));
 sky130_fd_sc_hd__a21o_1 _09093_ (.A1(net1042),
    .A2(_04380_),
    .B1(net574),
    .X(_04387_));
 sky130_fd_sc_hd__a21o_1 _09094_ (.A1(\tms1x00.O_pla_ands[13][5] ),
    .A2(_04381_),
    .B1(_04387_),
    .X(_01199_));
 sky130_fd_sc_hd__or2_1 _09095_ (.A(\tms1x00.O_pla_ands[13][6] ),
    .B(_04380_),
    .X(_04388_));
 sky130_fd_sc_hd__o211a_1 _09096_ (.A1(net1034),
    .A2(_04381_),
    .B1(_04388_),
    .C1(net508),
    .X(_01200_));
 sky130_fd_sc_hd__a21o_1 _09097_ (.A1(net1029),
    .A2(_04380_),
    .B1(net574),
    .X(_04389_));
 sky130_fd_sc_hd__a21o_1 _09098_ (.A1(\tms1x00.O_pla_ands[13][7] ),
    .A2(_04381_),
    .B1(_04389_),
    .X(_01201_));
 sky130_fd_sc_hd__or2_1 _09099_ (.A(\tms1x00.O_pla_ands[13][8] ),
    .B(_04380_),
    .X(_04390_));
 sky130_fd_sc_hd__o211a_1 _09100_ (.A1(net1021),
    .A2(_04381_),
    .B1(_04390_),
    .C1(net504),
    .X(_01202_));
 sky130_fd_sc_hd__a21o_1 _09101_ (.A1(net1011),
    .A2(_04380_),
    .B1(net574),
    .X(_04391_));
 sky130_fd_sc_hd__a21o_1 _09102_ (.A1(\tms1x00.O_pla_ands[13][9] ),
    .A2(_04381_),
    .B1(_04391_),
    .X(_01203_));
 sky130_fd_sc_hd__a31o_1 _09103_ (.A1(\tms1x00.ins_pla_ors[7][27] ),
    .A2(net371),
    .A3(net302),
    .B1(net394),
    .X(_04392_));
 sky130_fd_sc_hd__a21o_1 _09104_ (.A1(_03500_),
    .A2(_03673_),
    .B1(_04392_),
    .X(_01204_));
 sky130_fd_sc_hd__a31o_1 _09105_ (.A1(\tms1x00.ins_pla_ors[7][28] ),
    .A2(net371),
    .A3(net302),
    .B1(net394),
    .X(_04393_));
 sky130_fd_sc_hd__a21o_1 _09106_ (.A1(_03449_),
    .A2(_03673_),
    .B1(_04393_),
    .X(_01205_));
 sky130_fd_sc_hd__a31o_1 _09107_ (.A1(\tms1x00.ins_pla_ors[7][29] ),
    .A2(net371),
    .A3(net302),
    .B1(net394),
    .X(_04394_));
 sky130_fd_sc_hd__a21o_1 _09108_ (.A1(_03451_),
    .A2(_03673_),
    .B1(_04394_),
    .X(_01206_));
 sky130_fd_sc_hd__and3_4 _09109_ (.A(net740),
    .B(net360),
    .C(net597),
    .X(_04395_));
 sky130_fd_sc_hd__or3_4 _09110_ (.A(net735),
    .B(net358),
    .C(net595),
    .X(_04396_));
 sky130_fd_sc_hd__a21o_1 _09111_ (.A1(net980),
    .A2(_04395_),
    .B1(net576),
    .X(_04397_));
 sky130_fd_sc_hd__a21o_1 _09112_ (.A1(\tms1x00.O_pla_ands[10][0] ),
    .A2(_04396_),
    .B1(_04397_),
    .X(_01207_));
 sky130_fd_sc_hd__or2_1 _09113_ (.A(\tms1x00.O_pla_ands[10][1] ),
    .B(_04395_),
    .X(_04398_));
 sky130_fd_sc_hd__o211a_1 _09114_ (.A1(net932),
    .A2(_04396_),
    .B1(_04398_),
    .C1(net508),
    .X(_01208_));
 sky130_fd_sc_hd__or2_1 _09115_ (.A(\tms1x00.O_pla_ands[10][2] ),
    .B(_04395_),
    .X(_04399_));
 sky130_fd_sc_hd__o211a_1 _09116_ (.A1(net1069),
    .A2(_04396_),
    .B1(_04399_),
    .C1(net508),
    .X(_01209_));
 sky130_fd_sc_hd__a21o_1 _09117_ (.A1(net1061),
    .A2(_04395_),
    .B1(net577),
    .X(_04400_));
 sky130_fd_sc_hd__a21o_1 _09118_ (.A1(\tms1x00.O_pla_ands[10][3] ),
    .A2(_04396_),
    .B1(_04400_),
    .X(_01210_));
 sky130_fd_sc_hd__a21o_1 _09119_ (.A1(net1052),
    .A2(_04395_),
    .B1(net577),
    .X(_04401_));
 sky130_fd_sc_hd__a21o_1 _09120_ (.A1(\tms1x00.O_pla_ands[10][4] ),
    .A2(_04396_),
    .B1(_04401_),
    .X(_01211_));
 sky130_fd_sc_hd__or2_1 _09121_ (.A(\tms1x00.O_pla_ands[10][5] ),
    .B(_04395_),
    .X(_04402_));
 sky130_fd_sc_hd__o211a_1 _09122_ (.A1(net1042),
    .A2(_04396_),
    .B1(_04402_),
    .C1(net505),
    .X(_01212_));
 sky130_fd_sc_hd__or2_1 _09123_ (.A(\tms1x00.O_pla_ands[10][6] ),
    .B(_04395_),
    .X(_04403_));
 sky130_fd_sc_hd__o211a_1 _09124_ (.A1(net1035),
    .A2(_04396_),
    .B1(_04403_),
    .C1(net508),
    .X(_01213_));
 sky130_fd_sc_hd__a21o_1 _09125_ (.A1(net1029),
    .A2(_04395_),
    .B1(net577),
    .X(_04404_));
 sky130_fd_sc_hd__a21o_1 _09126_ (.A1(\tms1x00.O_pla_ands[10][7] ),
    .A2(_04396_),
    .B1(_04404_),
    .X(_01214_));
 sky130_fd_sc_hd__or2_1 _09127_ (.A(\tms1x00.O_pla_ands[10][8] ),
    .B(_04395_),
    .X(_04405_));
 sky130_fd_sc_hd__o211a_1 _09128_ (.A1(net1021),
    .A2(_04396_),
    .B1(_04405_),
    .C1(net504),
    .X(_01215_));
 sky130_fd_sc_hd__a21o_1 _09129_ (.A1(net1013),
    .A2(_04395_),
    .B1(net577),
    .X(_04406_));
 sky130_fd_sc_hd__a21o_1 _09130_ (.A1(\tms1x00.O_pla_ands[10][9] ),
    .A2(_04396_),
    .B1(_04406_),
    .X(_01216_));
 sky130_fd_sc_hd__and3_4 _09131_ (.A(net767),
    .B(net360),
    .C(net597),
    .X(_04407_));
 sky130_fd_sc_hd__or3_4 _09132_ (.A(net765),
    .B(net358),
    .C(net595),
    .X(_04408_));
 sky130_fd_sc_hd__or2_1 _09133_ (.A(\tms1x00.O_pla_ands[9][0] ),
    .B(_04407_),
    .X(_04409_));
 sky130_fd_sc_hd__o211a_1 _09134_ (.A1(net981),
    .A2(_04408_),
    .B1(_04409_),
    .C1(net498),
    .X(_01217_));
 sky130_fd_sc_hd__a21o_1 _09135_ (.A1(net931),
    .A2(_04407_),
    .B1(net563),
    .X(_04410_));
 sky130_fd_sc_hd__a21o_1 _09136_ (.A1(\tms1x00.O_pla_ands[9][1] ),
    .A2(_04408_),
    .B1(_04410_),
    .X(_01218_));
 sky130_fd_sc_hd__a21o_1 _09137_ (.A1(net1068),
    .A2(_04407_),
    .B1(net564),
    .X(_04411_));
 sky130_fd_sc_hd__a21o_1 _09138_ (.A1(\tms1x00.O_pla_ands[9][2] ),
    .A2(_04408_),
    .B1(_04411_),
    .X(_01219_));
 sky130_fd_sc_hd__or2_1 _09139_ (.A(\tms1x00.O_pla_ands[9][3] ),
    .B(_04407_),
    .X(_04412_));
 sky130_fd_sc_hd__o211a_1 _09140_ (.A1(net1059),
    .A2(_04408_),
    .B1(_04412_),
    .C1(net497),
    .X(_01220_));
 sky130_fd_sc_hd__a21o_1 _09141_ (.A1(net1050),
    .A2(_04407_),
    .B1(net563),
    .X(_04413_));
 sky130_fd_sc_hd__a21o_1 _09142_ (.A1(\tms1x00.O_pla_ands[9][4] ),
    .A2(_04408_),
    .B1(_04413_),
    .X(_01221_));
 sky130_fd_sc_hd__or2_1 _09143_ (.A(\tms1x00.O_pla_ands[9][5] ),
    .B(_04407_),
    .X(_04414_));
 sky130_fd_sc_hd__o211a_1 _09144_ (.A1(net1043),
    .A2(_04408_),
    .B1(_04414_),
    .C1(net497),
    .X(_01222_));
 sky130_fd_sc_hd__or2_1 _09145_ (.A(\tms1x00.O_pla_ands[9][6] ),
    .B(_04407_),
    .X(_04415_));
 sky130_fd_sc_hd__o211a_1 _09146_ (.A1(net1036),
    .A2(_04408_),
    .B1(_04415_),
    .C1(net497),
    .X(_01223_));
 sky130_fd_sc_hd__a21o_1 _09147_ (.A1(net1028),
    .A2(_04407_),
    .B1(net563),
    .X(_04416_));
 sky130_fd_sc_hd__a21o_1 _09148_ (.A1(\tms1x00.O_pla_ands[9][7] ),
    .A2(_04408_),
    .B1(_04416_),
    .X(_01224_));
 sky130_fd_sc_hd__or2_1 _09149_ (.A(\tms1x00.O_pla_ands[9][8] ),
    .B(_04407_),
    .X(_04417_));
 sky130_fd_sc_hd__o211a_1 _09150_ (.A1(net1020),
    .A2(_04408_),
    .B1(_04417_),
    .C1(net497),
    .X(_01225_));
 sky130_fd_sc_hd__a21o_1 _09151_ (.A1(net1012),
    .A2(_04407_),
    .B1(net563),
    .X(_04418_));
 sky130_fd_sc_hd__a21o_1 _09152_ (.A1(\tms1x00.O_pla_ands[9][9] ),
    .A2(_04408_),
    .B1(_04418_),
    .X(_01226_));
 sky130_fd_sc_hd__and3_4 _09153_ (.A(net876),
    .B(net360),
    .C(net597),
    .X(_04419_));
 sky130_fd_sc_hd__or3_4 _09154_ (.A(net869),
    .B(net358),
    .C(net595),
    .X(_04420_));
 sky130_fd_sc_hd__or2_1 _09155_ (.A(\tms1x00.O_pla_ands[11][0] ),
    .B(_04419_),
    .X(_04421_));
 sky130_fd_sc_hd__o211a_1 _09156_ (.A1(net981),
    .A2(_04420_),
    .B1(_04421_),
    .C1(net498),
    .X(_01227_));
 sky130_fd_sc_hd__a21o_1 _09157_ (.A1(net933),
    .A2(_04419_),
    .B1(net564),
    .X(_04422_));
 sky130_fd_sc_hd__a21o_1 _09158_ (.A1(\tms1x00.O_pla_ands[11][1] ),
    .A2(_04420_),
    .B1(_04422_),
    .X(_01228_));
 sky130_fd_sc_hd__or2_1 _09159_ (.A(\tms1x00.O_pla_ands[11][2] ),
    .B(_04419_),
    .X(_04423_));
 sky130_fd_sc_hd__o211a_1 _09160_ (.A1(net1067),
    .A2(_04420_),
    .B1(_04423_),
    .C1(net497),
    .X(_01229_));
 sky130_fd_sc_hd__a21o_1 _09161_ (.A1(net1059),
    .A2(_04419_),
    .B1(net561),
    .X(_04424_));
 sky130_fd_sc_hd__a21o_1 _09162_ (.A1(\tms1x00.O_pla_ands[11][3] ),
    .A2(_04420_),
    .B1(_04424_),
    .X(_01230_));
 sky130_fd_sc_hd__a21o_1 _09163_ (.A1(net1051),
    .A2(_04419_),
    .B1(net563),
    .X(_04425_));
 sky130_fd_sc_hd__a21o_1 _09164_ (.A1(\tms1x00.O_pla_ands[11][4] ),
    .A2(_04420_),
    .B1(_04425_),
    .X(_01231_));
 sky130_fd_sc_hd__or2_1 _09165_ (.A(\tms1x00.O_pla_ands[11][5] ),
    .B(_04419_),
    .X(_04426_));
 sky130_fd_sc_hd__o211a_1 _09166_ (.A1(net1043),
    .A2(_04420_),
    .B1(_04426_),
    .C1(net497),
    .X(_01232_));
 sky130_fd_sc_hd__or2_1 _09167_ (.A(\tms1x00.O_pla_ands[11][6] ),
    .B(_04419_),
    .X(_04427_));
 sky130_fd_sc_hd__o211a_1 _09168_ (.A1(net1036),
    .A2(_04420_),
    .B1(_04427_),
    .C1(net498),
    .X(_01233_));
 sky130_fd_sc_hd__a21o_1 _09169_ (.A1(net1028),
    .A2(_04419_),
    .B1(net563),
    .X(_04428_));
 sky130_fd_sc_hd__a21o_1 _09170_ (.A1(\tms1x00.O_pla_ands[11][7] ),
    .A2(_04420_),
    .B1(_04428_),
    .X(_01234_));
 sky130_fd_sc_hd__or2_1 _09171_ (.A(\tms1x00.O_pla_ands[11][8] ),
    .B(_04419_),
    .X(_04429_));
 sky130_fd_sc_hd__o211a_1 _09172_ (.A1(net1020),
    .A2(_04420_),
    .B1(_04429_),
    .C1(net497),
    .X(_01235_));
 sky130_fd_sc_hd__a21o_1 _09173_ (.A1(net1012),
    .A2(_04419_),
    .B1(net564),
    .X(_04430_));
 sky130_fd_sc_hd__a21o_1 _09174_ (.A1(\tms1x00.O_pla_ands[11][9] ),
    .A2(_04420_),
    .B1(_04430_),
    .X(_01236_));
 sky130_fd_sc_hd__nor2_2 _09175_ (.A(net380),
    .B(_03545_),
    .Y(_04431_));
 sky130_fd_sc_hd__nand2_2 _09176_ (.A(net386),
    .B(net320),
    .Y(_04432_));
 sky130_fd_sc_hd__a22o_1 _09177_ (.A1(\tms1x00.ins_pla_ors[3][2] ),
    .A2(_04431_),
    .B1(_04432_),
    .B2(_03429_),
    .X(_01237_));
 sky130_fd_sc_hd__a22o_1 _09178_ (.A1(\tms1x00.ins_pla_ors[3][3] ),
    .A2(_04431_),
    .B1(_04432_),
    .B2(_03534_),
    .X(_01238_));
 sky130_fd_sc_hd__a21o_1 _09179_ (.A1(net388),
    .A2(net320),
    .B1(_03536_),
    .X(_04433_));
 sky130_fd_sc_hd__o31a_1 _09180_ (.A1(\tms1x00.ins_pla_ors[3][7] ),
    .A2(net382),
    .A3(_03545_),
    .B1(_04433_),
    .X(_01239_));
 sky130_fd_sc_hd__a22o_1 _09181_ (.A1(\tms1x00.ins_pla_ors[3][12] ),
    .A2(_04431_),
    .B1(_04432_),
    .B2(_03588_),
    .X(_01240_));
 sky130_fd_sc_hd__mux2_1 _09182_ (.A0(net955),
    .A1(\tms1x00.ins_pla_ors[3][14] ),
    .S(net321),
    .X(_04434_));
 sky130_fd_sc_hd__o21a_1 _09183_ (.A1(net379),
    .A2(_04434_),
    .B1(net387),
    .X(_01241_));
 sky130_fd_sc_hd__mux2_1 _09184_ (.A0(net101),
    .A1(\tms1x00.ins_pla_ors[3][21] ),
    .S(net321),
    .X(_04435_));
 sky130_fd_sc_hd__o21a_1 _09185_ (.A1(net548),
    .A2(_04435_),
    .B1(net372),
    .X(_01242_));
 sky130_fd_sc_hd__a221o_1 _09186_ (.A1(_03467_),
    .A2(_03545_),
    .B1(_04431_),
    .B2(\tms1x00.ins_pla_ors[3][24] ),
    .C1(net395),
    .X(_01243_));
 sky130_fd_sc_hd__mux2_1 _09187_ (.A0(net105),
    .A1(\tms1x00.ins_pla_ors[3][25] ),
    .S(net320),
    .X(_04436_));
 sky130_fd_sc_hd__o21a_1 _09188_ (.A1(net379),
    .A2(_04436_),
    .B1(net386),
    .X(_01244_));
 sky130_fd_sc_hd__a22o_1 _09189_ (.A1(\tms1x00.ins_pla_ors[3][29] ),
    .A2(_04431_),
    .B1(_04432_),
    .B2(_03452_),
    .X(_01245_));
 sky130_fd_sc_hd__nor2_4 _09190_ (.A(net380),
    .B(_03768_),
    .Y(_04437_));
 sky130_fd_sc_hd__nand2_1 _09191_ (.A(net372),
    .B(net293),
    .Y(_04438_));
 sky130_fd_sc_hd__nor2_1 _09192_ (.A(net394),
    .B(_03768_),
    .Y(_04439_));
 sky130_fd_sc_hd__nand2_4 _09193_ (.A(net386),
    .B(net293),
    .Y(_04440_));
 sky130_fd_sc_hd__a22o_1 _09194_ (.A1(\tms1x00.ins_pla_ors[6][7] ),
    .A2(_04437_),
    .B1(_04440_),
    .B2(_03437_),
    .X(_01246_));
 sky130_fd_sc_hd__a22o_1 _09195_ (.A1(\tms1x00.ins_pla_ors[6][8] ),
    .A2(_04437_),
    .B1(_04440_),
    .B2(_03439_),
    .X(_01247_));
 sky130_fd_sc_hd__o22a_1 _09196_ (.A1(\tms1x00.ins_pla_ors[6][12] ),
    .A2(_04438_),
    .B1(_04439_),
    .B2(_03485_),
    .X(_01248_));
 sky130_fd_sc_hd__o22a_1 _09197_ (.A1(\tms1x00.ins_pla_ors[6][16] ),
    .A2(_04438_),
    .B1(_04439_),
    .B2(_03441_),
    .X(_01249_));
 sky130_fd_sc_hd__o221a_1 _09198_ (.A1(_03444_),
    .A2(net293),
    .B1(_04438_),
    .B2(\tms1x00.ins_pla_ors[6][18] ),
    .C1(net386),
    .X(_01250_));
 sky130_fd_sc_hd__a221o_1 _09199_ (.A1(_03498_),
    .A2(_03768_),
    .B1(_04437_),
    .B2(\tms1x00.ins_pla_ors[6][25] ),
    .C1(net394),
    .X(_01251_));
 sky130_fd_sc_hd__mux2_1 _09200_ (.A0(net106),
    .A1(\tms1x00.ins_pla_ors[6][26] ),
    .S(net295),
    .X(_04441_));
 sky130_fd_sc_hd__a21o_1 _09201_ (.A1(net484),
    .A2(_04441_),
    .B1(net379),
    .X(_01252_));
 sky130_fd_sc_hd__a22o_1 _09202_ (.A1(\tms1x00.ins_pla_ors[6][27] ),
    .A2(_04437_),
    .B1(_04440_),
    .B2(_03636_),
    .X(_01253_));
 sky130_fd_sc_hd__a22o_1 _09203_ (.A1(\tms1x00.ins_pla_ors[6][28] ),
    .A2(_04437_),
    .B1(_04440_),
    .B2(_03450_),
    .X(_01254_));
 sky130_fd_sc_hd__a22o_1 _09204_ (.A1(\tms1x00.ins_pla_ors[6][29] ),
    .A2(_04437_),
    .B1(_04440_),
    .B2(_03452_),
    .X(_01255_));
 sky130_fd_sc_hd__nor2_4 _09205_ (.A(net381),
    .B(_03821_),
    .Y(_04442_));
 sky130_fd_sc_hd__nand2_2 _09206_ (.A(net373),
    .B(net282),
    .Y(_04443_));
 sky130_fd_sc_hd__o221a_1 _09207_ (.A1(_03574_),
    .A2(net280),
    .B1(_04443_),
    .B2(\tms1x00.ins_pla_ors[5][0] ),
    .C1(net385),
    .X(_01256_));
 sky130_fd_sc_hd__nor2_2 _09208_ (.A(net395),
    .B(_03821_),
    .Y(_04444_));
 sky130_fd_sc_hd__nand2_4 _09209_ (.A(net385),
    .B(net280),
    .Y(_04445_));
 sky130_fd_sc_hd__a22o_1 _09210_ (.A1(\tms1x00.ins_pla_ors[5][1] ),
    .A2(_04442_),
    .B1(_04445_),
    .B2(_03427_),
    .X(_01257_));
 sky130_fd_sc_hd__o22a_1 _09211_ (.A1(\tms1x00.ins_pla_ors[5][3] ),
    .A2(_04443_),
    .B1(_04444_),
    .B2(_03433_),
    .X(_01258_));
 sky130_fd_sc_hd__o22a_1 _09212_ (.A1(\tms1x00.ins_pla_ors[5][4] ),
    .A2(_04443_),
    .B1(_04444_),
    .B2(_03479_),
    .X(_01259_));
 sky130_fd_sc_hd__o22a_1 _09213_ (.A1(\tms1x00.ins_pla_ors[5][7] ),
    .A2(_04443_),
    .B1(_04444_),
    .B2(_03536_),
    .X(_01260_));
 sky130_fd_sc_hd__or3_1 _09214_ (.A(net1022),
    .B(net381),
    .C(net280),
    .X(_04446_));
 sky130_fd_sc_hd__o211a_1 _09215_ (.A1(\tms1x00.ins_pla_ors[5][8] ),
    .A2(_04443_),
    .B1(_04446_),
    .C1(net385),
    .X(_01261_));
 sky130_fd_sc_hd__mux2_1 _09216_ (.A0(net943),
    .A1(\tms1x00.ins_pla_ors[5][16] ),
    .S(net281),
    .X(_04447_));
 sky130_fd_sc_hd__o21a_1 _09217_ (.A1(net547),
    .A2(_04447_),
    .B1(net371),
    .X(_01262_));
 sky130_fd_sc_hd__mux2_1 _09218_ (.A0(net101),
    .A1(\tms1x00.ins_pla_ors[5][21] ),
    .S(net281),
    .X(_04448_));
 sky130_fd_sc_hd__o21a_1 _09219_ (.A1(net379),
    .A2(_04448_),
    .B1(net387),
    .X(_01263_));
 sky130_fd_sc_hd__a221o_1 _09220_ (.A1(_03467_),
    .A2(_03821_),
    .B1(_04442_),
    .B2(\tms1x00.ins_pla_ors[5][24] ),
    .C1(net394),
    .X(_01264_));
 sky130_fd_sc_hd__and3_1 _09221_ (.A(\tms1x00.ins_pla_ors[5][26] ),
    .B(net371),
    .C(net280),
    .X(_04449_));
 sky130_fd_sc_hd__a31o_1 _09222_ (.A1(net371),
    .A2(_03447_),
    .A3(_04445_),
    .B1(_04449_),
    .X(_01265_));
 sky130_fd_sc_hd__a22o_1 _09223_ (.A1(\tms1x00.ins_pla_ors[5][27] ),
    .A2(_04442_),
    .B1(_04445_),
    .B2(_03636_),
    .X(_01266_));
 sky130_fd_sc_hd__a22o_1 _09224_ (.A1(\tms1x00.ins_pla_ors[5][28] ),
    .A2(_04442_),
    .B1(_04445_),
    .B2(_03450_),
    .X(_01267_));
 sky130_fd_sc_hd__a22o_1 _09225_ (.A1(\tms1x00.ins_pla_ors[5][29] ),
    .A2(_04442_),
    .B1(_04445_),
    .B2(_03452_),
    .X(_01268_));
 sky130_fd_sc_hd__nor2_4 _09226_ (.A(net380),
    .B(_03502_),
    .Y(_04450_));
 sky130_fd_sc_hd__nand2_1 _09227_ (.A(net372),
    .B(net330),
    .Y(_04451_));
 sky130_fd_sc_hd__nor2_1 _09228_ (.A(net395),
    .B(_03502_),
    .Y(_04452_));
 sky130_fd_sc_hd__nand2_4 _09229_ (.A(net385),
    .B(net330),
    .Y(_04453_));
 sky130_fd_sc_hd__a22o_1 _09230_ (.A1(\tms1x00.ins_pla_ors[4][5] ),
    .A2(_04450_),
    .B1(_04453_),
    .B2(_03712_),
    .X(_01269_));
 sky130_fd_sc_hd__a22o_1 _09231_ (.A1(\tms1x00.ins_pla_ors[4][6] ),
    .A2(_04450_),
    .B1(_04453_),
    .B2(_03435_),
    .X(_01270_));
 sky130_fd_sc_hd__a22o_1 _09232_ (.A1(\tms1x00.ins_pla_ors[4][8] ),
    .A2(_04450_),
    .B1(_04453_),
    .B2(net353),
    .X(_01271_));
 sky130_fd_sc_hd__o22a_1 _09233_ (.A1(\tms1x00.ins_pla_ors[4][11] ),
    .A2(_04451_),
    .B1(_04452_),
    .B2(_03580_),
    .X(_01272_));
 sky130_fd_sc_hd__mux2_1 _09234_ (.A0(net957),
    .A1(\tms1x00.ins_pla_ors[4][14] ),
    .S(net330),
    .X(_04454_));
 sky130_fd_sc_hd__o21a_1 _09235_ (.A1(net538),
    .A2(_04454_),
    .B1(net371),
    .X(_01273_));
 sky130_fd_sc_hd__o22a_1 _09236_ (.A1(\tms1x00.ins_pla_ors[4][16] ),
    .A2(_04451_),
    .B1(_04452_),
    .B2(_03441_),
    .X(_01274_));
 sky130_fd_sc_hd__mux2_1 _09237_ (.A0(net941),
    .A1(\tms1x00.ins_pla_ors[4][17] ),
    .S(_03503_),
    .X(_04455_));
 sky130_fd_sc_hd__o21a_1 _09238_ (.A1(net379),
    .A2(_04455_),
    .B1(net387),
    .X(_01275_));
 sky130_fd_sc_hd__o221a_1 _09239_ (.A1(_03444_),
    .A2(net331),
    .B1(_04451_),
    .B2(\tms1x00.ins_pla_ors[4][18] ),
    .C1(net385),
    .X(_01276_));
 sky130_fd_sc_hd__mux2_1 _09240_ (.A0(net104),
    .A1(\tms1x00.ins_pla_ors[4][24] ),
    .S(_03503_),
    .X(_04456_));
 sky130_fd_sc_hd__o21a_1 _09241_ (.A1(net380),
    .A2(_04456_),
    .B1(net387),
    .X(_01277_));
 sky130_fd_sc_hd__a221o_1 _09242_ (.A1(_03498_),
    .A2(_03502_),
    .B1(_04450_),
    .B2(\tms1x00.ins_pla_ors[4][25] ),
    .C1(net394),
    .X(_01278_));
 sky130_fd_sc_hd__and3_1 _09243_ (.A(\tms1x00.ins_pla_ors[4][26] ),
    .B(net371),
    .C(net330),
    .X(_04457_));
 sky130_fd_sc_hd__a31o_1 _09244_ (.A1(net371),
    .A2(_03447_),
    .A3(_04453_),
    .B1(_04457_),
    .X(_01279_));
 sky130_fd_sc_hd__a22o_1 _09245_ (.A1(\tms1x00.ins_pla_ors[4][27] ),
    .A2(_04450_),
    .B1(_04453_),
    .B2(_03636_),
    .X(_01280_));
 sky130_fd_sc_hd__a22o_1 _09246_ (.A1(\tms1x00.ins_pla_ors[4][28] ),
    .A2(_04450_),
    .B1(_04453_),
    .B2(_03450_),
    .X(_01281_));
 sky130_fd_sc_hd__a22o_1 _09247_ (.A1(\tms1x00.ins_pla_ors[4][29] ),
    .A2(_04450_),
    .B1(_04453_),
    .B2(_03452_),
    .X(_01282_));
 sky130_fd_sc_hd__and3_4 _09248_ (.A(net795),
    .B(net359),
    .C(net709),
    .X(_04458_));
 sky130_fd_sc_hd__or3_4 _09249_ (.A(net781),
    .B(net358),
    .C(net706),
    .X(_04459_));
 sky130_fd_sc_hd__or2_1 _09250_ (.A(\tms1x00.O_pla_ands[7][0] ),
    .B(_04458_),
    .X(_04460_));
 sky130_fd_sc_hd__o211a_1 _09251_ (.A1(net977),
    .A2(_04459_),
    .B1(_04460_),
    .C1(net476),
    .X(_01283_));
 sky130_fd_sc_hd__a21o_1 _09252_ (.A1(net929),
    .A2(_04458_),
    .B1(net531),
    .X(_04461_));
 sky130_fd_sc_hd__a21o_1 _09253_ (.A1(\tms1x00.O_pla_ands[7][1] ),
    .A2(_04459_),
    .B1(_04461_),
    .X(_01284_));
 sky130_fd_sc_hd__or2_1 _09254_ (.A(\tms1x00.O_pla_ands[7][2] ),
    .B(_04458_),
    .X(_04462_));
 sky130_fd_sc_hd__o211a_1 _09255_ (.A1(net1067),
    .A2(_04459_),
    .B1(_04462_),
    .C1(net476),
    .X(_01285_));
 sky130_fd_sc_hd__a21o_1 _09256_ (.A1(net1056),
    .A2(_04458_),
    .B1(net533),
    .X(_04463_));
 sky130_fd_sc_hd__a21o_1 _09257_ (.A1(\tms1x00.O_pla_ands[7][3] ),
    .A2(_04459_),
    .B1(_04463_),
    .X(_01286_));
 sky130_fd_sc_hd__or2_1 _09258_ (.A(\tms1x00.O_pla_ands[7][4] ),
    .B(_04458_),
    .X(_04464_));
 sky130_fd_sc_hd__o211a_1 _09259_ (.A1(net1051),
    .A2(_04459_),
    .B1(_04464_),
    .C1(net475),
    .X(_01287_));
 sky130_fd_sc_hd__a21o_1 _09260_ (.A1(net1040),
    .A2(_04458_),
    .B1(net531),
    .X(_04465_));
 sky130_fd_sc_hd__a21o_1 _09261_ (.A1(\tms1x00.O_pla_ands[7][5] ),
    .A2(_04459_),
    .B1(_04465_),
    .X(_01288_));
 sky130_fd_sc_hd__a21o_1 _09262_ (.A1(net1031),
    .A2(_04458_),
    .B1(net531),
    .X(_04466_));
 sky130_fd_sc_hd__a21o_1 _09263_ (.A1(\tms1x00.O_pla_ands[7][6] ),
    .A2(_04459_),
    .B1(_04466_),
    .X(_01289_));
 sky130_fd_sc_hd__or2_1 _09264_ (.A(\tms1x00.O_pla_ands[7][7] ),
    .B(_04458_),
    .X(_04467_));
 sky130_fd_sc_hd__o211a_1 _09265_ (.A1(net1025),
    .A2(_04459_),
    .B1(_04467_),
    .C1(net475),
    .X(_01290_));
 sky130_fd_sc_hd__or2_1 _09266_ (.A(\tms1x00.O_pla_ands[7][8] ),
    .B(_04458_),
    .X(_04468_));
 sky130_fd_sc_hd__o211a_1 _09267_ (.A1(net1019),
    .A2(_04459_),
    .B1(_04468_),
    .C1(net475),
    .X(_01291_));
 sky130_fd_sc_hd__a21o_1 _09268_ (.A1(net1009),
    .A2(_04458_),
    .B1(net531),
    .X(_04469_));
 sky130_fd_sc_hd__a21o_1 _09269_ (.A1(\tms1x00.O_pla_ands[7][9] ),
    .A2(_04459_),
    .B1(_04469_),
    .X(_01292_));
 sky130_fd_sc_hd__and3_4 _09270_ (.A(net849),
    .B(_03356_),
    .C(net597),
    .X(_04470_));
 sky130_fd_sc_hd__or3_4 _09271_ (.A(net843),
    .B(net358),
    .C(net595),
    .X(_04471_));
 sky130_fd_sc_hd__a21o_1 _09272_ (.A1(net981),
    .A2(_04470_),
    .B1(net575),
    .X(_04472_));
 sky130_fd_sc_hd__a21o_1 _09273_ (.A1(\tms1x00.O_pla_ands[8][0] ),
    .A2(_04471_),
    .B1(_04472_),
    .X(_01293_));
 sky130_fd_sc_hd__or2_1 _09274_ (.A(\tms1x00.O_pla_ands[8][1] ),
    .B(_04470_),
    .X(_04473_));
 sky130_fd_sc_hd__o211a_1 _09275_ (.A1(net931),
    .A2(_04471_),
    .B1(_04473_),
    .C1(net504),
    .X(_01294_));
 sky130_fd_sc_hd__a21o_1 _09276_ (.A1(net1068),
    .A2(_04470_),
    .B1(net575),
    .X(_04474_));
 sky130_fd_sc_hd__a21o_1 _09277_ (.A1(\tms1x00.O_pla_ands[8][2] ),
    .A2(_04471_),
    .B1(_04474_),
    .X(_01295_));
 sky130_fd_sc_hd__or2_1 _09278_ (.A(\tms1x00.O_pla_ands[8][3] ),
    .B(_04470_),
    .X(_04475_));
 sky130_fd_sc_hd__o211a_1 _09279_ (.A1(net1061),
    .A2(_04471_),
    .B1(_04475_),
    .C1(net508),
    .X(_01296_));
 sky130_fd_sc_hd__a21o_1 _09280_ (.A1(net1052),
    .A2(_04470_),
    .B1(net575),
    .X(_04476_));
 sky130_fd_sc_hd__a21o_1 _09281_ (.A1(\tms1x00.O_pla_ands[8][4] ),
    .A2(_04471_),
    .B1(_04476_),
    .X(_01297_));
 sky130_fd_sc_hd__or2_1 _09282_ (.A(\tms1x00.O_pla_ands[8][5] ),
    .B(_04470_),
    .X(_04477_));
 sky130_fd_sc_hd__o211a_1 _09283_ (.A1(net1042),
    .A2(_04471_),
    .B1(_04477_),
    .C1(net504),
    .X(_01298_));
 sky130_fd_sc_hd__or2_1 _09284_ (.A(\tms1x00.O_pla_ands[8][6] ),
    .B(_04470_),
    .X(_04478_));
 sky130_fd_sc_hd__o211a_1 _09285_ (.A1(net1034),
    .A2(_04471_),
    .B1(_04478_),
    .C1(net504),
    .X(_01299_));
 sky130_fd_sc_hd__a21o_1 _09286_ (.A1(net1029),
    .A2(_04470_),
    .B1(net575),
    .X(_04479_));
 sky130_fd_sc_hd__a21o_1 _09287_ (.A1(\tms1x00.O_pla_ands[8][7] ),
    .A2(_04471_),
    .B1(_04479_),
    .X(_01300_));
 sky130_fd_sc_hd__or2_1 _09288_ (.A(\tms1x00.O_pla_ands[8][8] ),
    .B(_04470_),
    .X(_04480_));
 sky130_fd_sc_hd__o211a_1 _09289_ (.A1(net1021),
    .A2(_04471_),
    .B1(_04480_),
    .C1(net504),
    .X(_01301_));
 sky130_fd_sc_hd__a21o_1 _09290_ (.A1(net117),
    .A2(_04470_),
    .B1(net575),
    .X(_04481_));
 sky130_fd_sc_hd__a21o_1 _09291_ (.A1(\tms1x00.O_pla_ands[8][9] ),
    .A2(_04471_),
    .B1(_04481_),
    .X(_01302_));
 sky130_fd_sc_hd__and3_4 _09292_ (.A(net741),
    .B(net359),
    .C(net709),
    .X(_04482_));
 sky130_fd_sc_hd__or3_4 _09293_ (.A(net733),
    .B(net357),
    .C(net706),
    .X(_04483_));
 sky130_fd_sc_hd__a21o_1 _09294_ (.A1(net981),
    .A2(_04482_),
    .B1(net563),
    .X(_04484_));
 sky130_fd_sc_hd__a21o_1 _09295_ (.A1(\tms1x00.O_pla_ands[2][0] ),
    .A2(_04483_),
    .B1(_04484_),
    .X(_01303_));
 sky130_fd_sc_hd__or2_1 _09296_ (.A(\tms1x00.O_pla_ands[2][1] ),
    .B(_04482_),
    .X(_04485_));
 sky130_fd_sc_hd__o211a_1 _09297_ (.A1(net933),
    .A2(_04483_),
    .B1(_04485_),
    .C1(net495),
    .X(_01304_));
 sky130_fd_sc_hd__or2_1 _09298_ (.A(\tms1x00.O_pla_ands[2][2] ),
    .B(_04482_),
    .X(_04486_));
 sky130_fd_sc_hd__o211a_1 _09299_ (.A1(net1067),
    .A2(_04483_),
    .B1(_04486_),
    .C1(net494),
    .X(_01305_));
 sky130_fd_sc_hd__a21o_1 _09300_ (.A1(net1059),
    .A2(_04482_),
    .B1(net563),
    .X(_04487_));
 sky130_fd_sc_hd__a21o_1 _09301_ (.A1(\tms1x00.O_pla_ands[2][3] ),
    .A2(_04483_),
    .B1(_04487_),
    .X(_01306_));
 sky130_fd_sc_hd__a21o_1 _09302_ (.A1(net1051),
    .A2(_04482_),
    .B1(net559),
    .X(_04488_));
 sky130_fd_sc_hd__a21o_1 _09303_ (.A1(\tms1x00.O_pla_ands[2][4] ),
    .A2(_04483_),
    .B1(_04488_),
    .X(_01307_));
 sky130_fd_sc_hd__or2_1 _09304_ (.A(\tms1x00.O_pla_ands[2][5] ),
    .B(_04482_),
    .X(_04489_));
 sky130_fd_sc_hd__o211a_1 _09305_ (.A1(net1043),
    .A2(_04483_),
    .B1(_04489_),
    .C1(net494),
    .X(_01308_));
 sky130_fd_sc_hd__a21o_1 _09306_ (.A1(net1036),
    .A2(_04482_),
    .B1(net559),
    .X(_04490_));
 sky130_fd_sc_hd__a21o_1 _09307_ (.A1(\tms1x00.O_pla_ands[2][6] ),
    .A2(_04483_),
    .B1(_04490_),
    .X(_01309_));
 sky130_fd_sc_hd__or2_1 _09308_ (.A(\tms1x00.O_pla_ands[2][7] ),
    .B(_04482_),
    .X(_04491_));
 sky130_fd_sc_hd__o211a_1 _09309_ (.A1(net1028),
    .A2(_04483_),
    .B1(_04491_),
    .C1(net497),
    .X(_01310_));
 sky130_fd_sc_hd__or2_1 _09310_ (.A(\tms1x00.O_pla_ands[2][8] ),
    .B(_04482_),
    .X(_04492_));
 sky130_fd_sc_hd__o211a_1 _09311_ (.A1(net1019),
    .A2(_04483_),
    .B1(_04492_),
    .C1(net494),
    .X(_01311_));
 sky130_fd_sc_hd__a21o_1 _09312_ (.A1(net1012),
    .A2(_04482_),
    .B1(net559),
    .X(_04493_));
 sky130_fd_sc_hd__a21o_1 _09313_ (.A1(\tms1x00.O_pla_ands[2][9] ),
    .A2(_04483_),
    .B1(_04493_),
    .X(_01312_));
 sky130_fd_sc_hd__or3_4 _09314_ (.A(net748),
    .B(net361),
    .C(net710),
    .X(_04494_));
 sky130_fd_sc_hd__mux2_1 _09315_ (.A0(net976),
    .A1(\tms1x00.O_pla_ands[25][0] ),
    .S(_04494_),
    .X(_01313_));
 sky130_fd_sc_hd__mux2_1 _09316_ (.A0(net927),
    .A1(\tms1x00.O_pla_ands[25][1] ),
    .S(_04494_),
    .X(_01314_));
 sky130_fd_sc_hd__mux2_1 _09317_ (.A0(net1063),
    .A1(\tms1x00.O_pla_ands[25][2] ),
    .S(_04494_),
    .X(_01315_));
 sky130_fd_sc_hd__mux2_1 _09318_ (.A0(net1054),
    .A1(\tms1x00.O_pla_ands[25][3] ),
    .S(_04494_),
    .X(_01316_));
 sky130_fd_sc_hd__mux2_1 _09319_ (.A0(net1046),
    .A1(\tms1x00.O_pla_ands[25][4] ),
    .S(_04494_),
    .X(_01317_));
 sky130_fd_sc_hd__mux2_1 _09320_ (.A0(net1038),
    .A1(\tms1x00.O_pla_ands[25][5] ),
    .S(_04494_),
    .X(_01318_));
 sky130_fd_sc_hd__mux2_1 _09321_ (.A0(net1030),
    .A1(\tms1x00.O_pla_ands[25][6] ),
    .S(_04494_),
    .X(_01319_));
 sky130_fd_sc_hd__mux2_1 _09322_ (.A0(net1024),
    .A1(\tms1x00.O_pla_ands[25][7] ),
    .S(_04494_),
    .X(_01320_));
 sky130_fd_sc_hd__mux2_1 _09323_ (.A0(net1015),
    .A1(\tms1x00.O_pla_ands[25][8] ),
    .S(_04494_),
    .X(_01321_));
 sky130_fd_sc_hd__mux2_1 _09324_ (.A0(net1007),
    .A1(\tms1x00.O_pla_ands[25][9] ),
    .S(_04494_),
    .X(_01322_));
 sky130_fd_sc_hd__and3_4 _09325_ (.A(net628),
    .B(net360),
    .C(net709),
    .X(_04495_));
 sky130_fd_sc_hd__or3_4 _09326_ (.A(net622),
    .B(net357),
    .C(net707),
    .X(_04496_));
 sky130_fd_sc_hd__a21o_1 _09327_ (.A1(net981),
    .A2(_04495_),
    .B1(net560),
    .X(_04497_));
 sky130_fd_sc_hd__a21o_1 _09328_ (.A1(\tms1x00.O_pla_ands[6][0] ),
    .A2(_04496_),
    .B1(_04497_),
    .X(_01323_));
 sky130_fd_sc_hd__or2_1 _09329_ (.A(\tms1x00.O_pla_ands[6][1] ),
    .B(_04495_),
    .X(_04498_));
 sky130_fd_sc_hd__o211a_1 _09330_ (.A1(net933),
    .A2(_04496_),
    .B1(_04498_),
    .C1(net496),
    .X(_01324_));
 sky130_fd_sc_hd__or2_1 _09331_ (.A(\tms1x00.O_pla_ands[6][2] ),
    .B(_04495_),
    .X(_04499_));
 sky130_fd_sc_hd__o211a_1 _09332_ (.A1(net1067),
    .A2(_04496_),
    .B1(_04499_),
    .C1(net496),
    .X(_01325_));
 sky130_fd_sc_hd__a21o_1 _09333_ (.A1(net1059),
    .A2(_04495_),
    .B1(net558),
    .X(_04500_));
 sky130_fd_sc_hd__a21o_1 _09334_ (.A1(\tms1x00.O_pla_ands[6][3] ),
    .A2(_04496_),
    .B1(_04500_),
    .X(_01326_));
 sky130_fd_sc_hd__or2_1 _09335_ (.A(\tms1x00.O_pla_ands[6][4] ),
    .B(_04495_),
    .X(_04501_));
 sky130_fd_sc_hd__o211a_1 _09336_ (.A1(net1051),
    .A2(_04496_),
    .B1(_04501_),
    .C1(net496),
    .X(_01327_));
 sky130_fd_sc_hd__a21o_1 _09337_ (.A1(net1043),
    .A2(_04495_),
    .B1(net558),
    .X(_04502_));
 sky130_fd_sc_hd__a21o_1 _09338_ (.A1(\tms1x00.O_pla_ands[6][5] ),
    .A2(_04496_),
    .B1(_04502_),
    .X(_01328_));
 sky130_fd_sc_hd__a21o_1 _09339_ (.A1(net1036),
    .A2(_04495_),
    .B1(net558),
    .X(_04503_));
 sky130_fd_sc_hd__a21o_1 _09340_ (.A1(\tms1x00.O_pla_ands[6][6] ),
    .A2(_04496_),
    .B1(_04503_),
    .X(_01329_));
 sky130_fd_sc_hd__or2_1 _09341_ (.A(\tms1x00.O_pla_ands[6][7] ),
    .B(_04495_),
    .X(_04504_));
 sky130_fd_sc_hd__o211a_1 _09342_ (.A1(net1028),
    .A2(_04496_),
    .B1(_04504_),
    .C1(net496),
    .X(_01330_));
 sky130_fd_sc_hd__or2_1 _09343_ (.A(\tms1x00.O_pla_ands[6][8] ),
    .B(_04495_),
    .X(_04505_));
 sky130_fd_sc_hd__o211a_1 _09344_ (.A1(net1019),
    .A2(_04496_),
    .B1(_04505_),
    .C1(net496),
    .X(_01331_));
 sky130_fd_sc_hd__a21o_1 _09345_ (.A1(net1012),
    .A2(_04495_),
    .B1(net558),
    .X(_04506_));
 sky130_fd_sc_hd__a21o_1 _09346_ (.A1(\tms1x00.O_pla_ands[6][9] ),
    .A2(_04496_),
    .B1(_04506_),
    .X(_01332_));
 sky130_fd_sc_hd__or3_4 _09347_ (.A(net722),
    .B(net361),
    .C(net710),
    .X(_04507_));
 sky130_fd_sc_hd__mux2_1 _09348_ (.A0(net976),
    .A1(\tms1x00.O_pla_ands[26][0] ),
    .S(_04507_),
    .X(_01333_));
 sky130_fd_sc_hd__mux2_1 _09349_ (.A0(net927),
    .A1(\tms1x00.O_pla_ands[26][1] ),
    .S(_04507_),
    .X(_01334_));
 sky130_fd_sc_hd__mux2_1 _09350_ (.A0(net1063),
    .A1(\tms1x00.O_pla_ands[26][2] ),
    .S(_04507_),
    .X(_01335_));
 sky130_fd_sc_hd__mux2_1 _09351_ (.A0(net1054),
    .A1(\tms1x00.O_pla_ands[26][3] ),
    .S(_04507_),
    .X(_01336_));
 sky130_fd_sc_hd__mux2_1 _09352_ (.A0(net1046),
    .A1(\tms1x00.O_pla_ands[26][4] ),
    .S(_04507_),
    .X(_01337_));
 sky130_fd_sc_hd__mux2_1 _09353_ (.A0(net1038),
    .A1(\tms1x00.O_pla_ands[26][5] ),
    .S(_04507_),
    .X(_01338_));
 sky130_fd_sc_hd__mux2_1 _09354_ (.A0(net1030),
    .A1(\tms1x00.O_pla_ands[26][6] ),
    .S(_04507_),
    .X(_01339_));
 sky130_fd_sc_hd__mux2_1 _09355_ (.A0(net1024),
    .A1(\tms1x00.O_pla_ands[26][7] ),
    .S(_04507_),
    .X(_01340_));
 sky130_fd_sc_hd__mux2_1 _09356_ (.A0(net1016),
    .A1(\tms1x00.O_pla_ands[26][8] ),
    .S(_04507_),
    .X(_01341_));
 sky130_fd_sc_hd__mux2_1 _09357_ (.A0(net1007),
    .A1(\tms1x00.O_pla_ands[26][9] ),
    .S(_04507_),
    .X(_01342_));
 sky130_fd_sc_hd__and3_4 _09358_ (.A(net902),
    .B(net359),
    .C(net709),
    .X(_04508_));
 sky130_fd_sc_hd__or3_4 _09359_ (.A(net896),
    .B(net357),
    .C(net706),
    .X(_04509_));
 sky130_fd_sc_hd__or2_1 _09360_ (.A(\tms1x00.O_pla_ands[5][0] ),
    .B(_04508_),
    .X(_04510_));
 sky130_fd_sc_hd__o211a_1 _09361_ (.A1(net981),
    .A2(_04509_),
    .B1(_04510_),
    .C1(net494),
    .X(_01343_));
 sky130_fd_sc_hd__a21o_1 _09362_ (.A1(net933),
    .A2(_04508_),
    .B1(net559),
    .X(_04511_));
 sky130_fd_sc_hd__a21o_1 _09363_ (.A1(\tms1x00.O_pla_ands[5][1] ),
    .A2(_04509_),
    .B1(_04511_),
    .X(_01344_));
 sky130_fd_sc_hd__a21o_1 _09364_ (.A1(net1067),
    .A2(_04508_),
    .B1(net532),
    .X(_04512_));
 sky130_fd_sc_hd__a21o_1 _09365_ (.A1(\tms1x00.O_pla_ands[5][2] ),
    .A2(_04509_),
    .B1(_04512_),
    .X(_01345_));
 sky130_fd_sc_hd__or2_1 _09366_ (.A(\tms1x00.O_pla_ands[5][3] ),
    .B(_04508_),
    .X(_04513_));
 sky130_fd_sc_hd__o211a_1 _09367_ (.A1(net1059),
    .A2(_04509_),
    .B1(_04513_),
    .C1(net495),
    .X(_01346_));
 sky130_fd_sc_hd__or2_1 _09368_ (.A(\tms1x00.O_pla_ands[5][4] ),
    .B(_04508_),
    .X(_04514_));
 sky130_fd_sc_hd__o211a_1 _09369_ (.A1(net1051),
    .A2(_04509_),
    .B1(_04514_),
    .C1(net494),
    .X(_01347_));
 sky130_fd_sc_hd__a21o_1 _09370_ (.A1(net1043),
    .A2(_04508_),
    .B1(net559),
    .X(_04515_));
 sky130_fd_sc_hd__a21o_1 _09371_ (.A1(\tms1x00.O_pla_ands[5][5] ),
    .A2(_04509_),
    .B1(_04515_),
    .X(_01348_));
 sky130_fd_sc_hd__a21o_1 _09372_ (.A1(net1036),
    .A2(_04508_),
    .B1(net559),
    .X(_04516_));
 sky130_fd_sc_hd__a21o_1 _09373_ (.A1(\tms1x00.O_pla_ands[5][6] ),
    .A2(_04509_),
    .B1(_04516_),
    .X(_01349_));
 sky130_fd_sc_hd__or2_1 _09374_ (.A(\tms1x00.O_pla_ands[5][7] ),
    .B(_04508_),
    .X(_04517_));
 sky130_fd_sc_hd__o211a_1 _09375_ (.A1(net1028),
    .A2(_04509_),
    .B1(_04517_),
    .C1(net494),
    .X(_01350_));
 sky130_fd_sc_hd__or2_1 _09376_ (.A(\tms1x00.O_pla_ands[5][8] ),
    .B(_04508_),
    .X(_04518_));
 sky130_fd_sc_hd__o211a_1 _09377_ (.A1(net1019),
    .A2(_04509_),
    .B1(_04518_),
    .C1(net494),
    .X(_01351_));
 sky130_fd_sc_hd__a21o_1 _09378_ (.A1(net1009),
    .A2(_04508_),
    .B1(net532),
    .X(_04519_));
 sky130_fd_sc_hd__a21o_1 _09379_ (.A1(\tms1x00.O_pla_ands[5][9] ),
    .A2(_04509_),
    .B1(_04519_),
    .X(_01352_));
 sky130_fd_sc_hd__or3_4 _09380_ (.A(net776),
    .B(net361),
    .C(_03353_),
    .X(_04520_));
 sky130_fd_sc_hd__mux2_1 _09381_ (.A0(net976),
    .A1(\tms1x00.O_pla_ands[23][0] ),
    .S(_04520_),
    .X(_01353_));
 sky130_fd_sc_hd__mux2_1 _09382_ (.A0(net927),
    .A1(\tms1x00.O_pla_ands[23][1] ),
    .S(_04520_),
    .X(_01354_));
 sky130_fd_sc_hd__mux2_1 _09383_ (.A0(net1064),
    .A1(\tms1x00.O_pla_ands[23][2] ),
    .S(_04520_),
    .X(_01355_));
 sky130_fd_sc_hd__mux2_1 _09384_ (.A0(net1055),
    .A1(\tms1x00.O_pla_ands[23][3] ),
    .S(_04520_),
    .X(_01356_));
 sky130_fd_sc_hd__mux2_1 _09385_ (.A0(net1046),
    .A1(\tms1x00.O_pla_ands[23][4] ),
    .S(_04520_),
    .X(_01357_));
 sky130_fd_sc_hd__mux2_1 _09386_ (.A0(net1038),
    .A1(\tms1x00.O_pla_ands[23][5] ),
    .S(_04520_),
    .X(_01358_));
 sky130_fd_sc_hd__mux2_1 _09387_ (.A0(net1030),
    .A1(\tms1x00.O_pla_ands[23][6] ),
    .S(_04520_),
    .X(_01359_));
 sky130_fd_sc_hd__mux2_1 _09388_ (.A0(net1024),
    .A1(\tms1x00.O_pla_ands[23][7] ),
    .S(_04520_),
    .X(_01360_));
 sky130_fd_sc_hd__mux2_1 _09389_ (.A0(net1017),
    .A1(\tms1x00.O_pla_ands[23][8] ),
    .S(_04520_),
    .X(_01361_));
 sky130_fd_sc_hd__mux2_1 _09390_ (.A0(net1007),
    .A1(\tms1x00.O_pla_ands[23][9] ),
    .S(_04520_),
    .X(_01362_));
 sky130_fd_sc_hd__or3_4 _09391_ (.A(net610),
    .B(_03351_),
    .C(_03353_),
    .X(_04521_));
 sky130_fd_sc_hd__mux2_1 _09392_ (.A0(net976),
    .A1(\tms1x00.O_pla_ands[22][0] ),
    .S(_04521_),
    .X(_01363_));
 sky130_fd_sc_hd__mux2_1 _09393_ (.A0(net928),
    .A1(\tms1x00.O_pla_ands[22][1] ),
    .S(_04521_),
    .X(_01364_));
 sky130_fd_sc_hd__mux2_1 _09394_ (.A0(net1064),
    .A1(\tms1x00.O_pla_ands[22][2] ),
    .S(_04521_),
    .X(_01365_));
 sky130_fd_sc_hd__mux2_1 _09395_ (.A0(net1055),
    .A1(\tms1x00.O_pla_ands[22][3] ),
    .S(_04521_),
    .X(_01366_));
 sky130_fd_sc_hd__mux2_1 _09396_ (.A0(net1047),
    .A1(\tms1x00.O_pla_ands[22][4] ),
    .S(_04521_),
    .X(_01367_));
 sky130_fd_sc_hd__mux2_1 _09397_ (.A0(net1039),
    .A1(\tms1x00.O_pla_ands[22][5] ),
    .S(_04521_),
    .X(_01368_));
 sky130_fd_sc_hd__mux2_1 _09398_ (.A0(net1030),
    .A1(\tms1x00.O_pla_ands[22][6] ),
    .S(_04521_),
    .X(_01369_));
 sky130_fd_sc_hd__mux2_1 _09399_ (.A0(net1024),
    .A1(\tms1x00.O_pla_ands[22][7] ),
    .S(_04521_),
    .X(_01370_));
 sky130_fd_sc_hd__mux2_1 _09400_ (.A0(net1017),
    .A1(\tms1x00.O_pla_ands[22][8] ),
    .S(_04521_),
    .X(_01371_));
 sky130_fd_sc_hd__mux2_1 _09401_ (.A0(net1008),
    .A1(\tms1x00.O_pla_ands[22][9] ),
    .S(_04521_),
    .X(_01372_));
 sky130_fd_sc_hd__and2_1 _09402_ (.A(\tms1x00.wb_step ),
    .B(net637),
    .X(_01373_));
 sky130_fd_sc_hd__nand2b_2 _09403_ (.A_N(\tms1x00.cycle[1] ),
    .B(\tms1x00.cycle[2] ),
    .Y(_04522_));
 sky130_fd_sc_hd__nor2_4 _09404_ (.A(\tms1x00.cycle[0] ),
    .B(net593),
    .Y(_04523_));
 sky130_fd_sc_hd__or2_4 _09405_ (.A(\tms1x00.cycle[0] ),
    .B(net593),
    .X(_04524_));
 sky130_fd_sc_hd__nor2_8 _09406_ (.A(net458),
    .B(_04524_),
    .Y(_04525_));
 sky130_fd_sc_hd__nand2_8 _09407_ (.A(net631),
    .B(_04525_),
    .Y(_04526_));
 sky130_fd_sc_hd__mux2_1 _09408_ (.A0(\tms1x00.Y[0] ),
    .A1(net146),
    .S(_04526_),
    .X(_01374_));
 sky130_fd_sc_hd__mux2_1 _09409_ (.A0(\tms1x00.Y[1] ),
    .A1(net147),
    .S(_04526_),
    .X(_01375_));
 sky130_fd_sc_hd__mux2_1 _09410_ (.A0(net654),
    .A1(net148),
    .S(_04526_),
    .X(_01376_));
 sky130_fd_sc_hd__mux2_1 _09411_ (.A0(net652),
    .A1(net149),
    .S(_04526_),
    .X(_01377_));
 sky130_fd_sc_hd__mux2_1 _09412_ (.A0(\tms1x00.X[0] ),
    .A1(net150),
    .S(_04526_),
    .X(_01378_));
 sky130_fd_sc_hd__mux2_1 _09413_ (.A0(\tms1x00.X[1] ),
    .A1(net151),
    .S(_04526_),
    .X(_01379_));
 sky130_fd_sc_hd__mux2_1 _09414_ (.A0(\tms1x00.X[2] ),
    .A1(net152),
    .S(_04526_),
    .X(_01380_));
 sky130_fd_sc_hd__nor2_2 _09415_ (.A(\tms1x00.cycle[2] ),
    .B(\tms1x00.cycle[1] ),
    .Y(_04527_));
 sky130_fd_sc_hd__nand2_4 _09416_ (.A(_03374_),
    .B(_04527_),
    .Y(_04528_));
 sky130_fd_sc_hd__mux2_1 _09417_ (.A0(\tms1x00.PC[0] ),
    .A1(\tms1x00.rom_addr[0] ),
    .S(net339),
    .X(_01381_));
 sky130_fd_sc_hd__mux2_1 _09418_ (.A0(\tms1x00.PC[1] ),
    .A1(\tms1x00.rom_addr[1] ),
    .S(_04528_),
    .X(_01382_));
 sky130_fd_sc_hd__mux2_1 _09419_ (.A0(\tms1x00.PC[2] ),
    .A1(net158),
    .S(net339),
    .X(_01383_));
 sky130_fd_sc_hd__mux2_1 _09420_ (.A0(\tms1x00.PC[3] ),
    .A1(net159),
    .S(net339),
    .X(_01384_));
 sky130_fd_sc_hd__mux2_1 _09421_ (.A0(\tms1x00.PC[4] ),
    .A1(net160),
    .S(net339),
    .X(_01385_));
 sky130_fd_sc_hd__mux2_1 _09422_ (.A0(\tms1x00.PC[5] ),
    .A1(net161),
    .S(net339),
    .X(_01386_));
 sky130_fd_sc_hd__mux2_1 _09423_ (.A0(\tms1x00.PA[0] ),
    .A1(net162),
    .S(net339),
    .X(_01387_));
 sky130_fd_sc_hd__mux2_1 _09424_ (.A0(\tms1x00.PA[1] ),
    .A1(net163),
    .S(net339),
    .X(_01388_));
 sky130_fd_sc_hd__mux2_1 _09425_ (.A0(\tms1x00.PA[2] ),
    .A1(net164),
    .S(net339),
    .X(_01389_));
 sky130_fd_sc_hd__mux2_1 _09426_ (.A0(\tms1x00.PA[3] ),
    .A1(net165),
    .S(_04528_),
    .X(_01390_));
 sky130_fd_sc_hd__mux2_1 _09427_ (.A0(\tms1x00.CA ),
    .A1(net166),
    .S(net339),
    .X(_01391_));
 sky130_fd_sc_hd__mux2_1 _09428_ (.A0(net1),
    .A1(chip_sel_override),
    .S(net145),
    .X(_04529_));
 sky130_fd_sc_hd__mux2_1 _09429_ (.A0(net705),
    .A1(_04529_),
    .S(net591),
    .X(_01392_));
 sky130_fd_sc_hd__nand2_8 _09430_ (.A(\tms1x00.status ),
    .B(net669),
    .Y(_04530_));
 sky130_fd_sc_hd__or4_1 _09431_ (.A(_01622_),
    .B(_01624_),
    .C(net593),
    .D(_04530_),
    .X(_04531_));
 sky130_fd_sc_hd__or2_4 _09432_ (.A(net458),
    .B(_04531_),
    .X(_04532_));
 sky130_fd_sc_hd__nor2_1 _09433_ (.A(\tms1x00.CL ),
    .B(_04532_),
    .Y(_04533_));
 sky130_fd_sc_hd__and2_4 _09434_ (.A(net633),
    .B(_04533_),
    .X(_04534_));
 sky130_fd_sc_hd__mux2_1 _09435_ (.A0(\tms1x00.SR[0] ),
    .A1(\tms1x00.PC[0] ),
    .S(_04534_),
    .X(_01393_));
 sky130_fd_sc_hd__mux2_1 _09436_ (.A0(\tms1x00.SR[1] ),
    .A1(\tms1x00.PC[1] ),
    .S(_04534_),
    .X(_01394_));
 sky130_fd_sc_hd__mux2_1 _09437_ (.A0(\tms1x00.SR[2] ),
    .A1(\tms1x00.PC[2] ),
    .S(_04534_),
    .X(_01395_));
 sky130_fd_sc_hd__mux2_1 _09438_ (.A0(\tms1x00.SR[3] ),
    .A1(\tms1x00.PC[3] ),
    .S(_04534_),
    .X(_01396_));
 sky130_fd_sc_hd__mux2_1 _09439_ (.A0(\tms1x00.SR[4] ),
    .A1(\tms1x00.PC[4] ),
    .S(_04534_),
    .X(_01397_));
 sky130_fd_sc_hd__mux2_1 _09440_ (.A0(\tms1x00.SR[5] ),
    .A1(\tms1x00.PC[5] ),
    .S(_04534_),
    .X(_01398_));
 sky130_fd_sc_hd__nor2_2 _09441_ (.A(_01639_),
    .B(_01640_),
    .Y(_04535_));
 sky130_fd_sc_hd__or2_2 _09442_ (.A(\tms1x00.rom_addr[0] ),
    .B(\tms1x00.rom_addr[1] ),
    .X(_04536_));
 sky130_fd_sc_hd__mux4_1 _09443_ (.A0(net10),
    .A1(net40),
    .A2(net17),
    .A3(net26),
    .S0(\tms1x00.rom_addr[0] ),
    .S1(\tms1x00.rom_addr[1] ),
    .X(_04537_));
 sky130_fd_sc_hd__nand2_1 _09444_ (.A(_01630_),
    .B(net632),
    .Y(_04538_));
 sky130_fd_sc_hd__a22o_1 _09445_ (.A1(_04525_),
    .A2(_04537_),
    .B1(_04538_),
    .B2(_04526_),
    .X(_01399_));
 sky130_fd_sc_hd__mux4_1 _09446_ (.A0(net21),
    .A1(net41),
    .A2(net18),
    .A3(net27),
    .S0(\tms1x00.rom_addr[0] ),
    .S1(\tms1x00.rom_addr[1] ),
    .X(_04539_));
 sky130_fd_sc_hd__nand2_2 _09447_ (.A(_01629_),
    .B(net637),
    .Y(_04540_));
 sky130_fd_sc_hd__a22o_1 _09448_ (.A1(_04525_),
    .A2(_04539_),
    .B1(_04540_),
    .B2(_04526_),
    .X(_01400_));
 sky130_fd_sc_hd__o21a_1 _09449_ (.A1(_01640_),
    .A2(net19),
    .B1(_01639_),
    .X(_04541_));
 sky130_fd_sc_hd__a221o_1 _09450_ (.A1(_01640_),
    .A2(net11),
    .B1(_04535_),
    .B2(net28),
    .C1(_04541_),
    .X(_04542_));
 sky130_fd_sc_hd__o21ai_1 _09451_ (.A1(net32),
    .A2(_04536_),
    .B1(_04542_),
    .Y(_04543_));
 sky130_fd_sc_hd__nand2_1 _09452_ (.A(net362),
    .B(_04543_),
    .Y(_04544_));
 sky130_fd_sc_hd__o211a_1 _09453_ (.A1(net692),
    .A2(net362),
    .B1(_04544_),
    .C1(net631),
    .X(_01401_));
 sky130_fd_sc_hd__o21a_1 _09454_ (.A1(_01640_),
    .A2(net20),
    .B1(_01639_),
    .X(_04545_));
 sky130_fd_sc_hd__a221o_1 _09455_ (.A1(_01640_),
    .A2(net12),
    .B1(_04535_),
    .B2(net29),
    .C1(_04545_),
    .X(_04546_));
 sky130_fd_sc_hd__o21ai_1 _09456_ (.A1(net35),
    .A2(_04536_),
    .B1(_04546_),
    .Y(_04547_));
 sky130_fd_sc_hd__nand2_1 _09457_ (.A(net362),
    .B(_04547_),
    .Y(_04548_));
 sky130_fd_sc_hd__o211a_1 _09458_ (.A1(net686),
    .A2(net362),
    .B1(_04548_),
    .C1(net631),
    .X(_01402_));
 sky130_fd_sc_hd__o21a_1 _09459_ (.A1(_01639_),
    .A2(net13),
    .B1(_01640_),
    .X(_04549_));
 sky130_fd_sc_hd__a221o_1 _09460_ (.A1(_01639_),
    .A2(net22),
    .B1(_04535_),
    .B2(net30),
    .C1(_04549_),
    .X(_04550_));
 sky130_fd_sc_hd__o21ai_1 _09461_ (.A1(net36),
    .A2(_04536_),
    .B1(_04550_),
    .Y(_04551_));
 sky130_fd_sc_hd__nand2_1 _09462_ (.A(net362),
    .B(_04551_),
    .Y(_04552_));
 sky130_fd_sc_hd__o211a_1 _09463_ (.A1(net682),
    .A2(net362),
    .B1(_04552_),
    .C1(net631),
    .X(_01403_));
 sky130_fd_sc_hd__mux4_1 _09464_ (.A0(net37),
    .A1(net14),
    .A2(net23),
    .A3(net31),
    .S0(\tms1x00.rom_addr[0] ),
    .S1(\tms1x00.rom_addr[1] ),
    .X(_04553_));
 sky130_fd_sc_hd__nand2_1 _09465_ (.A(_01625_),
    .B(net632),
    .Y(_04554_));
 sky130_fd_sc_hd__a22o_1 _09466_ (.A1(net362),
    .A2(_04553_),
    .B1(_04554_),
    .B2(_04526_),
    .X(_01404_));
 sky130_fd_sc_hd__o21a_1 _09467_ (.A1(_01639_),
    .A2(net15),
    .B1(_01640_),
    .X(_04555_));
 sky130_fd_sc_hd__a221o_1 _09468_ (.A1(_01639_),
    .A2(net24),
    .B1(_04535_),
    .B2(net33),
    .C1(_04555_),
    .X(_04556_));
 sky130_fd_sc_hd__o21ai_1 _09469_ (.A1(net38),
    .A2(_04536_),
    .B1(_04556_),
    .Y(_04557_));
 sky130_fd_sc_hd__nand2_1 _09470_ (.A(net362),
    .B(_04557_),
    .Y(_04558_));
 sky130_fd_sc_hd__o211a_1 _09471_ (.A1(net672),
    .A2(net362),
    .B1(_04558_),
    .C1(net632),
    .X(_01405_));
 sky130_fd_sc_hd__o21a_1 _09472_ (.A1(_01640_),
    .A2(net25),
    .B1(_01639_),
    .X(_04559_));
 sky130_fd_sc_hd__a221o_1 _09473_ (.A1(_01640_),
    .A2(net16),
    .B1(_04535_),
    .B2(net34),
    .C1(_04559_),
    .X(_04560_));
 sky130_fd_sc_hd__o21ai_1 _09474_ (.A1(net39),
    .A2(_04536_),
    .B1(_04560_),
    .Y(_04561_));
 sky130_fd_sc_hd__nand2_1 _09475_ (.A(net362),
    .B(_04561_),
    .Y(_04562_));
 sky130_fd_sc_hd__o211a_1 _09476_ (.A1(net668),
    .A2(_04525_),
    .B1(_04562_),
    .C1(net632),
    .X(_01406_));
 sky130_fd_sc_hd__nand2_1 _09477_ (.A(_01622_),
    .B(net458),
    .Y(_04563_));
 sky130_fd_sc_hd__and3_1 _09478_ (.A(net632),
    .B(_04305_),
    .C(_04563_),
    .X(_01407_));
 sky130_fd_sc_hd__a21o_1 _09479_ (.A1(\tms1x00.cycle[0] ),
    .A2(_03373_),
    .B1(\tms1x00.cycle[1] ),
    .X(_04564_));
 sky130_fd_sc_hd__o211a_1 _09480_ (.A1(_04305_),
    .A2(_04527_),
    .B1(_04564_),
    .C1(net633),
    .X(_01408_));
 sky130_fd_sc_hd__nand2_1 _09481_ (.A(\tms1x00.cycle[2] ),
    .B(_04305_),
    .Y(_04565_));
 sky130_fd_sc_hd__a21oi_1 _09482_ (.A1(_04306_),
    .A2(_04565_),
    .B1(net592),
    .Y(_01409_));
 sky130_fd_sc_hd__nand2b_1 _09483_ (.A_N(net655),
    .B(net656),
    .Y(_04566_));
 sky130_fd_sc_hd__nor2_1 _09484_ (.A(net655),
    .B(net656),
    .Y(_04567_));
 sky130_fd_sc_hd__and2b_1 _09485_ (.A_N(net653),
    .B(_04567_),
    .X(_04568_));
 sky130_fd_sc_hd__or3_1 _09486_ (.A(net653),
    .B(net655),
    .C(net656),
    .X(_04569_));
 sky130_fd_sc_hd__nor2_1 _09487_ (.A(net653),
    .B(_04566_),
    .Y(_04570_));
 sky130_fd_sc_hd__nor4_4 _09488_ (.A(_03376_),
    .B(_03378_),
    .C(_03394_),
    .D(net340),
    .Y(_04571_));
 sky130_fd_sc_hd__nand3_1 _09489_ (.A(net648),
    .B(_04570_),
    .C(net242),
    .Y(_04572_));
 sky130_fd_sc_hd__inv_2 _09490_ (.A(_04572_),
    .Y(_04573_));
 sky130_fd_sc_hd__or3_4 _09491_ (.A(_03376_),
    .B(net340),
    .C(_04310_),
    .X(_04574_));
 sky130_fd_sc_hd__or3b_1 _09492_ (.A(net240),
    .B(net650),
    .C_N(_04570_),
    .X(_04575_));
 sky130_fd_sc_hd__o211a_1 _09493_ (.A1(net129),
    .A2(_04573_),
    .B1(_04575_),
    .C1(net635),
    .X(_01410_));
 sky130_fd_sc_hd__nor3b_2 _09494_ (.A(net654),
    .B(net656),
    .C_N(net655),
    .Y(_04576_));
 sky130_fd_sc_hd__nand3_1 _09495_ (.A(net649),
    .B(net243),
    .C(_04576_),
    .Y(_04577_));
 sky130_fd_sc_hd__inv_2 _09496_ (.A(_04577_),
    .Y(_04578_));
 sky130_fd_sc_hd__or3b_1 _09497_ (.A(net651),
    .B(net241),
    .C_N(_04576_),
    .X(_04579_));
 sky130_fd_sc_hd__o211a_1 _09498_ (.A1(net130),
    .A2(_04578_),
    .B1(_04579_),
    .C1(net636),
    .X(_01411_));
 sky130_fd_sc_hd__and3b_1 _09499_ (.A_N(net654),
    .B(net655),
    .C(net656),
    .X(_04580_));
 sky130_fd_sc_hd__nand3_1 _09500_ (.A(net649),
    .B(net243),
    .C(_04580_),
    .Y(_04581_));
 sky130_fd_sc_hd__inv_2 _09501_ (.A(_04581_),
    .Y(_04582_));
 sky130_fd_sc_hd__or3b_1 _09502_ (.A(net652),
    .B(net241),
    .C_N(_04580_),
    .X(_04583_));
 sky130_fd_sc_hd__o211a_1 _09503_ (.A1(net131),
    .A2(_04582_),
    .B1(_04583_),
    .C1(net635),
    .X(_01412_));
 sky130_fd_sc_hd__nand2_1 _09504_ (.A(net653),
    .B(_04567_),
    .Y(_04584_));
 sky130_fd_sc_hd__a41o_1 _09505_ (.A1(net648),
    .A2(net653),
    .A3(_04567_),
    .A4(net242),
    .B1(net132),
    .X(_04585_));
 sky130_fd_sc_hd__o311a_1 _09506_ (.A1(net650),
    .A2(net240),
    .A3(_04584_),
    .B1(_04585_),
    .C1(net634),
    .X(_01413_));
 sky130_fd_sc_hd__and3b_1 _09507_ (.A_N(net655),
    .B(net656),
    .C(net654),
    .X(_04586_));
 sky130_fd_sc_hd__inv_2 _09508_ (.A(_04586_),
    .Y(_04587_));
 sky130_fd_sc_hd__a31o_1 _09509_ (.A1(net649),
    .A2(net243),
    .A3(_04586_),
    .B1(net133),
    .X(_04588_));
 sky130_fd_sc_hd__o311a_1 _09510_ (.A1(net650),
    .A2(net241),
    .A3(_04587_),
    .B1(_04588_),
    .C1(net635),
    .X(_01414_));
 sky130_fd_sc_hd__and3b_1 _09511_ (.A_N(net656),
    .B(net655),
    .C(net654),
    .X(_04589_));
 sky130_fd_sc_hd__inv_2 _09512_ (.A(_04589_),
    .Y(_04590_));
 sky130_fd_sc_hd__a31o_1 _09513_ (.A1(net648),
    .A2(net243),
    .A3(_04589_),
    .B1(net134),
    .X(_04591_));
 sky130_fd_sc_hd__o311a_1 _09514_ (.A1(net650),
    .A2(net241),
    .A3(_04590_),
    .B1(_04591_),
    .C1(net635),
    .X(_01415_));
 sky130_fd_sc_hd__and3_1 _09515_ (.A(net653),
    .B(net655),
    .C(net656),
    .X(_04592_));
 sky130_fd_sc_hd__inv_2 _09516_ (.A(_04592_),
    .Y(_04593_));
 sky130_fd_sc_hd__a31o_1 _09517_ (.A1(net648),
    .A2(net242),
    .A3(_04592_),
    .B1(net135),
    .X(_04594_));
 sky130_fd_sc_hd__o311a_1 _09518_ (.A1(net650),
    .A2(net240),
    .A3(_04593_),
    .B1(_04594_),
    .C1(net634),
    .X(_01416_));
 sky130_fd_sc_hd__a31o_1 _09519_ (.A1(net651),
    .A2(_04568_),
    .A3(net242),
    .B1(net136),
    .X(_04595_));
 sky130_fd_sc_hd__o311a_1 _09520_ (.A1(net648),
    .A2(_04569_),
    .A3(net240),
    .B1(_04595_),
    .C1(net635),
    .X(_01417_));
 sky130_fd_sc_hd__a31o_1 _09521_ (.A1(net650),
    .A2(_04570_),
    .A3(net242),
    .B1(net137),
    .X(_04596_));
 sky130_fd_sc_hd__or4_1 _09522_ (.A(net648),
    .B(net653),
    .C(_04566_),
    .D(net240),
    .X(_04597_));
 sky130_fd_sc_hd__and3_1 _09523_ (.A(net634),
    .B(_04596_),
    .C(_04597_),
    .X(_01418_));
 sky130_fd_sc_hd__a31o_1 _09524_ (.A1(net652),
    .A2(net242),
    .A3(_04576_),
    .B1(net138),
    .X(_04598_));
 sky130_fd_sc_hd__or3b_1 _09525_ (.A(net648),
    .B(net240),
    .C_N(_04576_),
    .X(_04599_));
 sky130_fd_sc_hd__and3_1 _09526_ (.A(net635),
    .B(_04598_),
    .C(_04599_),
    .X(_01419_));
 sky130_fd_sc_hd__a31o_1 _09527_ (.A1(net652),
    .A2(net242),
    .A3(_04580_),
    .B1(net139),
    .X(_04600_));
 sky130_fd_sc_hd__or3b_1 _09528_ (.A(net649),
    .B(net240),
    .C_N(_04580_),
    .X(_04601_));
 sky130_fd_sc_hd__and3_1 _09529_ (.A(net635),
    .B(_04600_),
    .C(_04601_),
    .X(_01420_));
 sky130_fd_sc_hd__a41o_1 _09530_ (.A1(net650),
    .A2(net653),
    .A3(_04567_),
    .A4(net242),
    .B1(net140),
    .X(_04602_));
 sky130_fd_sc_hd__o311a_1 _09531_ (.A1(net648),
    .A2(net240),
    .A3(_04584_),
    .B1(_04602_),
    .C1(net634),
    .X(_01421_));
 sky130_fd_sc_hd__a31o_1 _09532_ (.A1(net650),
    .A2(net243),
    .A3(_04586_),
    .B1(net141),
    .X(_04603_));
 sky130_fd_sc_hd__o311a_1 _09533_ (.A1(net649),
    .A2(net241),
    .A3(_04587_),
    .B1(_04603_),
    .C1(net635),
    .X(_01422_));
 sky130_fd_sc_hd__a31o_1 _09534_ (.A1(net650),
    .A2(net243),
    .A3(_04589_),
    .B1(net142),
    .X(_04604_));
 sky130_fd_sc_hd__o311a_1 _09535_ (.A1(net649),
    .A2(net241),
    .A3(_04590_),
    .B1(_04604_),
    .C1(net635),
    .X(_01423_));
 sky130_fd_sc_hd__a31o_1 _09536_ (.A1(net650),
    .A2(net242),
    .A3(_04592_),
    .B1(net143),
    .X(_04605_));
 sky130_fd_sc_hd__o311a_1 _09537_ (.A1(net648),
    .A2(net240),
    .A3(_04593_),
    .B1(_04605_),
    .C1(net634),
    .X(_01424_));
 sky130_fd_sc_hd__and4_2 _09538_ (.A(net688),
    .B(_01628_),
    .C(_03377_),
    .D(_03388_),
    .X(_04606_));
 sky130_fd_sc_hd__or4_4 _09539_ (.A(_01629_),
    .B(net702),
    .C(_03378_),
    .D(_04303_),
    .X(_04607_));
 sky130_fd_sc_hd__or4_4 _09540_ (.A(net705),
    .B(_03378_),
    .C(_03400_),
    .D(_04303_),
    .X(_04608_));
 sky130_fd_sc_hd__a21oi_4 _09541_ (.A1(_04607_),
    .A2(_04608_),
    .B1(net340),
    .Y(_04609_));
 sky130_fd_sc_hd__a21o_2 _09542_ (.A1(_04607_),
    .A2(_04608_),
    .B1(net340),
    .X(_04610_));
 sky130_fd_sc_hd__a21o_1 _09543_ (.A1(\tms1x00.A[0] ),
    .A2(_04606_),
    .B1(_04610_),
    .X(_04611_));
 sky130_fd_sc_hd__o211a_1 _09544_ (.A1(\tms1x00.O_latch[0] ),
    .A2(_04609_),
    .B1(_04611_),
    .C1(net636),
    .X(_01425_));
 sky130_fd_sc_hd__a21o_1 _09545_ (.A1(\tms1x00.A[1] ),
    .A2(_04606_),
    .B1(_04610_),
    .X(_04612_));
 sky130_fd_sc_hd__o211a_1 _09546_ (.A1(net664),
    .A2(_04609_),
    .B1(_04612_),
    .C1(net636),
    .X(_01426_));
 sky130_fd_sc_hd__a21o_1 _09547_ (.A1(\tms1x00.A[2] ),
    .A2(_04606_),
    .B1(_04610_),
    .X(_04613_));
 sky130_fd_sc_hd__o211a_1 _09548_ (.A1(net661),
    .A2(_04609_),
    .B1(_04613_),
    .C1(net636),
    .X(_01427_));
 sky130_fd_sc_hd__a21o_1 _09549_ (.A1(\tms1x00.A[3] ),
    .A2(_04606_),
    .B1(_04610_),
    .X(_04614_));
 sky130_fd_sc_hd__o211a_1 _09550_ (.A1(net660),
    .A2(_04609_),
    .B1(_04614_),
    .C1(net636),
    .X(_01428_));
 sky130_fd_sc_hd__a21o_1 _09551_ (.A1(\tms1x00.SL ),
    .A2(_04606_),
    .B1(_04610_),
    .X(_04615_));
 sky130_fd_sc_hd__o211a_1 _09552_ (.A1(net658),
    .A2(_04609_),
    .B1(_04615_),
    .C1(net637),
    .X(_01429_));
 sky130_fd_sc_hd__nor3_4 _09553_ (.A(_03376_),
    .B(_03378_),
    .C(_03400_),
    .Y(_04616_));
 sky130_fd_sc_hd__nor2_4 _09554_ (.A(_04305_),
    .B(net593),
    .Y(_04617_));
 sky130_fd_sc_hd__a221oi_1 _09555_ (.A1(_01616_),
    .A2(_04532_),
    .B1(_04616_),
    .B2(_04617_),
    .C1(net592),
    .Y(_01430_));
 sky130_fd_sc_hd__nand2_1 _09556_ (.A(\tms1x00.P[3] ),
    .B(\tms1x00.N[3] ),
    .Y(_04618_));
 sky130_fd_sc_hd__or2_1 _09557_ (.A(\tms1x00.P[3] ),
    .B(\tms1x00.N[3] ),
    .X(_04619_));
 sky130_fd_sc_hd__nand2_2 _09558_ (.A(_04618_),
    .B(_04619_),
    .Y(_04620_));
 sky130_fd_sc_hd__and2_2 _09559_ (.A(\tms1x00.N[2] ),
    .B(\tms1x00.P[2] ),
    .X(_04621_));
 sky130_fd_sc_hd__nor2_2 _09560_ (.A(\tms1x00.N[2] ),
    .B(\tms1x00.P[2] ),
    .Y(_04622_));
 sky130_fd_sc_hd__nor2_2 _09561_ (.A(_04621_),
    .B(_04622_),
    .Y(_04623_));
 sky130_fd_sc_hd__and2_2 _09562_ (.A(\tms1x00.N[1] ),
    .B(\tms1x00.P[1] ),
    .X(_04624_));
 sky130_fd_sc_hd__nor2_1 _09563_ (.A(\tms1x00.N[1] ),
    .B(\tms1x00.P[1] ),
    .Y(_04625_));
 sky130_fd_sc_hd__nor2_4 _09564_ (.A(_04624_),
    .B(_04625_),
    .Y(_04626_));
 sky130_fd_sc_hd__or4_1 _09565_ (.A(net444),
    .B(net424),
    .C(net409),
    .D(net407),
    .X(_04627_));
 sky130_fd_sc_hd__or4_1 _09566_ (.A(net440),
    .B(net438),
    .C(net432),
    .D(net422),
    .X(_04628_));
 sky130_fd_sc_hd__or4_1 _09567_ (.A(net454),
    .B(net430),
    .C(net415),
    .D(net411),
    .X(_04629_));
 sky130_fd_sc_hd__or4_1 _09568_ (.A(net446),
    .B(net442),
    .C(net436),
    .D(net434),
    .X(_04630_));
 sky130_fd_sc_hd__or4_4 _09569_ (.A(_04627_),
    .B(_04628_),
    .C(_04629_),
    .D(_04630_),
    .X(_04631_));
 sky130_fd_sc_hd__or2_1 _09570_ (.A(net452),
    .B(net412),
    .X(_04632_));
 sky130_fd_sc_hd__or4_1 _09571_ (.A(net456),
    .B(net450),
    .C(net416),
    .D(net402),
    .X(_04633_));
 sky130_fd_sc_hd__or4_1 _09572_ (.A(net429),
    .B(net426),
    .C(net404),
    .D(net398),
    .X(_04634_));
 sky130_fd_sc_hd__or4_1 _09573_ (.A(net449),
    .B(net420),
    .C(net418),
    .D(net400),
    .X(_04635_));
 sky130_fd_sc_hd__or4_4 _09574_ (.A(_04632_),
    .B(_04633_),
    .C(_04634_),
    .D(_04635_),
    .X(_04636_));
 sky130_fd_sc_hd__nor2_8 _09575_ (.A(_04631_),
    .B(_04636_),
    .Y(_04637_));
 sky130_fd_sc_hd__or2_1 _09576_ (.A(_04631_),
    .B(_04636_),
    .X(_04638_));
 sky130_fd_sc_hd__a22o_1 _09577_ (.A1(\tms1x00.ins_pla_ors[12][28] ),
    .A2(net446),
    .B1(net428),
    .B2(\tms1x00.ins_pla_ors[12][29] ),
    .X(_04639_));
 sky130_fd_sc_hd__a22o_1 _09578_ (.A1(\tms1x00.ins_pla_ors[12][4] ),
    .A2(net442),
    .B1(net402),
    .B2(\tms1x00.ins_pla_ors[12][5] ),
    .X(_04640_));
 sky130_fd_sc_hd__a22o_1 _09579_ (.A1(\tms1x00.ins_pla_ors[12][7] ),
    .A2(net450),
    .B1(net400),
    .B2(\tms1x00.ins_pla_ors[12][6] ),
    .X(_04641_));
 sky130_fd_sc_hd__a22o_1 _09580_ (.A1(\tms1x00.ins_pla_ors[12][2] ),
    .A2(net438),
    .B1(net432),
    .B2(\tms1x00.ins_pla_ors[12][3] ),
    .X(_04642_));
 sky130_fd_sc_hd__a221o_4 _09581_ (.A1(\tms1x00.ins_pla_ors[12][23] ),
    .A2(net427),
    .B1(net417),
    .B2(\tms1x00.ins_pla_ors[12][22] ),
    .C1(_04639_),
    .X(_04643_));
 sky130_fd_sc_hd__a221o_2 _09582_ (.A1(\tms1x00.ins_pla_ors[12][26] ),
    .A2(net454),
    .B1(net422),
    .B2(\tms1x00.ins_pla_ors[12][27] ),
    .C1(_04640_),
    .X(_04644_));
 sky130_fd_sc_hd__a22o_1 _09583_ (.A1(\tms1x00.ins_pla_ors[12][20] ),
    .A2(net452),
    .B1(net418),
    .B2(\tms1x00.ins_pla_ors[12][21] ),
    .X(_04645_));
 sky130_fd_sc_hd__a221o_2 _09584_ (.A1(\tms1x00.ins_pla_ors[12][15] ),
    .A2(net410),
    .B1(net408),
    .B2(\tms1x00.ins_pla_ors[12][14] ),
    .C1(_04645_),
    .X(_04646_));
 sky130_fd_sc_hd__a221o_2 _09585_ (.A1(\tms1x00.ins_pla_ors[12][0] ),
    .A2(net440),
    .B1(net434),
    .B2(\tms1x00.ins_pla_ors[12][1] ),
    .C1(_04642_),
    .X(_04647_));
 sky130_fd_sc_hd__nor4_4 _09586_ (.A(_04643_),
    .B(_04644_),
    .C(_04646_),
    .D(_04647_),
    .Y(_04648_));
 sky130_fd_sc_hd__a22o_1 _09587_ (.A1(\tms1x00.ins_pla_ors[12][16] ),
    .A2(net444),
    .B1(net412),
    .B2(\tms1x00.ins_pla_ors[12][17] ),
    .X(_04649_));
 sky130_fd_sc_hd__a221o_1 _09588_ (.A1(\tms1x00.ins_pla_ors[12][18] ),
    .A2(net430),
    .B1(net406),
    .B2(\tms1x00.ins_pla_ors[12][19] ),
    .C1(_04649_),
    .X(_04650_));
 sky130_fd_sc_hd__a22o_1 _09589_ (.A1(\tms1x00.ins_pla_ors[12][24] ),
    .A2(net456),
    .B1(net404),
    .B2(\tms1x00.ins_pla_ors[12][25] ),
    .X(_04651_));
 sky130_fd_sc_hd__a221o_1 _09590_ (.A1(\tms1x00.ins_pla_ors[12][13] ),
    .A2(net436),
    .B1(net424),
    .B2(\tms1x00.ins_pla_ors[12][12] ),
    .C1(_04651_),
    .X(_04652_));
 sky130_fd_sc_hd__a22o_1 _09591_ (.A1(\tms1x00.ins_pla_ors[12][9] ),
    .A2(net414),
    .B1(net398),
    .B2(\tms1x00.ins_pla_ors[12][8] ),
    .X(_04653_));
 sky130_fd_sc_hd__a221o_1 _09592_ (.A1(\tms1x00.ins_pla_ors[12][11] ),
    .A2(net448),
    .B1(net420),
    .B2(\tms1x00.ins_pla_ors[12][10] ),
    .C1(_04641_),
    .X(_04654_));
 sky130_fd_sc_hd__nor4_2 _09593_ (.A(_04650_),
    .B(_04652_),
    .C(_04653_),
    .D(_04654_),
    .Y(_04655_));
 sky130_fd_sc_hd__and4_1 _09594_ (.A(\tms1x00.N[0] ),
    .B(_04638_),
    .C(_04648_),
    .D(_04655_),
    .X(_04656_));
 sky130_fd_sc_hd__a31o_1 _09595_ (.A1(_04638_),
    .A2(_04648_),
    .A3(_04655_),
    .B1(\tms1x00.N[0] ),
    .X(_04657_));
 sky130_fd_sc_hd__nand2b_1 _09596_ (.A_N(_04656_),
    .B(_04657_),
    .Y(_04658_));
 sky130_fd_sc_hd__a21o_2 _09597_ (.A1(\tms1x00.P[0] ),
    .A2(_04657_),
    .B1(_04656_),
    .X(_04659_));
 sky130_fd_sc_hd__a21oi_4 _09598_ (.A1(_04626_),
    .A2(_04659_),
    .B1(_04624_),
    .Y(_04660_));
 sky130_fd_sc_hd__or3b_2 _09599_ (.A(_04620_),
    .B(_04660_),
    .C_N(_04623_),
    .X(_04661_));
 sky130_fd_sc_hd__nand2_1 _09600_ (.A(_04619_),
    .B(_04621_),
    .Y(_04662_));
 sky130_fd_sc_hd__a22o_1 _09601_ (.A1(\tms1x00.ins_pla_ors[11][0] ),
    .A2(net440),
    .B1(net424),
    .B2(\tms1x00.ins_pla_ors[11][12] ),
    .X(_04663_));
 sky130_fd_sc_hd__a22o_2 _09602_ (.A1(\tms1x00.ins_pla_ors[11][13] ),
    .A2(net436),
    .B1(net408),
    .B2(\tms1x00.ins_pla_ors[11][14] ),
    .X(_04664_));
 sky130_fd_sc_hd__a22o_1 _09603_ (.A1(\tms1x00.ins_pla_ors[11][3] ),
    .A2(net432),
    .B1(net422),
    .B2(\tms1x00.ins_pla_ors[11][27] ),
    .X(_04665_));
 sky130_fd_sc_hd__a22o_1 _09604_ (.A1(\tms1x00.ins_pla_ors[11][4] ),
    .A2(net442),
    .B1(net416),
    .B2(\tms1x00.ins_pla_ors[11][22] ),
    .X(_04666_));
 sky130_fd_sc_hd__a22o_1 _09605_ (.A1(\tms1x00.ins_pla_ors[11][18] ),
    .A2(net430),
    .B1(net412),
    .B2(\tms1x00.ins_pla_ors[11][17] ),
    .X(_04667_));
 sky130_fd_sc_hd__a22o_1 _09606_ (.A1(\tms1x00.ins_pla_ors[11][11] ),
    .A2(net448),
    .B1(net434),
    .B2(\tms1x00.ins_pla_ors[11][1] ),
    .X(_04668_));
 sky130_fd_sc_hd__a221o_1 _09607_ (.A1(\tms1x00.ins_pla_ors[11][29] ),
    .A2(net429),
    .B1(net402),
    .B2(\tms1x00.ins_pla_ors[11][5] ),
    .C1(_04668_),
    .X(_04669_));
 sky130_fd_sc_hd__a22o_1 _09608_ (.A1(\tms1x00.ins_pla_ors[11][24] ),
    .A2(net456),
    .B1(net414),
    .B2(\tms1x00.ins_pla_ors[11][9] ),
    .X(_04670_));
 sky130_fd_sc_hd__a221o_1 _09609_ (.A1(\tms1x00.ins_pla_ors[11][7] ),
    .A2(net450),
    .B1(net398),
    .B2(\tms1x00.ins_pla_ors[11][8] ),
    .C1(_04670_),
    .X(_04671_));
 sky130_fd_sc_hd__a22o_1 _09610_ (.A1(\tms1x00.ins_pla_ors[11][26] ),
    .A2(net454),
    .B1(net452),
    .B2(\tms1x00.ins_pla_ors[11][20] ),
    .X(_04672_));
 sky130_fd_sc_hd__a221o_1 _09611_ (.A1(\tms1x00.ins_pla_ors[11][28] ),
    .A2(net447),
    .B1(net418),
    .B2(\tms1x00.ins_pla_ors[11][21] ),
    .C1(_04666_),
    .X(_04673_));
 sky130_fd_sc_hd__a221o_1 _09612_ (.A1(\tms1x00.ins_pla_ors[11][16] ),
    .A2(net444),
    .B1(net400),
    .B2(\tms1x00.ins_pla_ors[11][6] ),
    .C1(_04667_),
    .X(_04674_));
 sky130_fd_sc_hd__a221o_1 _09613_ (.A1(\tms1x00.ins_pla_ors[11][23] ),
    .A2(net426),
    .B1(net404),
    .B2(\tms1x00.ins_pla_ors[11][25] ),
    .C1(_04672_),
    .X(_04675_));
 sky130_fd_sc_hd__a221o_2 _09614_ (.A1(\tms1x00.ins_pla_ors[11][2] ),
    .A2(net438),
    .B1(net420),
    .B2(\tms1x00.ins_pla_ors[11][10] ),
    .C1(_04663_),
    .X(_04676_));
 sky130_fd_sc_hd__or4_2 _09615_ (.A(_04673_),
    .B(_04674_),
    .C(_04675_),
    .D(_04676_),
    .X(_04677_));
 sky130_fd_sc_hd__a221o_1 _09616_ (.A1(\tms1x00.ins_pla_ors[11][15] ),
    .A2(net410),
    .B1(net406),
    .B2(\tms1x00.ins_pla_ors[11][19] ),
    .C1(_04665_),
    .X(_04678_));
 sky130_fd_sc_hd__or4_2 _09617_ (.A(_04664_),
    .B(_04669_),
    .C(_04671_),
    .D(_04678_),
    .X(_04679_));
 sky130_fd_sc_hd__o211a_1 _09618_ (.A1(_04677_),
    .A2(_04679_),
    .B1(_04618_),
    .C1(_04662_),
    .X(_04680_));
 sky130_fd_sc_hd__a22o_1 _09619_ (.A1(\tms1x00.ins_pla_ors[10][29] ),
    .A2(net429),
    .B1(net402),
    .B2(\tms1x00.ins_pla_ors[10][5] ),
    .X(_04681_));
 sky130_fd_sc_hd__a22o_1 _09620_ (.A1(\tms1x00.ins_pla_ors[10][3] ),
    .A2(net432),
    .B1(net422),
    .B2(\tms1x00.ins_pla_ors[10][27] ),
    .X(_04682_));
 sky130_fd_sc_hd__a22o_1 _09621_ (.A1(\tms1x00.ins_pla_ors[10][18] ),
    .A2(net430),
    .B1(net412),
    .B2(\tms1x00.ins_pla_ors[10][17] ),
    .X(_04683_));
 sky130_fd_sc_hd__a22o_1 _09622_ (.A1(\tms1x00.ins_pla_ors[10][4] ),
    .A2(net442),
    .B1(net416),
    .B2(\tms1x00.ins_pla_ors[10][22] ),
    .X(_04684_));
 sky130_fd_sc_hd__a22o_1 _09623_ (.A1(\tms1x00.ins_pla_ors[10][11] ),
    .A2(net448),
    .B1(net434),
    .B2(\tms1x00.ins_pla_ors[10][1] ),
    .X(_04685_));
 sky130_fd_sc_hd__a22o_1 _09624_ (.A1(\tms1x00.ins_pla_ors[10][24] ),
    .A2(net456),
    .B1(net414),
    .B2(\tms1x00.ins_pla_ors[10][9] ),
    .X(_04686_));
 sky130_fd_sc_hd__a22o_1 _09625_ (.A1(\tms1x00.ins_pla_ors[10][7] ),
    .A2(net450),
    .B1(net398),
    .B2(\tms1x00.ins_pla_ors[10][8] ),
    .X(_04687_));
 sky130_fd_sc_hd__or4_1 _09626_ (.A(_04681_),
    .B(_04685_),
    .C(_04686_),
    .D(_04687_),
    .X(_04688_));
 sky130_fd_sc_hd__a22o_1 _09627_ (.A1(\tms1x00.ins_pla_ors[10][26] ),
    .A2(net454),
    .B1(net452),
    .B2(\tms1x00.ins_pla_ors[10][20] ),
    .X(_04689_));
 sky130_fd_sc_hd__a22o_1 _09628_ (.A1(\tms1x00.ins_pla_ors[10][2] ),
    .A2(net438),
    .B1(net420),
    .B2(\tms1x00.ins_pla_ors[10][10] ),
    .X(_04690_));
 sky130_fd_sc_hd__a221o_1 _09629_ (.A1(\tms1x00.ins_pla_ors[10][28] ),
    .A2(net447),
    .B1(net418),
    .B2(\tms1x00.ins_pla_ors[10][21] ),
    .C1(_04684_),
    .X(_04691_));
 sky130_fd_sc_hd__a221o_1 _09630_ (.A1(\tms1x00.ins_pla_ors[10][16] ),
    .A2(net444),
    .B1(net400),
    .B2(\tms1x00.ins_pla_ors[10][6] ),
    .C1(_04683_),
    .X(_04692_));
 sky130_fd_sc_hd__a221o_1 _09631_ (.A1(\tms1x00.ins_pla_ors[10][23] ),
    .A2(net426),
    .B1(net404),
    .B2(\tms1x00.ins_pla_ors[10][25] ),
    .C1(_04689_),
    .X(_04693_));
 sky130_fd_sc_hd__a221o_1 _09632_ (.A1(\tms1x00.ins_pla_ors[10][0] ),
    .A2(net440),
    .B1(net424),
    .B2(\tms1x00.ins_pla_ors[10][12] ),
    .C1(_04690_),
    .X(_04694_));
 sky130_fd_sc_hd__or4_1 _09633_ (.A(_04691_),
    .B(_04692_),
    .C(_04693_),
    .D(_04694_),
    .X(_04695_));
 sky130_fd_sc_hd__a221o_1 _09634_ (.A1(\tms1x00.ins_pla_ors[10][15] ),
    .A2(net410),
    .B1(net406),
    .B2(\tms1x00.ins_pla_ors[10][19] ),
    .C1(_04682_),
    .X(_04696_));
 sky130_fd_sc_hd__a221o_2 _09635_ (.A1(\tms1x00.ins_pla_ors[10][13] ),
    .A2(net436),
    .B1(net408),
    .B2(\tms1x00.ins_pla_ors[10][14] ),
    .C1(_04696_),
    .X(_04697_));
 sky130_fd_sc_hd__or3_2 _09636_ (.A(_04688_),
    .B(_04695_),
    .C(_04697_),
    .X(_04698_));
 sky130_fd_sc_hd__and2_1 _09637_ (.A(\tms1x00.N[0] ),
    .B(\tms1x00.P[0] ),
    .X(_04699_));
 sky130_fd_sc_hd__nor2_1 _09638_ (.A(\tms1x00.N[0] ),
    .B(\tms1x00.P[0] ),
    .Y(_04700_));
 sky130_fd_sc_hd__o221a_1 _09639_ (.A1(_04621_),
    .A2(_04622_),
    .B1(_04699_),
    .B2(_04700_),
    .C1(_04620_),
    .X(_04701_));
 sky130_fd_sc_hd__and3b_1 _09640_ (.A_N(_04626_),
    .B(_04698_),
    .C(_04701_),
    .X(_04702_));
 sky130_fd_sc_hd__a21oi_2 _09641_ (.A1(_04661_),
    .A2(_04680_),
    .B1(_04702_),
    .Y(_04703_));
 sky130_fd_sc_hd__a22o_1 _09642_ (.A1(\tms1x00.ins_pla_ors[15][28] ),
    .A2(net447),
    .B1(net426),
    .B2(\tms1x00.ins_pla_ors[15][23] ),
    .X(_04704_));
 sky130_fd_sc_hd__a221o_2 _09643_ (.A1(\tms1x00.ins_pla_ors[15][16] ),
    .A2(net444),
    .B1(net416),
    .B2(\tms1x00.ins_pla_ors[15][22] ),
    .C1(_04704_),
    .X(_04705_));
 sky130_fd_sc_hd__a22o_1 _09644_ (.A1(\tms1x00.ins_pla_ors[15][21] ),
    .A2(net418),
    .B1(net412),
    .B2(\tms1x00.ins_pla_ors[15][17] ),
    .X(_04706_));
 sky130_fd_sc_hd__a221o_1 _09645_ (.A1(\tms1x00.ins_pla_ors[15][0] ),
    .A2(net440),
    .B1(net436),
    .B2(\tms1x00.ins_pla_ors[15][13] ),
    .C1(_04706_),
    .X(_04707_));
 sky130_fd_sc_hd__a22o_1 _09646_ (.A1(\tms1x00.ins_pla_ors[15][26] ),
    .A2(net454),
    .B1(net420),
    .B2(\tms1x00.ins_pla_ors[15][10] ),
    .X(_04708_));
 sky130_fd_sc_hd__a21o_1 _09647_ (.A1(\tms1x00.ins_pla_ors[15][15] ),
    .A2(net410),
    .B1(_04708_),
    .X(_04709_));
 sky130_fd_sc_hd__a22o_1 _09648_ (.A1(\tms1x00.ins_pla_ors[15][14] ),
    .A2(net408),
    .B1(net406),
    .B2(\tms1x00.ins_pla_ors[15][19] ),
    .X(_04710_));
 sky130_fd_sc_hd__a221o_1 _09649_ (.A1(\tms1x00.ins_pla_ors[15][25] ),
    .A2(net404),
    .B1(net400),
    .B2(\tms1x00.ins_pla_ors[15][6] ),
    .C1(_04710_),
    .X(_04711_));
 sky130_fd_sc_hd__or4_2 _09650_ (.A(_04705_),
    .B(_04707_),
    .C(_04709_),
    .D(_04711_),
    .X(_04712_));
 sky130_fd_sc_hd__a22o_1 _09651_ (.A1(\tms1x00.ins_pla_ors[15][18] ),
    .A2(net430),
    .B1(net424),
    .B2(\tms1x00.ins_pla_ors[15][12] ),
    .X(_04713_));
 sky130_fd_sc_hd__a221o_1 _09652_ (.A1(\tms1x00.ins_pla_ors[15][24] ),
    .A2(net456),
    .B1(net398),
    .B2(\tms1x00.ins_pla_ors[15][8] ),
    .C1(_04713_),
    .X(_04714_));
 sky130_fd_sc_hd__a21bo_1 _09653_ (.A1(\tms1x00.ins_pla_ors[15][1] ),
    .A2(net434),
    .B1_N(_04608_),
    .X(_04715_));
 sky130_fd_sc_hd__a221o_1 _09654_ (.A1(\tms1x00.ins_pla_ors[15][7] ),
    .A2(net450),
    .B1(net432),
    .B2(\tms1x00.ins_pla_ors[15][3] ),
    .C1(_04715_),
    .X(_04716_));
 sky130_fd_sc_hd__a22o_1 _09655_ (.A1(\tms1x00.ins_pla_ors[15][20] ),
    .A2(net452),
    .B1(net422),
    .B2(\tms1x00.ins_pla_ors[15][27] ),
    .X(_04717_));
 sky130_fd_sc_hd__a221o_1 _09656_ (.A1(\tms1x00.ins_pla_ors[15][29] ),
    .A2(net429),
    .B1(net414),
    .B2(\tms1x00.ins_pla_ors[15][9] ),
    .C1(_04717_),
    .X(_04718_));
 sky130_fd_sc_hd__a22o_1 _09657_ (.A1(\tms1x00.ins_pla_ors[15][11] ),
    .A2(net448),
    .B1(net442),
    .B2(\tms1x00.ins_pla_ors[15][4] ),
    .X(_04719_));
 sky130_fd_sc_hd__a221o_1 _09658_ (.A1(\tms1x00.ins_pla_ors[15][2] ),
    .A2(net438),
    .B1(net402),
    .B2(\tms1x00.ins_pla_ors[15][5] ),
    .C1(_04719_),
    .X(_04720_));
 sky130_fd_sc_hd__or4_1 _09659_ (.A(_04714_),
    .B(_04716_),
    .C(_04718_),
    .D(_04720_),
    .X(_04721_));
 sky130_fd_sc_hd__o21bai_2 _09660_ (.A1(_04712_),
    .A2(_04721_),
    .B1_N(net340),
    .Y(_04722_));
 sky130_fd_sc_hd__and2b_1 _09661_ (.A_N(_04722_),
    .B(_04608_),
    .X(_04723_));
 sky130_fd_sc_hd__a221o_1 _09662_ (.A1(\tms1x00.SL ),
    .A2(_04722_),
    .B1(_04723_),
    .B2(_04703_),
    .C1(net592),
    .X(_01431_));
 sky130_fd_sc_hd__a211o_1 _09663_ (.A1(_04661_),
    .A2(_04680_),
    .B1(_04702_),
    .C1(net340),
    .X(_04724_));
 sky130_fd_sc_hd__a21oi_1 _09664_ (.A1(\tms1x00.status ),
    .A2(net340),
    .B1(net592),
    .Y(_04725_));
 sky130_fd_sc_hd__nand2_1 _09665_ (.A(_04724_),
    .B(_04725_),
    .Y(_01432_));
 sky130_fd_sc_hd__a211o_1 _09666_ (.A1(\tms1x00.CA ),
    .A2(net705),
    .B1(_04532_),
    .C1(\tms1x00.CL ),
    .X(_04726_));
 sky130_fd_sc_hd__o211a_1 _09667_ (.A1(\tms1x00.CS ),
    .A2(_04533_),
    .B1(_04726_),
    .C1(net633),
    .X(_01433_));
 sky130_fd_sc_hd__or4_4 _09668_ (.A(_01638_),
    .B(_03378_),
    .C(_03400_),
    .D(_04303_),
    .X(_04727_));
 sky130_fd_sc_hd__nor2_2 _09669_ (.A(net340),
    .B(_04727_),
    .Y(_04728_));
 sky130_fd_sc_hd__o21a_1 _09670_ (.A1(\tms1x00.CB ),
    .A2(_04728_),
    .B1(net637),
    .X(_04729_));
 sky130_fd_sc_hd__a21boi_1 _09671_ (.A1(\tms1x00.CB ),
    .A2(_04728_),
    .B1_N(_04729_),
    .Y(_01434_));
 sky130_fd_sc_hd__nor2_2 _09672_ (.A(\tms1x00.CL ),
    .B(_04530_),
    .Y(_04730_));
 sky130_fd_sc_hd__nand2_8 _09673_ (.A(\tms1x00.CL ),
    .B(_04616_),
    .Y(_04731_));
 sky130_fd_sc_hd__inv_2 _09674_ (.A(_04731_),
    .Y(_04732_));
 sky130_fd_sc_hd__a22o_1 _09675_ (.A1(\tms1x00.CB ),
    .A2(_04730_),
    .B1(_04732_),
    .B2(\tms1x00.CS ),
    .X(_04733_));
 sky130_fd_sc_hd__o21ai_1 _09676_ (.A1(_04730_),
    .A2(_04732_),
    .B1(_04617_),
    .Y(_04734_));
 sky130_fd_sc_hd__a32o_1 _09677_ (.A1(net705),
    .A2(_04617_),
    .A3(_04733_),
    .B1(_04734_),
    .B2(\tms1x00.CA ),
    .X(_04735_));
 sky130_fd_sc_hd__and2_1 _09678_ (.A(net633),
    .B(_04735_),
    .X(_01435_));
 sky130_fd_sc_hd__nand2_1 _09679_ (.A(\tms1x00.cycle[0] ),
    .B(_01625_),
    .Y(_04736_));
 sky130_fd_sc_hd__or4b_1 _09680_ (.A(\tms1x00.cycle[2] ),
    .B(net668),
    .C(net672),
    .D_N(\tms1x00.cycle[1] ),
    .X(_04737_));
 sky130_fd_sc_hd__or4_4 _09681_ (.A(_01626_),
    .B(net458),
    .C(_04736_),
    .D(_04737_),
    .X(_04738_));
 sky130_fd_sc_hd__nand2_2 _09682_ (.A(_04532_),
    .B(_04738_),
    .Y(_04739_));
 sky130_fd_sc_hd__or2_1 _09683_ (.A(\tms1x00.PA[0] ),
    .B(_04532_),
    .X(_04740_));
 sky130_fd_sc_hd__o221a_1 _09684_ (.A1(net686),
    .A2(_04738_),
    .B1(_04739_),
    .B2(\tms1x00.PB[0] ),
    .C1(_04740_),
    .X(_04741_));
 sky130_fd_sc_hd__or2_1 _09685_ (.A(net591),
    .B(_04741_),
    .X(_01436_));
 sky130_fd_sc_hd__or2_1 _09686_ (.A(\tms1x00.PA[1] ),
    .B(_04532_),
    .X(_04742_));
 sky130_fd_sc_hd__o221a_1 _09687_ (.A1(net691),
    .A2(_04738_),
    .B1(_04739_),
    .B2(\tms1x00.PB[1] ),
    .C1(_04742_),
    .X(_04743_));
 sky130_fd_sc_hd__or2_1 _09688_ (.A(net591),
    .B(_04743_),
    .X(_01437_));
 sky130_fd_sc_hd__or2_1 _09689_ (.A(\tms1x00.PA[2] ),
    .B(_04532_),
    .X(_04744_));
 sky130_fd_sc_hd__o221a_1 _09690_ (.A1(net696),
    .A2(_04738_),
    .B1(_04739_),
    .B2(\tms1x00.PB[2] ),
    .C1(_04744_),
    .X(_04745_));
 sky130_fd_sc_hd__or2_1 _09691_ (.A(net591),
    .B(_04745_),
    .X(_01438_));
 sky130_fd_sc_hd__or2_1 _09692_ (.A(\tms1x00.PA[3] ),
    .B(_04532_),
    .X(_04746_));
 sky130_fd_sc_hd__o221a_1 _09693_ (.A1(net700),
    .A2(_04738_),
    .B1(_04739_),
    .B2(\tms1x00.PB[3] ),
    .C1(_04746_),
    .X(_04747_));
 sky130_fd_sc_hd__or2_1 _09694_ (.A(net591),
    .B(_04747_),
    .X(_01439_));
 sky130_fd_sc_hd__o21ai_4 _09695_ (.A1(_04616_),
    .A2(_04730_),
    .B1(_04617_),
    .Y(_04748_));
 sky130_fd_sc_hd__mux2_1 _09696_ (.A0(\tms1x00.PB[0] ),
    .A1(\tms1x00.PA[0] ),
    .S(_04748_),
    .X(_04749_));
 sky130_fd_sc_hd__or2_1 _09697_ (.A(net591),
    .B(_04749_),
    .X(_01440_));
 sky130_fd_sc_hd__mux2_1 _09698_ (.A0(\tms1x00.PB[1] ),
    .A1(\tms1x00.PA[1] ),
    .S(_04748_),
    .X(_04750_));
 sky130_fd_sc_hd__or2_1 _09699_ (.A(net591),
    .B(_04750_),
    .X(_01441_));
 sky130_fd_sc_hd__mux2_1 _09700_ (.A0(\tms1x00.PB[2] ),
    .A1(\tms1x00.PA[2] ),
    .S(_04748_),
    .X(_04751_));
 sky130_fd_sc_hd__or2_1 _09701_ (.A(net591),
    .B(_04751_),
    .X(_01442_));
 sky130_fd_sc_hd__mux2_1 _09702_ (.A0(\tms1x00.PB[3] ),
    .A1(\tms1x00.PA[3] ),
    .S(_04748_),
    .X(_04752_));
 sky130_fd_sc_hd__or2_1 _09703_ (.A(net591),
    .B(_04752_),
    .X(_01443_));
 sky130_fd_sc_hd__nor2_8 _09704_ (.A(\tms1x00.cycle[0] ),
    .B(net339),
    .Y(_04753_));
 sky130_fd_sc_hd__a22o_1 _09705_ (.A1(\tms1x00.ins_pla_ors[3][1] ),
    .A2(net435),
    .B1(net433),
    .B2(\tms1x00.ins_pla_ors[3][3] ),
    .X(_04754_));
 sky130_fd_sc_hd__a221o_1 _09706_ (.A1(\tms1x00.ins_pla_ors[3][28] ),
    .A2(net446),
    .B1(net399),
    .B2(\tms1x00.ins_pla_ors[3][8] ),
    .C1(_04754_),
    .X(_04755_));
 sky130_fd_sc_hd__a22o_1 _09707_ (.A1(\tms1x00.ins_pla_ors[3][16] ),
    .A2(net445),
    .B1(net421),
    .B2(\tms1x00.ins_pla_ors[3][10] ),
    .X(_04756_));
 sky130_fd_sc_hd__a221o_1 _09708_ (.A1(\tms1x00.ins_pla_ors[3][0] ),
    .A2(net441),
    .B1(net437),
    .B2(\tms1x00.ins_pla_ors[3][13] ),
    .C1(_04756_),
    .X(_04757_));
 sky130_fd_sc_hd__a22o_2 _09709_ (.A1(\tms1x00.ins_pla_ors[3][7] ),
    .A2(net451),
    .B1(net449),
    .B2(\tms1x00.ins_pla_ors[3][11] ),
    .X(_04758_));
 sky130_fd_sc_hd__a221o_1 _09710_ (.A1(\tms1x00.ins_pla_ors[3][20] ),
    .A2(net453),
    .B1(net413),
    .B2(\tms1x00.ins_pla_ors[3][17] ),
    .C1(_04758_),
    .X(_04759_));
 sky130_fd_sc_hd__a22o_1 _09711_ (.A1(\tms1x00.ins_pla_ors[3][26] ),
    .A2(net455),
    .B1(net419),
    .B2(\tms1x00.ins_pla_ors[3][21] ),
    .X(_04760_));
 sky130_fd_sc_hd__a221o_1 _09712_ (.A1(\tms1x00.ins_pla_ors[3][9] ),
    .A2(net415),
    .B1(net403),
    .B2(\tms1x00.ins_pla_ors[3][5] ),
    .C1(_04760_),
    .X(_04761_));
 sky130_fd_sc_hd__or4_1 _09713_ (.A(_04755_),
    .B(_04757_),
    .C(_04759_),
    .D(_04761_),
    .X(_04762_));
 sky130_fd_sc_hd__a22o_1 _09714_ (.A1(\tms1x00.ins_pla_ors[3][22] ),
    .A2(net417),
    .B1(net411),
    .B2(\tms1x00.ins_pla_ors[3][15] ),
    .X(_04763_));
 sky130_fd_sc_hd__a221o_1 _09715_ (.A1(\tms1x00.ins_pla_ors[3][18] ),
    .A2(net431),
    .B1(net409),
    .B2(\tms1x00.ins_pla_ors[3][14] ),
    .C1(_04763_),
    .X(_04764_));
 sky130_fd_sc_hd__a221o_1 _09716_ (.A1(\tms1x00.ins_pla_ors[3][27] ),
    .A2(net423),
    .B1(net405),
    .B2(\tms1x00.ins_pla_ors[3][25] ),
    .C1(_04764_),
    .X(_04765_));
 sky130_fd_sc_hd__a22o_1 _09717_ (.A1(\tms1x00.ins_pla_ors[3][4] ),
    .A2(net443),
    .B1(net439),
    .B2(\tms1x00.ins_pla_ors[3][2] ),
    .X(_04766_));
 sky130_fd_sc_hd__a221o_1 _09718_ (.A1(\tms1x00.ins_pla_ors[3][23] ),
    .A2(net427),
    .B1(net425),
    .B2(\tms1x00.ins_pla_ors[3][12] ),
    .C1(_04766_),
    .X(_04767_));
 sky130_fd_sc_hd__a22o_1 _09719_ (.A1(\tms1x00.ins_pla_ors[3][24] ),
    .A2(net457),
    .B1(net401),
    .B2(\tms1x00.ins_pla_ors[3][6] ),
    .X(_04768_));
 sky130_fd_sc_hd__a221o_1 _09720_ (.A1(\tms1x00.ins_pla_ors[3][29] ),
    .A2(net428),
    .B1(net407),
    .B2(\tms1x00.ins_pla_ors[3][19] ),
    .C1(_04768_),
    .X(_04769_));
 sky130_fd_sc_hd__or4_4 _09721_ (.A(_04762_),
    .B(_04765_),
    .C(_04767_),
    .D(_04769_),
    .X(_04770_));
 sky130_fd_sc_hd__nor2_2 _09722_ (.A(_04637_),
    .B(_04770_),
    .Y(_04771_));
 sky130_fd_sc_hd__a22o_1 _09723_ (.A1(\tms1x00.ins_pla_ors[4][18] ),
    .A2(net431),
    .B1(net428),
    .B2(\tms1x00.ins_pla_ors[4][29] ),
    .X(_04772_));
 sky130_fd_sc_hd__a221o_1 _09724_ (.A1(\tms1x00.ins_pla_ors[4][20] ),
    .A2(net453),
    .B1(net417),
    .B2(\tms1x00.ins_pla_ors[4][22] ),
    .C1(_04772_),
    .X(_04773_));
 sky130_fd_sc_hd__a22o_1 _09725_ (.A1(\tms1x00.ins_pla_ors[4][4] ),
    .A2(net443),
    .B1(net437),
    .B2(\tms1x00.ins_pla_ors[4][13] ),
    .X(_04774_));
 sky130_fd_sc_hd__a221o_1 _09726_ (.A1(\tms1x00.ins_pla_ors[4][21] ),
    .A2(net419),
    .B1(net403),
    .B2(\tms1x00.ins_pla_ors[4][5] ),
    .C1(_04774_),
    .X(_04775_));
 sky130_fd_sc_hd__a22o_1 _09727_ (.A1(\tms1x00.ins_pla_ors[4][28] ),
    .A2(net446),
    .B1(net445),
    .B2(\tms1x00.ins_pla_ors[4][16] ),
    .X(_04776_));
 sky130_fd_sc_hd__a221o_1 _09728_ (.A1(\tms1x00.ins_pla_ors[4][12] ),
    .A2(net425),
    .B1(net409),
    .B2(\tms1x00.ins_pla_ors[4][14] ),
    .C1(_04776_),
    .X(_04777_));
 sky130_fd_sc_hd__a22o_1 _09729_ (.A1(\tms1x00.ins_pla_ors[4][1] ),
    .A2(net435),
    .B1(net413),
    .B2(\tms1x00.ins_pla_ors[4][17] ),
    .X(_04778_));
 sky130_fd_sc_hd__a221o_1 _09730_ (.A1(\tms1x00.ins_pla_ors[4][24] ),
    .A2(net457),
    .B1(net449),
    .B2(\tms1x00.ins_pla_ors[4][11] ),
    .C1(_04778_),
    .X(_04779_));
 sky130_fd_sc_hd__or4_1 _09731_ (.A(_04773_),
    .B(_04775_),
    .C(_04777_),
    .D(_04779_),
    .X(_04780_));
 sky130_fd_sc_hd__a22o_1 _09732_ (.A1(\tms1x00.ins_pla_ors[4][26] ),
    .A2(net455),
    .B1(net411),
    .B2(\tms1x00.ins_pla_ors[4][15] ),
    .X(_04781_));
 sky130_fd_sc_hd__a221o_1 _09733_ (.A1(\tms1x00.ins_pla_ors[4][27] ),
    .A2(net423),
    .B1(net399),
    .B2(\tms1x00.ins_pla_ors[4][8] ),
    .C1(_04781_),
    .X(_04782_));
 sky130_fd_sc_hd__a221o_1 _09734_ (.A1(\tms1x00.ins_pla_ors[4][3] ),
    .A2(net433),
    .B1(net401),
    .B2(\tms1x00.ins_pla_ors[4][6] ),
    .C1(_04782_),
    .X(_04783_));
 sky130_fd_sc_hd__a22o_1 _09735_ (.A1(\tms1x00.ins_pla_ors[4][7] ),
    .A2(net451),
    .B1(net405),
    .B2(\tms1x00.ins_pla_ors[4][25] ),
    .X(_04784_));
 sky130_fd_sc_hd__a221o_1 _09736_ (.A1(\tms1x00.ins_pla_ors[4][2] ),
    .A2(net439),
    .B1(net427),
    .B2(\tms1x00.ins_pla_ors[4][23] ),
    .C1(_04784_),
    .X(_04785_));
 sky130_fd_sc_hd__a22o_1 _09737_ (.A1(\tms1x00.ins_pla_ors[4][0] ),
    .A2(net441),
    .B1(net407),
    .B2(\tms1x00.ins_pla_ors[4][19] ),
    .X(_04786_));
 sky130_fd_sc_hd__a221o_2 _09738_ (.A1(\tms1x00.ins_pla_ors[4][10] ),
    .A2(net421),
    .B1(net415),
    .B2(\tms1x00.ins_pla_ors[4][9] ),
    .C1(_04786_),
    .X(_04787_));
 sky130_fd_sc_hd__or4_2 _09739_ (.A(_04780_),
    .B(_04783_),
    .C(_04785_),
    .D(_04787_),
    .X(_04788_));
 sky130_fd_sc_hd__nor2_2 _09740_ (.A(_04637_),
    .B(_04788_),
    .Y(_04789_));
 sky130_fd_sc_hd__a22o_1 _09741_ (.A1(\tms1x00.ins_pla_ors[2][13] ),
    .A2(net437),
    .B1(net435),
    .B2(\tms1x00.ins_pla_ors[2][1] ),
    .X(_04790_));
 sky130_fd_sc_hd__a221o_1 _09742_ (.A1(\tms1x00.ins_pla_ors[2][28] ),
    .A2(net446),
    .B1(net441),
    .B2(\tms1x00.ins_pla_ors[2][0] ),
    .C1(_04790_),
    .X(_04791_));
 sky130_fd_sc_hd__a22o_1 _09743_ (.A1(\tms1x00.ins_pla_ors[2][3] ),
    .A2(net433),
    .B1(net403),
    .B2(\tms1x00.ins_pla_ors[2][5] ),
    .X(_04792_));
 sky130_fd_sc_hd__a221o_1 _09744_ (.A1(\tms1x00.ins_pla_ors[2][4] ),
    .A2(net443),
    .B1(net415),
    .B2(\tms1x00.ins_pla_ors[2][9] ),
    .C1(_04792_),
    .X(_04793_));
 sky130_fd_sc_hd__a22o_1 _09745_ (.A1(\tms1x00.ins_pla_ors[2][7] ),
    .A2(net451),
    .B1(net439),
    .B2(\tms1x00.ins_pla_ors[2][2] ),
    .X(_04794_));
 sky130_fd_sc_hd__a221o_1 _09746_ (.A1(\tms1x00.ins_pla_ors[2][20] ),
    .A2(net453),
    .B1(net413),
    .B2(\tms1x00.ins_pla_ors[2][17] ),
    .C1(_04794_),
    .X(_04795_));
 sky130_fd_sc_hd__a22o_1 _09747_ (.A1(\tms1x00.ins_pla_ors[2][26] ),
    .A2(net455),
    .B1(net419),
    .B2(\tms1x00.ins_pla_ors[2][21] ),
    .X(_04796_));
 sky130_fd_sc_hd__a221o_1 _09748_ (.A1(\tms1x00.ins_pla_ors[2][11] ),
    .A2(net449),
    .B1(net427),
    .B2(\tms1x00.ins_pla_ors[2][23] ),
    .C1(_04796_),
    .X(_04797_));
 sky130_fd_sc_hd__or4_1 _09749_ (.A(_04791_),
    .B(_04793_),
    .C(_04795_),
    .D(_04797_),
    .X(_04798_));
 sky130_fd_sc_hd__a22o_1 _09750_ (.A1(\tms1x00.ins_pla_ors[2][22] ),
    .A2(net417),
    .B1(net411),
    .B2(\tms1x00.ins_pla_ors[2][15] ),
    .X(_04799_));
 sky130_fd_sc_hd__a221o_1 _09751_ (.A1(\tms1x00.ins_pla_ors[2][18] ),
    .A2(net431),
    .B1(net407),
    .B2(\tms1x00.ins_pla_ors[2][19] ),
    .C1(_04799_),
    .X(_04800_));
 sky130_fd_sc_hd__a221o_1 _09752_ (.A1(\tms1x00.ins_pla_ors[2][27] ),
    .A2(net423),
    .B1(net405),
    .B2(\tms1x00.ins_pla_ors[2][25] ),
    .C1(_04800_),
    .X(_04801_));
 sky130_fd_sc_hd__a22o_1 _09753_ (.A1(\tms1x00.ins_pla_ors[2][29] ),
    .A2(net428),
    .B1(net425),
    .B2(\tms1x00.ins_pla_ors[2][12] ),
    .X(_04802_));
 sky130_fd_sc_hd__a221o_1 _09754_ (.A1(\tms1x00.ins_pla_ors[2][10] ),
    .A2(net421),
    .B1(net399),
    .B2(\tms1x00.ins_pla_ors[2][8] ),
    .C1(_04802_),
    .X(_04803_));
 sky130_fd_sc_hd__a22o_1 _09755_ (.A1(\tms1x00.ins_pla_ors[2][16] ),
    .A2(net445),
    .B1(net409),
    .B2(\tms1x00.ins_pla_ors[2][14] ),
    .X(_04804_));
 sky130_fd_sc_hd__a221o_1 _09756_ (.A1(\tms1x00.ins_pla_ors[2][24] ),
    .A2(net457),
    .B1(net401),
    .B2(\tms1x00.ins_pla_ors[2][6] ),
    .C1(_04804_),
    .X(_04805_));
 sky130_fd_sc_hd__or4_4 _09757_ (.A(_04798_),
    .B(_04801_),
    .C(_04803_),
    .D(_04805_),
    .X(_04806_));
 sky130_fd_sc_hd__nor2_2 _09758_ (.A(_04637_),
    .B(_04806_),
    .Y(_04807_));
 sky130_fd_sc_hd__a22o_1 _09759_ (.A1(net656),
    .A2(_04771_),
    .B1(_04807_),
    .B2(_03384_),
    .X(_04808_));
 sky130_fd_sc_hd__a21o_1 _09760_ (.A1(net6),
    .A2(_04789_),
    .B1(_04808_),
    .X(_04809_));
 sky130_fd_sc_hd__mux2_1 _09761_ (.A0(\tms1x00.P[0] ),
    .A1(_04809_),
    .S(_04753_),
    .X(_01444_));
 sky130_fd_sc_hd__a22o_1 _09762_ (.A1(net655),
    .A2(_04771_),
    .B1(_04807_),
    .B2(_03390_),
    .X(_04810_));
 sky130_fd_sc_hd__a21o_1 _09763_ (.A1(net7),
    .A2(_04789_),
    .B1(_04810_),
    .X(_04811_));
 sky130_fd_sc_hd__mux2_1 _09764_ (.A0(\tms1x00.P[1] ),
    .A1(_04811_),
    .S(_04753_),
    .X(_01445_));
 sky130_fd_sc_hd__a22o_1 _09765_ (.A1(net653),
    .A2(_04771_),
    .B1(_04807_),
    .B2(_03396_),
    .X(_04812_));
 sky130_fd_sc_hd__a21o_1 _09766_ (.A1(net8),
    .A2(_04789_),
    .B1(_04812_),
    .X(_04813_));
 sky130_fd_sc_hd__mux2_1 _09767_ (.A0(\tms1x00.P[2] ),
    .A1(_04813_),
    .S(_04753_),
    .X(_01446_));
 sky130_fd_sc_hd__a22o_1 _09768_ (.A1(net651),
    .A2(_04771_),
    .B1(_04807_),
    .B2(_03402_),
    .X(_04814_));
 sky130_fd_sc_hd__a21o_1 _09769_ (.A1(net9),
    .A2(_04789_),
    .B1(_04814_),
    .X(_04815_));
 sky130_fd_sc_hd__mux2_1 _09770_ (.A0(\tms1x00.P[3] ),
    .A1(_04815_),
    .S(_04753_),
    .X(_01447_));
 sky130_fd_sc_hd__a211oi_4 _09771_ (.A1(_04530_),
    .A2(_04731_),
    .B1(_01622_),
    .C1(_04522_),
    .Y(_04816_));
 sky130_fd_sc_hd__o22a_1 _09772_ (.A1(net701),
    .A2(_04530_),
    .B1(_04731_),
    .B2(\tms1x00.SR[0] ),
    .X(_04817_));
 sky130_fd_sc_hd__o221a_1 _09773_ (.A1(\tms1x00.PC[0] ),
    .A2(_04816_),
    .B1(_04817_),
    .B2(net593),
    .C1(_04524_),
    .X(_04818_));
 sky130_fd_sc_hd__and4_1 _09774_ (.A(\tms1x00.PC[3] ),
    .B(\tms1x00.PC[2] ),
    .C(\tms1x00.PC[1] ),
    .D(\tms1x00.PC[0] ),
    .X(_04819_));
 sky130_fd_sc_hd__or3_1 _09775_ (.A(\tms1x00.PC[5] ),
    .B(_01615_),
    .C(_04819_),
    .X(_04820_));
 sky130_fd_sc_hd__o21ai_1 _09776_ (.A1(_01615_),
    .A2(_04819_),
    .B1(\tms1x00.PC[5] ),
    .Y(_04821_));
 sky130_fd_sc_hd__a31o_1 _09777_ (.A1(_04523_),
    .A2(_04820_),
    .A3(_04821_),
    .B1(net458),
    .X(_04822_));
 sky130_fd_sc_hd__o221a_1 _09778_ (.A1(\tms1x00.PC[0] ),
    .A2(_03373_),
    .B1(_04818_),
    .B2(_04822_),
    .C1(net631),
    .X(_01448_));
 sky130_fd_sc_hd__o22a_1 _09779_ (.A1(net697),
    .A2(_04530_),
    .B1(_04731_),
    .B2(\tms1x00.SR[1] ),
    .X(_04823_));
 sky130_fd_sc_hd__o221a_1 _09780_ (.A1(\tms1x00.PC[1] ),
    .A2(_04816_),
    .B1(_04823_),
    .B2(net593),
    .C1(_04524_),
    .X(_04824_));
 sky130_fd_sc_hd__a211o_1 _09781_ (.A1(\tms1x00.PC[0] ),
    .A2(_04523_),
    .B1(_04824_),
    .C1(net458),
    .X(_04825_));
 sky130_fd_sc_hd__o211a_1 _09782_ (.A1(\tms1x00.PC[1] ),
    .A2(_03373_),
    .B1(_04825_),
    .C1(net631),
    .X(_01449_));
 sky130_fd_sc_hd__o22a_1 _09783_ (.A1(net692),
    .A2(_04530_),
    .B1(_04731_),
    .B2(\tms1x00.SR[2] ),
    .X(_04826_));
 sky130_fd_sc_hd__o221a_1 _09784_ (.A1(\tms1x00.PC[2] ),
    .A2(_04816_),
    .B1(_04826_),
    .B2(net593),
    .C1(_04524_),
    .X(_04827_));
 sky130_fd_sc_hd__a211o_1 _09785_ (.A1(\tms1x00.PC[1] ),
    .A2(_04523_),
    .B1(_04827_),
    .C1(net458),
    .X(_04828_));
 sky130_fd_sc_hd__o211a_1 _09786_ (.A1(\tms1x00.PC[2] ),
    .A2(_03373_),
    .B1(_04828_),
    .C1(net631),
    .X(_01450_));
 sky130_fd_sc_hd__o22a_1 _09787_ (.A1(net686),
    .A2(_04530_),
    .B1(_04731_),
    .B2(\tms1x00.SR[3] ),
    .X(_04829_));
 sky130_fd_sc_hd__o221a_1 _09788_ (.A1(\tms1x00.PC[3] ),
    .A2(_04816_),
    .B1(_04829_),
    .B2(net593),
    .C1(_04524_),
    .X(_04830_));
 sky130_fd_sc_hd__a211o_1 _09789_ (.A1(\tms1x00.PC[2] ),
    .A2(_04523_),
    .B1(_04830_),
    .C1(net458),
    .X(_04831_));
 sky130_fd_sc_hd__o211a_1 _09790_ (.A1(\tms1x00.PC[3] ),
    .A2(_03373_),
    .B1(_04831_),
    .C1(net631),
    .X(_01451_));
 sky130_fd_sc_hd__o22a_1 _09791_ (.A1(net681),
    .A2(_04530_),
    .B1(_04731_),
    .B2(\tms1x00.SR[4] ),
    .X(_04832_));
 sky130_fd_sc_hd__o221a_1 _09792_ (.A1(\tms1x00.PC[4] ),
    .A2(_04816_),
    .B1(_04832_),
    .B2(net593),
    .C1(_04524_),
    .X(_04833_));
 sky130_fd_sc_hd__a211o_1 _09793_ (.A1(\tms1x00.PC[3] ),
    .A2(_04523_),
    .B1(_04833_),
    .C1(net458),
    .X(_04834_));
 sky130_fd_sc_hd__o211a_1 _09794_ (.A1(\tms1x00.PC[4] ),
    .A2(_03373_),
    .B1(_04834_),
    .C1(net632),
    .X(_01452_));
 sky130_fd_sc_hd__o22a_1 _09795_ (.A1(net679),
    .A2(_04530_),
    .B1(_04731_),
    .B2(\tms1x00.SR[5] ),
    .X(_04835_));
 sky130_fd_sc_hd__o221a_1 _09796_ (.A1(\tms1x00.PC[5] ),
    .A2(_04816_),
    .B1(_04835_),
    .B2(net593),
    .C1(_04524_),
    .X(_04836_));
 sky130_fd_sc_hd__a211o_1 _09797_ (.A1(\tms1x00.PC[4] ),
    .A2(_04523_),
    .B1(_04836_),
    .C1(net458),
    .X(_04837_));
 sky130_fd_sc_hd__o211a_1 _09798_ (.A1(\tms1x00.PC[5] ),
    .A2(_03373_),
    .B1(_04837_),
    .C1(net631),
    .X(_01453_));
 sky130_fd_sc_hd__a22o_1 _09799_ (.A1(\tms1x00.ins_pla_ors[14][11] ),
    .A2(net448),
    .B1(net406),
    .B2(\tms1x00.ins_pla_ors[14][19] ),
    .X(_04838_));
 sky130_fd_sc_hd__a221o_1 _09800_ (.A1(\tms1x00.ins_pla_ors[14][12] ),
    .A2(net424),
    .B1(net408),
    .B2(\tms1x00.ins_pla_ors[14][14] ),
    .C1(_04838_),
    .X(_04839_));
 sky130_fd_sc_hd__a22o_1 _09801_ (.A1(\tms1x00.ins_pla_ors[14][2] ),
    .A2(net438),
    .B1(net402),
    .B2(\tms1x00.ins_pla_ors[14][5] ),
    .X(_04840_));
 sky130_fd_sc_hd__a22o_1 _09802_ (.A1(\tms1x00.ins_pla_ors[14][7] ),
    .A2(net450),
    .B1(net398),
    .B2(\tms1x00.ins_pla_ors[14][8] ),
    .X(_04841_));
 sky130_fd_sc_hd__a22o_1 _09803_ (.A1(\tms1x00.ins_pla_ors[14][10] ),
    .A2(net420),
    .B1(net418),
    .B2(\tms1x00.ins_pla_ors[14][21] ),
    .X(_04842_));
 sky130_fd_sc_hd__a22o_1 _09804_ (.A1(\tms1x00.ins_pla_ors[14][20] ),
    .A2(net452),
    .B1(net412),
    .B2(\tms1x00.ins_pla_ors[14][17] ),
    .X(_04843_));
 sky130_fd_sc_hd__a22o_1 _09805_ (.A1(\tms1x00.ins_pla_ors[14][16] ),
    .A2(net444),
    .B1(net414),
    .B2(\tms1x00.ins_pla_ors[14][9] ),
    .X(_04844_));
 sky130_fd_sc_hd__a22o_1 _09806_ (.A1(\tms1x00.ins_pla_ors[14][3] ),
    .A2(net432),
    .B1(net404),
    .B2(\tms1x00.ins_pla_ors[14][25] ),
    .X(_04845_));
 sky130_fd_sc_hd__a221o_1 _09807_ (.A1(\tms1x00.ins_pla_ors[14][26] ),
    .A2(net454),
    .B1(net416),
    .B2(\tms1x00.ins_pla_ors[14][22] ),
    .C1(_04842_),
    .X(_04846_));
 sky130_fd_sc_hd__a221o_1 _09808_ (.A1(\tms1x00.ins_pla_ors[14][4] ),
    .A2(net442),
    .B1(net436),
    .B2(\tms1x00.ins_pla_ors[14][13] ),
    .C1(_04841_),
    .X(_04847_));
 sky130_fd_sc_hd__a221o_2 _09809_ (.A1(\tms1x00.ins_pla_ors[14][28] ),
    .A2(net447),
    .B1(net428),
    .B2(\tms1x00.ins_pla_ors[14][29] ),
    .C1(_04843_),
    .X(_04848_));
 sky130_fd_sc_hd__a221o_1 _09810_ (.A1(\tms1x00.ins_pla_ors[14][0] ),
    .A2(net440),
    .B1(net434),
    .B2(\tms1x00.ins_pla_ors[14][1] ),
    .C1(_04844_),
    .X(_04849_));
 sky130_fd_sc_hd__or4_1 _09811_ (.A(_04846_),
    .B(_04847_),
    .C(_04848_),
    .D(_04849_),
    .X(_04850_));
 sky130_fd_sc_hd__a22o_1 _09812_ (.A1(\tms1x00.ins_pla_ors[14][24] ),
    .A2(net456),
    .B1(net400),
    .B2(\tms1x00.ins_pla_ors[14][6] ),
    .X(_04851_));
 sky130_fd_sc_hd__a221o_1 _09813_ (.A1(\tms1x00.ins_pla_ors[14][18] ),
    .A2(net430),
    .B1(net410),
    .B2(\tms1x00.ins_pla_ors[14][15] ),
    .C1(_04845_),
    .X(_04852_));
 sky130_fd_sc_hd__a221o_1 _09814_ (.A1(\tms1x00.ins_pla_ors[14][23] ),
    .A2(net426),
    .B1(net422),
    .B2(\tms1x00.ins_pla_ors[14][27] ),
    .C1(_04840_),
    .X(_04853_));
 sky130_fd_sc_hd__or4_1 _09815_ (.A(_04839_),
    .B(_04851_),
    .C(_04852_),
    .D(_04853_),
    .X(_04854_));
 sky130_fd_sc_hd__o21ba_4 _09816_ (.A1(_04850_),
    .A2(_04854_),
    .B1_N(_04306_),
    .X(_04855_));
 sky130_fd_sc_hd__xnor2_2 _09817_ (.A(\tms1x00.P[0] ),
    .B(_04658_),
    .Y(_04856_));
 sky130_fd_sc_hd__mux2_1 _09818_ (.A0(net656),
    .A1(_04856_),
    .S(_04855_),
    .X(_04857_));
 sky130_fd_sc_hd__and2_1 _09819_ (.A(net634),
    .B(_04857_),
    .X(_01454_));
 sky130_fd_sc_hd__xor2_2 _09820_ (.A(_04626_),
    .B(_04659_),
    .X(_04858_));
 sky130_fd_sc_hd__mux2_1 _09821_ (.A0(net655),
    .A1(_04858_),
    .S(_04855_),
    .X(_04859_));
 sky130_fd_sc_hd__and2_1 _09822_ (.A(net634),
    .B(_04859_),
    .X(_01455_));
 sky130_fd_sc_hd__xnor2_2 _09823_ (.A(_04623_),
    .B(_04660_),
    .Y(_04860_));
 sky130_fd_sc_hd__mux2_1 _09824_ (.A0(net653),
    .A1(_04860_),
    .S(_04855_),
    .X(_04861_));
 sky130_fd_sc_hd__and2_1 _09825_ (.A(net634),
    .B(_04861_),
    .X(_01456_));
 sky130_fd_sc_hd__o21ba_1 _09826_ (.A1(_04622_),
    .A2(_04660_),
    .B1_N(_04621_),
    .X(_04862_));
 sky130_fd_sc_hd__xnor2_2 _09827_ (.A(_04620_),
    .B(_04862_),
    .Y(_04863_));
 sky130_fd_sc_hd__o21ai_1 _09828_ (.A1(net651),
    .A2(_04855_),
    .B1(net634),
    .Y(_04864_));
 sky130_fd_sc_hd__a21oi_1 _09829_ (.A1(_04855_),
    .A2(_04863_),
    .B1(_04864_),
    .Y(_01457_));
 sky130_fd_sc_hd__nand2_1 _09830_ (.A(\tms1x00.X[2] ),
    .B(_04309_),
    .Y(_04865_));
 sky130_fd_sc_hd__o211a_1 _09831_ (.A1(net702),
    .A2(_04309_),
    .B1(_04865_),
    .C1(net144),
    .X(_04866_));
 sky130_fd_sc_hd__mux2_1 _09832_ (.A0(_04866_),
    .A1(\tms1x00.X[2] ),
    .S(_04312_),
    .X(_04867_));
 sky130_fd_sc_hd__and2_1 _09833_ (.A(net636),
    .B(_04867_),
    .X(_01458_));
 sky130_fd_sc_hd__a22o_1 _09834_ (.A1(\tms1x00.ins_pla_ors[5][3] ),
    .A2(net433),
    .B1(net421),
    .B2(\tms1x00.ins_pla_ors[5][10] ),
    .X(_04868_));
 sky130_fd_sc_hd__a221o_2 _09835_ (.A1(\tms1x00.ins_pla_ors[5][13] ),
    .A2(net437),
    .B1(net435),
    .B2(\tms1x00.ins_pla_ors[5][1] ),
    .C1(_04868_),
    .X(_04869_));
 sky130_fd_sc_hd__a22o_1 _09836_ (.A1(\tms1x00.ins_pla_ors[5][24] ),
    .A2(net457),
    .B1(net413),
    .B2(\tms1x00.ins_pla_ors[5][17] ),
    .X(_04870_));
 sky130_fd_sc_hd__a221o_1 _09837_ (.A1(\tms1x00.ins_pla_ors[5][11] ),
    .A2(net449),
    .B1(net428),
    .B2(\tms1x00.ins_pla_ors[5][29] ),
    .C1(_04870_),
    .X(_04871_));
 sky130_fd_sc_hd__a22o_1 _09838_ (.A1(\tms1x00.ins_pla_ors[5][16] ),
    .A2(net445),
    .B1(net419),
    .B2(\tms1x00.ins_pla_ors[5][21] ),
    .X(_04872_));
 sky130_fd_sc_hd__a221o_1 _09839_ (.A1(\tms1x00.ins_pla_ors[5][27] ),
    .A2(net423),
    .B1(net415),
    .B2(\tms1x00.ins_pla_ors[5][9] ),
    .C1(_04872_),
    .X(_04873_));
 sky130_fd_sc_hd__a22o_1 _09840_ (.A1(\tms1x00.ins_pla_ors[5][7] ),
    .A2(net451),
    .B1(net441),
    .B2(\tms1x00.ins_pla_ors[5][0] ),
    .X(_04874_));
 sky130_fd_sc_hd__a221o_2 _09841_ (.A1(\tms1x00.ins_pla_ors[5][4] ),
    .A2(net443),
    .B1(net402),
    .B2(\tms1x00.ins_pla_ors[5][5] ),
    .C1(_04874_),
    .X(_04875_));
 sky130_fd_sc_hd__or4_1 _09842_ (.A(_04869_),
    .B(_04871_),
    .C(_04873_),
    .D(_04875_),
    .X(_04876_));
 sky130_fd_sc_hd__a22o_1 _09843_ (.A1(\tms1x00.ins_pla_ors[5][18] ),
    .A2(net431),
    .B1(net401),
    .B2(\tms1x00.ins_pla_ors[5][6] ),
    .X(_04877_));
 sky130_fd_sc_hd__a221o_1 _09844_ (.A1(\tms1x00.ins_pla_ors[5][12] ),
    .A2(net425),
    .B1(net409),
    .B2(\tms1x00.ins_pla_ors[5][14] ),
    .C1(_04877_),
    .X(_04878_));
 sky130_fd_sc_hd__a221o_1 _09845_ (.A1(\tms1x00.ins_pla_ors[5][26] ),
    .A2(net455),
    .B1(net405),
    .B2(\tms1x00.ins_pla_ors[5][25] ),
    .C1(_04878_),
    .X(_04879_));
 sky130_fd_sc_hd__a22o_1 _09846_ (.A1(\tms1x00.ins_pla_ors[5][2] ),
    .A2(net439),
    .B1(net427),
    .B2(\tms1x00.ins_pla_ors[5][23] ),
    .X(_04880_));
 sky130_fd_sc_hd__a221o_1 _09847_ (.A1(\tms1x00.ins_pla_ors[5][20] ),
    .A2(net453),
    .B1(net399),
    .B2(\tms1x00.ins_pla_ors[5][8] ),
    .C1(_04880_),
    .X(_04881_));
 sky130_fd_sc_hd__a22o_1 _09848_ (.A1(\tms1x00.ins_pla_ors[5][22] ),
    .A2(net417),
    .B1(net411),
    .B2(\tms1x00.ins_pla_ors[5][15] ),
    .X(_04882_));
 sky130_fd_sc_hd__a221o_1 _09849_ (.A1(\tms1x00.ins_pla_ors[5][28] ),
    .A2(net446),
    .B1(net407),
    .B2(\tms1x00.ins_pla_ors[5][19] ),
    .C1(_04882_),
    .X(_04883_));
 sky130_fd_sc_hd__or4_4 _09850_ (.A(_04876_),
    .B(_04879_),
    .C(_04881_),
    .D(_04883_),
    .X(_04884_));
 sky130_fd_sc_hd__nor2_2 _09851_ (.A(_04637_),
    .B(_04884_),
    .Y(_04885_));
 sky130_fd_sc_hd__a22o_1 _09852_ (.A1(\tms1x00.ins_pla_ors[6][28] ),
    .A2(net447),
    .B1(net409),
    .B2(\tms1x00.ins_pla_ors[6][14] ),
    .X(_04886_));
 sky130_fd_sc_hd__a22o_1 _09853_ (.A1(\tms1x00.ins_pla_ors[6][23] ),
    .A2(net427),
    .B1(net403),
    .B2(\tms1x00.ins_pla_ors[6][5] ),
    .X(_04887_));
 sky130_fd_sc_hd__a221o_1 _09854_ (.A1(\tms1x00.ins_pla_ors[6][4] ),
    .A2(net443),
    .B1(net437),
    .B2(\tms1x00.ins_pla_ors[6][13] ),
    .C1(_04887_),
    .X(_04888_));
 sky130_fd_sc_hd__a22o_1 _09855_ (.A1(\tms1x00.ins_pla_ors[6][0] ),
    .A2(net441),
    .B1(net415),
    .B2(\tms1x00.ins_pla_ors[6][9] ),
    .X(_04889_));
 sky130_fd_sc_hd__a221o_1 _09856_ (.A1(\tms1x00.ins_pla_ors[6][2] ),
    .A2(net439),
    .B1(net435),
    .B2(\tms1x00.ins_pla_ors[6][1] ),
    .C1(_04889_),
    .X(_04890_));
 sky130_fd_sc_hd__a22o_1 _09857_ (.A1(\tms1x00.ins_pla_ors[6][24] ),
    .A2(net457),
    .B1(net421),
    .B2(\tms1x00.ins_pla_ors[6][10] ),
    .X(_04891_));
 sky130_fd_sc_hd__a221o_1 _09858_ (.A1(\tms1x00.ins_pla_ors[6][7] ),
    .A2(net451),
    .B1(net399),
    .B2(\tms1x00.ins_pla_ors[6][8] ),
    .C1(_04891_),
    .X(_04892_));
 sky130_fd_sc_hd__a22o_1 _09859_ (.A1(\tms1x00.ins_pla_ors[6][21] ),
    .A2(net419),
    .B1(net413),
    .B2(\tms1x00.ins_pla_ors[6][17] ),
    .X(_04893_));
 sky130_fd_sc_hd__a221o_4 _09860_ (.A1(\tms1x00.ins_pla_ors[6][26] ),
    .A2(net455),
    .B1(net453),
    .B2(\tms1x00.ins_pla_ors[6][20] ),
    .C1(_04893_),
    .X(_04894_));
 sky130_fd_sc_hd__or4_1 _09861_ (.A(_04888_),
    .B(_04890_),
    .C(_04892_),
    .D(_04894_),
    .X(_04895_));
 sky130_fd_sc_hd__a22o_1 _09862_ (.A1(\tms1x00.ins_pla_ors[6][16] ),
    .A2(net445),
    .B1(net401),
    .B2(\tms1x00.ins_pla_ors[6][6] ),
    .X(_04896_));
 sky130_fd_sc_hd__a22o_1 _09863_ (.A1(\tms1x00.ins_pla_ors[6][11] ),
    .A2(net449),
    .B1(net430),
    .B2(\tms1x00.ins_pla_ors[6][18] ),
    .X(_04897_));
 sky130_fd_sc_hd__a221o_1 _09864_ (.A1(\tms1x00.ins_pla_ors[6][12] ),
    .A2(net425),
    .B1(net411),
    .B2(\tms1x00.ins_pla_ors[6][15] ),
    .C1(_04897_),
    .X(_04898_));
 sky130_fd_sc_hd__a221o_1 _09865_ (.A1(\tms1x00.ins_pla_ors[6][29] ),
    .A2(net428),
    .B1(net417),
    .B2(\tms1x00.ins_pla_ors[6][22] ),
    .C1(_04886_),
    .X(_04899_));
 sky130_fd_sc_hd__a22o_1 _09866_ (.A1(\tms1x00.ins_pla_ors[6][3] ),
    .A2(net433),
    .B1(net405),
    .B2(\tms1x00.ins_pla_ors[6][25] ),
    .X(_04900_));
 sky130_fd_sc_hd__a221o_1 _09867_ (.A1(\tms1x00.ins_pla_ors[6][27] ),
    .A2(net423),
    .B1(net407),
    .B2(\tms1x00.ins_pla_ors[6][19] ),
    .C1(_04900_),
    .X(_04901_));
 sky130_fd_sc_hd__or4_2 _09868_ (.A(_04896_),
    .B(_04898_),
    .C(_04899_),
    .D(_04901_),
    .X(_04902_));
 sky130_fd_sc_hd__or3_4 _09869_ (.A(_04637_),
    .B(_04895_),
    .C(_04902_),
    .X(_04903_));
 sky130_fd_sc_hd__nor2_1 _09870_ (.A(\tms1x00.A[0] ),
    .B(_04903_),
    .Y(_04904_));
 sky130_fd_sc_hd__a22o_1 _09871_ (.A1(\tms1x00.ins_pla_ors[7][27] ),
    .A2(net423),
    .B1(net407),
    .B2(\tms1x00.ins_pla_ors[7][19] ),
    .X(_04905_));
 sky130_fd_sc_hd__a22o_1 _09872_ (.A1(\tms1x00.ins_pla_ors[7][23] ),
    .A2(net427),
    .B1(net403),
    .B2(\tms1x00.ins_pla_ors[7][5] ),
    .X(_04906_));
 sky130_fd_sc_hd__a221o_1 _09873_ (.A1(\tms1x00.ins_pla_ors[7][4] ),
    .A2(net443),
    .B1(net437),
    .B2(\tms1x00.ins_pla_ors[7][13] ),
    .C1(_04906_),
    .X(_04907_));
 sky130_fd_sc_hd__a22o_1 _09874_ (.A1(\tms1x00.ins_pla_ors[7][0] ),
    .A2(net441),
    .B1(net415),
    .B2(\tms1x00.ins_pla_ors[7][9] ),
    .X(_04908_));
 sky130_fd_sc_hd__a221o_1 _09875_ (.A1(\tms1x00.ins_pla_ors[7][2] ),
    .A2(net439),
    .B1(net435),
    .B2(\tms1x00.ins_pla_ors[7][1] ),
    .C1(_04908_),
    .X(_04909_));
 sky130_fd_sc_hd__a22o_1 _09876_ (.A1(\tms1x00.ins_pla_ors[7][24] ),
    .A2(net457),
    .B1(net421),
    .B2(\tms1x00.ins_pla_ors[7][10] ),
    .X(_04910_));
 sky130_fd_sc_hd__a221o_1 _09877_ (.A1(\tms1x00.ins_pla_ors[7][7] ),
    .A2(net451),
    .B1(net399),
    .B2(\tms1x00.ins_pla_ors[7][8] ),
    .C1(_04910_),
    .X(_04911_));
 sky130_fd_sc_hd__a22o_1 _09878_ (.A1(\tms1x00.ins_pla_ors[7][21] ),
    .A2(net419),
    .B1(net413),
    .B2(\tms1x00.ins_pla_ors[7][17] ),
    .X(_04912_));
 sky130_fd_sc_hd__a221o_4 _09879_ (.A1(\tms1x00.ins_pla_ors[7][26] ),
    .A2(net455),
    .B1(net453),
    .B2(\tms1x00.ins_pla_ors[7][20] ),
    .C1(_04912_),
    .X(_04913_));
 sky130_fd_sc_hd__or4_1 _09880_ (.A(_04907_),
    .B(_04909_),
    .C(_04911_),
    .D(_04913_),
    .X(_04914_));
 sky130_fd_sc_hd__a22o_1 _09881_ (.A1(\tms1x00.ins_pla_ors[7][16] ),
    .A2(net445),
    .B1(net401),
    .B2(\tms1x00.ins_pla_ors[7][6] ),
    .X(_04915_));
 sky130_fd_sc_hd__a22o_1 _09882_ (.A1(\tms1x00.ins_pla_ors[7][29] ),
    .A2(net429),
    .B1(net417),
    .B2(\tms1x00.ins_pla_ors[7][22] ),
    .X(_04916_));
 sky130_fd_sc_hd__a22o_1 _09883_ (.A1(\tms1x00.ins_pla_ors[7][11] ),
    .A2(net449),
    .B1(net431),
    .B2(\tms1x00.ins_pla_ors[7][18] ),
    .X(_04917_));
 sky130_fd_sc_hd__a221o_1 _09884_ (.A1(\tms1x00.ins_pla_ors[7][12] ),
    .A2(net425),
    .B1(net411),
    .B2(\tms1x00.ins_pla_ors[7][15] ),
    .C1(_04917_),
    .X(_04918_));
 sky130_fd_sc_hd__a221o_1 _09885_ (.A1(\tms1x00.ins_pla_ors[7][28] ),
    .A2(net446),
    .B1(net409),
    .B2(\tms1x00.ins_pla_ors[7][14] ),
    .C1(_04916_),
    .X(_04919_));
 sky130_fd_sc_hd__a221o_1 _09886_ (.A1(\tms1x00.ins_pla_ors[7][3] ),
    .A2(net433),
    .B1(net405),
    .B2(\tms1x00.ins_pla_ors[7][25] ),
    .C1(_04905_),
    .X(_04920_));
 sky130_fd_sc_hd__or4_2 _09887_ (.A(_04915_),
    .B(_04918_),
    .C(_04919_),
    .D(_04920_),
    .X(_04921_));
 sky130_fd_sc_hd__or3_2 _09888_ (.A(_04637_),
    .B(_04914_),
    .C(_04921_),
    .X(_04922_));
 sky130_fd_sc_hd__clkinv_2 _09889_ (.A(_04922_),
    .Y(_04923_));
 sky130_fd_sc_hd__a221o_1 _09890_ (.A1(\tms1x00.A[0] ),
    .A2(_04885_),
    .B1(_04923_),
    .B2(net6),
    .C1(_04904_),
    .X(_04924_));
 sky130_fd_sc_hd__a22o_1 _09891_ (.A1(\tms1x00.ins_pla_ors[9][3] ),
    .A2(net432),
    .B1(net418),
    .B2(\tms1x00.ins_pla_ors[9][21] ),
    .X(_04925_));
 sky130_fd_sc_hd__a221o_1 _09892_ (.A1(\tms1x00.ins_pla_ors[9][26] ),
    .A2(net454),
    .B1(net408),
    .B2(\tms1x00.ins_pla_ors[9][14] ),
    .C1(_04925_),
    .X(_04926_));
 sky130_fd_sc_hd__a22o_1 _09893_ (.A1(\tms1x00.ins_pla_ors[9][29] ),
    .A2(net429),
    .B1(net416),
    .B2(\tms1x00.ins_pla_ors[9][22] ),
    .X(_04927_));
 sky130_fd_sc_hd__a221o_1 _09894_ (.A1(\tms1x00.ins_pla_ors[9][20] ),
    .A2(net452),
    .B1(net398),
    .B2(\tms1x00.ins_pla_ors[9][8] ),
    .C1(_04927_),
    .X(_04928_));
 sky130_fd_sc_hd__a22o_1 _09895_ (.A1(\tms1x00.ins_pla_ors[9][27] ),
    .A2(net422),
    .B1(net400),
    .B2(\tms1x00.ins_pla_ors[9][6] ),
    .X(_04929_));
 sky130_fd_sc_hd__a221o_1 _09896_ (.A1(\tms1x00.ins_pla_ors[9][4] ),
    .A2(net442),
    .B1(net406),
    .B2(\tms1x00.ins_pla_ors[9][19] ),
    .C1(_04929_),
    .X(_04930_));
 sky130_fd_sc_hd__a22o_1 _09897_ (.A1(\tms1x00.ins_pla_ors[9][16] ),
    .A2(net444),
    .B1(net412),
    .B2(\tms1x00.ins_pla_ors[9][17] ),
    .X(_04931_));
 sky130_fd_sc_hd__a221o_1 _09898_ (.A1(\tms1x00.ins_pla_ors[9][7] ),
    .A2(net450),
    .B1(net440),
    .B2(\tms1x00.ins_pla_ors[9][0] ),
    .C1(_04931_),
    .X(_04932_));
 sky130_fd_sc_hd__or4_1 _09899_ (.A(_04926_),
    .B(_04928_),
    .C(_04930_),
    .D(_04932_),
    .X(_04933_));
 sky130_fd_sc_hd__a22o_1 _09900_ (.A1(\tms1x00.ins_pla_ors[9][2] ),
    .A2(net438),
    .B1(net430),
    .B2(\tms1x00.ins_pla_ors[9][18] ),
    .X(_04934_));
 sky130_fd_sc_hd__a221o_1 _09901_ (.A1(\tms1x00.ins_pla_ors[9][24] ),
    .A2(net456),
    .B1(net447),
    .B2(\tms1x00.ins_pla_ors[9][28] ),
    .C1(_04934_),
    .X(_04935_));
 sky130_fd_sc_hd__a221o_1 _09902_ (.A1(\tms1x00.ins_pla_ors[9][1] ),
    .A2(net434),
    .B1(net402),
    .B2(\tms1x00.ins_pla_ors[9][5] ),
    .C1(_04935_),
    .X(_04936_));
 sky130_fd_sc_hd__a22o_1 _09903_ (.A1(\tms1x00.ins_pla_ors[9][13] ),
    .A2(net436),
    .B1(net410),
    .B2(\tms1x00.ins_pla_ors[9][15] ),
    .X(_04937_));
 sky130_fd_sc_hd__a221o_1 _09904_ (.A1(\tms1x00.ins_pla_ors[9][10] ),
    .A2(net420),
    .B1(net404),
    .B2(\tms1x00.ins_pla_ors[9][25] ),
    .C1(_04937_),
    .X(_04938_));
 sky130_fd_sc_hd__a22o_1 _09905_ (.A1(\tms1x00.ins_pla_ors[9][12] ),
    .A2(net424),
    .B1(net414),
    .B2(\tms1x00.ins_pla_ors[9][9] ),
    .X(_04939_));
 sky130_fd_sc_hd__a221o_1 _09906_ (.A1(\tms1x00.ins_pla_ors[9][11] ),
    .A2(net448),
    .B1(net426),
    .B2(\tms1x00.ins_pla_ors[9][23] ),
    .C1(_04939_),
    .X(_04940_));
 sky130_fd_sc_hd__or4_4 _09907_ (.A(_04933_),
    .B(_04936_),
    .C(_04938_),
    .D(_04940_),
    .X(_04941_));
 sky130_fd_sc_hd__nor2_2 _09908_ (.A(_04637_),
    .B(_04941_),
    .Y(_04942_));
 sky130_fd_sc_hd__a22o_1 _09909_ (.A1(\tms1x00.ins_pla_ors[8][28] ),
    .A2(net447),
    .B1(net410),
    .B2(\tms1x00.ins_pla_ors[8][15] ),
    .X(_04943_));
 sky130_fd_sc_hd__a221o_1 _09910_ (.A1(\tms1x00.ins_pla_ors[8][24] ),
    .A2(net456),
    .B1(net454),
    .B2(\tms1x00.ins_pla_ors[8][26] ),
    .C1(_04943_),
    .X(_04944_));
 sky130_fd_sc_hd__a22o_1 _09911_ (.A1(\tms1x00.ins_pla_ors[8][7] ),
    .A2(net450),
    .B1(net430),
    .B2(\tms1x00.ins_pla_ors[8][18] ),
    .X(_04945_));
 sky130_fd_sc_hd__a221o_1 _09912_ (.A1(\tms1x00.ins_pla_ors[8][29] ),
    .A2(net429),
    .B1(net424),
    .B2(\tms1x00.ins_pla_ors[8][12] ),
    .C1(_04945_),
    .X(_04946_));
 sky130_fd_sc_hd__a22o_1 _09913_ (.A1(\tms1x00.ins_pla_ors[8][21] ),
    .A2(net418),
    .B1(net414),
    .B2(\tms1x00.ins_pla_ors[8][9] ),
    .X(_04947_));
 sky130_fd_sc_hd__a221o_1 _09914_ (.A1(\tms1x00.ins_pla_ors[8][10] ),
    .A2(net420),
    .B1(net402),
    .B2(\tms1x00.ins_pla_ors[8][5] ),
    .C1(_04947_),
    .X(_04948_));
 sky130_fd_sc_hd__a22o_1 _09915_ (.A1(\tms1x00.ins_pla_ors[8][11] ),
    .A2(net448),
    .B1(net436),
    .B2(\tms1x00.ins_pla_ors[8][13] ),
    .X(_04949_));
 sky130_fd_sc_hd__a221o_1 _09916_ (.A1(\tms1x00.ins_pla_ors[8][0] ),
    .A2(net440),
    .B1(net426),
    .B2(\tms1x00.ins_pla_ors[8][23] ),
    .C1(_04949_),
    .X(_04950_));
 sky130_fd_sc_hd__or4_2 _09917_ (.A(_04944_),
    .B(_04946_),
    .C(_04948_),
    .D(_04950_),
    .X(_04951_));
 sky130_fd_sc_hd__a22o_1 _09918_ (.A1(\tms1x00.ins_pla_ors[8][1] ),
    .A2(net434),
    .B1(net408),
    .B2(\tms1x00.ins_pla_ors[8][14] ),
    .X(_04952_));
 sky130_fd_sc_hd__a221o_1 _09919_ (.A1(\tms1x00.ins_pla_ors[8][3] ),
    .A2(net432),
    .B1(net406),
    .B2(\tms1x00.ins_pla_ors[8][19] ),
    .C1(_04952_),
    .X(_04953_));
 sky130_fd_sc_hd__a221o_1 _09920_ (.A1(\tms1x00.ins_pla_ors[8][17] ),
    .A2(net412),
    .B1(net404),
    .B2(\tms1x00.ins_pla_ors[8][25] ),
    .C1(_04953_),
    .X(_04954_));
 sky130_fd_sc_hd__a22o_1 _09921_ (.A1(\tms1x00.ins_pla_ors[8][4] ),
    .A2(net442),
    .B1(net438),
    .B2(\tms1x00.ins_pla_ors[8][2] ),
    .X(_04955_));
 sky130_fd_sc_hd__a221o_1 _09922_ (.A1(\tms1x00.ins_pla_ors[8][22] ),
    .A2(net416),
    .B1(net398),
    .B2(\tms1x00.ins_pla_ors[8][8] ),
    .C1(_04955_),
    .X(_04956_));
 sky130_fd_sc_hd__a22o_1 _09923_ (.A1(\tms1x00.ins_pla_ors[8][20] ),
    .A2(net452),
    .B1(net444),
    .B2(\tms1x00.ins_pla_ors[8][16] ),
    .X(_04957_));
 sky130_fd_sc_hd__a221o_1 _09924_ (.A1(\tms1x00.ins_pla_ors[8][27] ),
    .A2(net422),
    .B1(net400),
    .B2(\tms1x00.ins_pla_ors[8][6] ),
    .C1(_04957_),
    .X(_04958_));
 sky130_fd_sc_hd__or4_4 _09925_ (.A(_04951_),
    .B(_04954_),
    .C(_04956_),
    .D(_04958_),
    .X(_04959_));
 sky130_fd_sc_hd__o21ai_4 _09926_ (.A1(_04637_),
    .A2(_04959_),
    .B1(_04753_),
    .Y(_04960_));
 sky130_fd_sc_hd__a21o_1 _09927_ (.A1(_03384_),
    .A2(_04942_),
    .B1(_04960_),
    .X(_04961_));
 sky130_fd_sc_hd__o22a_1 _09928_ (.A1(\tms1x00.N[0] ),
    .A2(_04753_),
    .B1(_04924_),
    .B2(_04961_),
    .X(_01459_));
 sky130_fd_sc_hd__a21o_1 _09929_ (.A1(net7),
    .A2(_04923_),
    .B1(_04960_),
    .X(_04962_));
 sky130_fd_sc_hd__nor2_1 _09930_ (.A(\tms1x00.A[1] ),
    .B(_04903_),
    .Y(_04963_));
 sky130_fd_sc_hd__a221o_1 _09931_ (.A1(\tms1x00.A[1] ),
    .A2(_04885_),
    .B1(_04942_),
    .B2(_03390_),
    .C1(_04963_),
    .X(_04964_));
 sky130_fd_sc_hd__o22a_1 _09932_ (.A1(\tms1x00.N[1] ),
    .A2(_04753_),
    .B1(_04962_),
    .B2(_04964_),
    .X(_01460_));
 sky130_fd_sc_hd__nor2_1 _09933_ (.A(\tms1x00.A[2] ),
    .B(_04903_),
    .Y(_04965_));
 sky130_fd_sc_hd__a221o_1 _09934_ (.A1(\tms1x00.A[2] ),
    .A2(_04885_),
    .B1(_04923_),
    .B2(net8),
    .C1(_04965_),
    .X(_04966_));
 sky130_fd_sc_hd__a21o_1 _09935_ (.A1(_03396_),
    .A2(_04942_),
    .B1(_04960_),
    .X(_04967_));
 sky130_fd_sc_hd__o22a_1 _09936_ (.A1(\tms1x00.N[2] ),
    .A2(_04753_),
    .B1(_04966_),
    .B2(_04967_),
    .X(_01461_));
 sky130_fd_sc_hd__a21o_1 _09937_ (.A1(net9),
    .A2(_04923_),
    .B1(_04960_),
    .X(_04968_));
 sky130_fd_sc_hd__nor2_1 _09938_ (.A(\tms1x00.A[3] ),
    .B(_04903_),
    .Y(_04969_));
 sky130_fd_sc_hd__a221o_1 _09939_ (.A1(\tms1x00.A[3] ),
    .A2(_04885_),
    .B1(_04942_),
    .B2(_03402_),
    .C1(_04969_),
    .X(_04970_));
 sky130_fd_sc_hd__o22a_1 _09940_ (.A1(\tms1x00.N[3] ),
    .A2(_04753_),
    .B1(_04968_),
    .B2(_04970_),
    .X(_01462_));
 sky130_fd_sc_hd__a22o_1 _09941_ (.A1(\tms1x00.ins_pla_ors[13][3] ),
    .A2(net432),
    .B1(net404),
    .B2(\tms1x00.ins_pla_ors[13][25] ),
    .X(_04971_));
 sky130_fd_sc_hd__a22o_1 _09942_ (.A1(\tms1x00.ins_pla_ors[13][2] ),
    .A2(net438),
    .B1(net402),
    .B2(\tms1x00.ins_pla_ors[13][5] ),
    .X(_04972_));
 sky130_fd_sc_hd__a221o_1 _09943_ (.A1(\tms1x00.ins_pla_ors[13][23] ),
    .A2(net426),
    .B1(net422),
    .B2(\tms1x00.ins_pla_ors[13][27] ),
    .C1(_04972_),
    .X(_04973_));
 sky130_fd_sc_hd__a221o_1 _09944_ (.A1(\tms1x00.ins_pla_ors[13][18] ),
    .A2(net430),
    .B1(net410),
    .B2(\tms1x00.ins_pla_ors[13][15] ),
    .C1(_04971_),
    .X(_04974_));
 sky130_fd_sc_hd__a22o_1 _09945_ (.A1(\tms1x00.ins_pla_ors[13][7] ),
    .A2(net450),
    .B1(net398),
    .B2(\tms1x00.ins_pla_ors[13][8] ),
    .X(_04975_));
 sky130_fd_sc_hd__a22o_1 _09946_ (.A1(\tms1x00.ins_pla_ors[13][10] ),
    .A2(net420),
    .B1(net418),
    .B2(\tms1x00.ins_pla_ors[13][21] ),
    .X(_04976_));
 sky130_fd_sc_hd__a22o_1 _09947_ (.A1(\tms1x00.ins_pla_ors[13][11] ),
    .A2(net448),
    .B1(net406),
    .B2(\tms1x00.ins_pla_ors[13][19] ),
    .X(_04977_));
 sky130_fd_sc_hd__a221o_1 _09948_ (.A1(\tms1x00.ins_pla_ors[13][12] ),
    .A2(net424),
    .B1(net408),
    .B2(\tms1x00.ins_pla_ors[13][14] ),
    .C1(_04977_),
    .X(_04978_));
 sky130_fd_sc_hd__a22o_1 _09949_ (.A1(\tms1x00.ins_pla_ors[13][20] ),
    .A2(net452),
    .B1(net412),
    .B2(\tms1x00.ins_pla_ors[13][17] ),
    .X(_04979_));
 sky130_fd_sc_hd__a22o_1 _09950_ (.A1(\tms1x00.ins_pla_ors[13][16] ),
    .A2(net444),
    .B1(net414),
    .B2(\tms1x00.ins_pla_ors[13][9] ),
    .X(_04980_));
 sky130_fd_sc_hd__a221o_1 _09951_ (.A1(\tms1x00.ins_pla_ors[13][26] ),
    .A2(net454),
    .B1(net416),
    .B2(\tms1x00.ins_pla_ors[13][22] ),
    .C1(_04976_),
    .X(_04981_));
 sky130_fd_sc_hd__a221o_1 _09952_ (.A1(\tms1x00.ins_pla_ors[13][4] ),
    .A2(net442),
    .B1(net436),
    .B2(\tms1x00.ins_pla_ors[13][13] ),
    .C1(_04975_),
    .X(_04982_));
 sky130_fd_sc_hd__a221o_2 _09953_ (.A1(\tms1x00.ins_pla_ors[13][28] ),
    .A2(net446),
    .B1(net428),
    .B2(\tms1x00.ins_pla_ors[13][29] ),
    .C1(_04979_),
    .X(_04983_));
 sky130_fd_sc_hd__a221o_1 _09954_ (.A1(\tms1x00.ins_pla_ors[13][0] ),
    .A2(net440),
    .B1(net434),
    .B2(\tms1x00.ins_pla_ors[13][1] ),
    .C1(_04980_),
    .X(_04984_));
 sky130_fd_sc_hd__or4_2 _09955_ (.A(_04981_),
    .B(_04982_),
    .C(_04983_),
    .D(_04984_),
    .X(_04985_));
 sky130_fd_sc_hd__a22o_1 _09956_ (.A1(\tms1x00.ins_pla_ors[13][24] ),
    .A2(net456),
    .B1(net400),
    .B2(\tms1x00.ins_pla_ors[13][6] ),
    .X(_04986_));
 sky130_fd_sc_hd__or4_2 _09957_ (.A(_04973_),
    .B(_04974_),
    .C(_04978_),
    .D(_04986_),
    .X(_04987_));
 sky130_fd_sc_hd__nor2_4 _09958_ (.A(_04985_),
    .B(_04987_),
    .Y(_04988_));
 sky130_fd_sc_hd__nor3_4 _09959_ (.A(net592),
    .B(net340),
    .C(_04988_),
    .Y(_04989_));
 sky130_fd_sc_hd__mux2_1 _09960_ (.A0(\tms1x00.A[0] ),
    .A1(_04856_),
    .S(_04989_),
    .X(_01463_));
 sky130_fd_sc_hd__mux2_1 _09961_ (.A0(\tms1x00.A[1] ),
    .A1(_04858_),
    .S(_04989_),
    .X(_01464_));
 sky130_fd_sc_hd__mux2_1 _09962_ (.A0(\tms1x00.A[2] ),
    .A1(_04860_),
    .S(_04989_),
    .X(_01465_));
 sky130_fd_sc_hd__nor2_1 _09963_ (.A(\tms1x00.A[3] ),
    .B(_04989_),
    .Y(_04990_));
 sky130_fd_sc_hd__a21oi_1 _09964_ (.A1(_04863_),
    .A2(_04989_),
    .B1(_04990_),
    .Y(_01466_));
 sky130_fd_sc_hd__or3_4 _09965_ (.A(net611),
    .B(net361),
    .C(net710),
    .X(_04991_));
 sky130_fd_sc_hd__mux2_1 _09966_ (.A0(net976),
    .A1(\tms1x00.O_pla_ands[30][0] ),
    .S(_04991_),
    .X(_01467_));
 sky130_fd_sc_hd__mux2_1 _09967_ (.A0(net927),
    .A1(\tms1x00.O_pla_ands[30][1] ),
    .S(_04991_),
    .X(_01468_));
 sky130_fd_sc_hd__mux2_1 _09968_ (.A0(net1063),
    .A1(\tms1x00.O_pla_ands[30][2] ),
    .S(_04991_),
    .X(_01469_));
 sky130_fd_sc_hd__mux2_1 _09969_ (.A0(net1054),
    .A1(\tms1x00.O_pla_ands[30][3] ),
    .S(_04991_),
    .X(_01470_));
 sky130_fd_sc_hd__mux2_1 _09970_ (.A0(net1046),
    .A1(\tms1x00.O_pla_ands[30][4] ),
    .S(_04991_),
    .X(_01471_));
 sky130_fd_sc_hd__mux2_1 _09971_ (.A0(net1039),
    .A1(\tms1x00.O_pla_ands[30][5] ),
    .S(_04991_),
    .X(_01472_));
 sky130_fd_sc_hd__mux2_1 _09972_ (.A0(net1032),
    .A1(\tms1x00.O_pla_ands[30][6] ),
    .S(_04991_),
    .X(_01473_));
 sky130_fd_sc_hd__mux2_1 _09973_ (.A0(net1024),
    .A1(\tms1x00.O_pla_ands[30][7] ),
    .S(_04991_),
    .X(_01474_));
 sky130_fd_sc_hd__mux2_1 _09974_ (.A0(net1016),
    .A1(\tms1x00.O_pla_ands[30][8] ),
    .S(_04991_),
    .X(_01475_));
 sky130_fd_sc_hd__mux2_1 _09975_ (.A0(net1008),
    .A1(\tms1x00.O_pla_ands[30][9] ),
    .S(_04991_),
    .X(_01476_));
 sky130_fd_sc_hd__and3_4 _09976_ (.A(net820),
    .B(net359),
    .C(net709),
    .X(_04992_));
 sky130_fd_sc_hd__or3_4 _09977_ (.A(net813),
    .B(net357),
    .C(net706),
    .X(_04993_));
 sky130_fd_sc_hd__a21o_1 _09978_ (.A1(net981),
    .A2(_04992_),
    .B1(net558),
    .X(_04994_));
 sky130_fd_sc_hd__a21o_1 _09979_ (.A1(\tms1x00.O_pla_ands[4][0] ),
    .A2(_04993_),
    .B1(_04994_),
    .X(_01477_));
 sky130_fd_sc_hd__or2_1 _09980_ (.A(\tms1x00.O_pla_ands[4][1] ),
    .B(_04992_),
    .X(_04995_));
 sky130_fd_sc_hd__o211a_1 _09981_ (.A1(net933),
    .A2(_04993_),
    .B1(_04995_),
    .C1(net494),
    .X(_01478_));
 sky130_fd_sc_hd__a21o_1 _09982_ (.A1(net1069),
    .A2(_04992_),
    .B1(net559),
    .X(_04996_));
 sky130_fd_sc_hd__a21o_1 _09983_ (.A1(\tms1x00.O_pla_ands[4][2] ),
    .A2(_04993_),
    .B1(_04996_),
    .X(_01479_));
 sky130_fd_sc_hd__or2_1 _09984_ (.A(\tms1x00.O_pla_ands[4][3] ),
    .B(_04992_),
    .X(_04997_));
 sky130_fd_sc_hd__o211a_1 _09985_ (.A1(net1059),
    .A2(_04993_),
    .B1(_04997_),
    .C1(net494),
    .X(_01480_));
 sky130_fd_sc_hd__or2_1 _09986_ (.A(\tms1x00.O_pla_ands[4][4] ),
    .B(_04992_),
    .X(_04998_));
 sky130_fd_sc_hd__o211a_1 _09987_ (.A1(net1051),
    .A2(_04993_),
    .B1(_04998_),
    .C1(net496),
    .X(_01481_));
 sky130_fd_sc_hd__a21o_1 _09988_ (.A1(net1043),
    .A2(_04992_),
    .B1(net559),
    .X(_04999_));
 sky130_fd_sc_hd__a21o_1 _09989_ (.A1(\tms1x00.O_pla_ands[4][5] ),
    .A2(_04993_),
    .B1(_04999_),
    .X(_01482_));
 sky130_fd_sc_hd__a21o_1 _09990_ (.A1(net1036),
    .A2(_04992_),
    .B1(net560),
    .X(_05000_));
 sky130_fd_sc_hd__a21o_1 _09991_ (.A1(\tms1x00.O_pla_ands[4][6] ),
    .A2(_04993_),
    .B1(_05000_),
    .X(_01483_));
 sky130_fd_sc_hd__or2_1 _09992_ (.A(\tms1x00.O_pla_ands[4][7] ),
    .B(_04992_),
    .X(_05001_));
 sky130_fd_sc_hd__o211a_1 _09993_ (.A1(net1028),
    .A2(_04993_),
    .B1(_05001_),
    .C1(net496),
    .X(_01484_));
 sky130_fd_sc_hd__or2_1 _09994_ (.A(\tms1x00.O_pla_ands[4][8] ),
    .B(_04992_),
    .X(_05002_));
 sky130_fd_sc_hd__o211a_1 _09995_ (.A1(net1019),
    .A2(_04993_),
    .B1(_05002_),
    .C1(net494),
    .X(_01485_));
 sky130_fd_sc_hd__a21o_1 _09996_ (.A1(net1012),
    .A2(_04992_),
    .B1(net558),
    .X(_05003_));
 sky130_fd_sc_hd__a21o_1 _09997_ (.A1(\tms1x00.O_pla_ands[4][9] ),
    .A2(_04993_),
    .B1(_05003_),
    .X(_01486_));
 sky130_fd_sc_hd__or3_4 _09998_ (.A(net884),
    .B(net361),
    .C(net710),
    .X(_05004_));
 sky130_fd_sc_hd__mux2_1 _09999_ (.A0(net976),
    .A1(\tms1x00.O_pla_ands[29][0] ),
    .S(_05004_),
    .X(_01487_));
 sky130_fd_sc_hd__mux2_1 _10000_ (.A0(net927),
    .A1(\tms1x00.O_pla_ands[29][1] ),
    .S(_05004_),
    .X(_01488_));
 sky130_fd_sc_hd__mux2_1 _10001_ (.A0(net1063),
    .A1(\tms1x00.O_pla_ands[29][2] ),
    .S(_05004_),
    .X(_01489_));
 sky130_fd_sc_hd__mux2_1 _10002_ (.A0(net1054),
    .A1(\tms1x00.O_pla_ands[29][3] ),
    .S(_05004_),
    .X(_01490_));
 sky130_fd_sc_hd__mux2_1 _10003_ (.A0(net1046),
    .A1(\tms1x00.O_pla_ands[29][4] ),
    .S(_05004_),
    .X(_01491_));
 sky130_fd_sc_hd__mux2_1 _10004_ (.A0(net1038),
    .A1(\tms1x00.O_pla_ands[29][5] ),
    .S(_05004_),
    .X(_01492_));
 sky130_fd_sc_hd__mux2_1 _10005_ (.A0(net1030),
    .A1(\tms1x00.O_pla_ands[29][6] ),
    .S(_05004_),
    .X(_01493_));
 sky130_fd_sc_hd__mux2_1 _10006_ (.A0(net1024),
    .A1(\tms1x00.O_pla_ands[29][7] ),
    .S(_05004_),
    .X(_01494_));
 sky130_fd_sc_hd__mux2_1 _10007_ (.A0(net1016),
    .A1(\tms1x00.O_pla_ands[29][8] ),
    .S(_05004_),
    .X(_01495_));
 sky130_fd_sc_hd__mux2_1 _10008_ (.A0(net1007),
    .A1(\tms1x00.O_pla_ands[29][9] ),
    .S(_05004_),
    .X(_01496_));
 sky130_fd_sc_hd__nor2_2 _10009_ (.A(net745),
    .B(net355),
    .Y(_05005_));
 sky130_fd_sc_hd__or2_4 _10010_ (.A(net746),
    .B(net356),
    .X(_05006_));
 sky130_fd_sc_hd__mux2_1 _10011_ (.A0(net982),
    .A1(\tms1x00.ins_pla_ors[9][0] ),
    .S(_05006_),
    .X(_05007_));
 sky130_fd_sc_hd__or2_1 _10012_ (.A(net540),
    .B(_05007_),
    .X(_01497_));
 sky130_fd_sc_hd__mux2_1 _10013_ (.A0(net934),
    .A1(\tms1x00.ins_pla_ors[9][1] ),
    .S(net237),
    .X(_05008_));
 sky130_fd_sc_hd__or2_1 _10014_ (.A(net540),
    .B(_05008_),
    .X(_01498_));
 sky130_fd_sc_hd__mux2_1 _10015_ (.A0(net1070),
    .A1(\tms1x00.ins_pla_ors[9][2] ),
    .S(net237),
    .X(_05009_));
 sky130_fd_sc_hd__or2_1 _10016_ (.A(net540),
    .B(_05009_),
    .X(_01499_));
 sky130_fd_sc_hd__mux2_1 _10017_ (.A0(net1053),
    .A1(\tms1x00.ins_pla_ors[9][4] ),
    .S(net237),
    .X(_05010_));
 sky130_fd_sc_hd__or2_1 _10018_ (.A(net543),
    .B(_05010_),
    .X(_01500_));
 sky130_fd_sc_hd__mux2_1 _10019_ (.A0(net1044),
    .A1(\tms1x00.ins_pla_ors[9][5] ),
    .S(net237),
    .X(_05011_));
 sky130_fd_sc_hd__or2_1 _10020_ (.A(net543),
    .B(_05011_),
    .X(_01501_));
 sky130_fd_sc_hd__mux2_1 _10021_ (.A0(net1037),
    .A1(\tms1x00.ins_pla_ors[9][6] ),
    .S(net237),
    .X(_05012_));
 sky130_fd_sc_hd__or2_1 _10022_ (.A(net539),
    .B(_05012_),
    .X(_01502_));
 sky130_fd_sc_hd__mux2_1 _10023_ (.A0(net1029),
    .A1(\tms1x00.ins_pla_ors[9][7] ),
    .S(_05006_),
    .X(_05013_));
 sky130_fd_sc_hd__or2_1 _10024_ (.A(net540),
    .B(_05013_),
    .X(_01503_));
 sky130_fd_sc_hd__mux2_1 _10025_ (.A0(net1022),
    .A1(\tms1x00.ins_pla_ors[9][8] ),
    .S(_05006_),
    .X(_05014_));
 sky130_fd_sc_hd__or2_1 _10026_ (.A(net540),
    .B(_05014_),
    .X(_01504_));
 sky130_fd_sc_hd__nor2_2 _10027_ (.A(net519),
    .B(net238),
    .Y(_05015_));
 sky130_fd_sc_hd__nand2_8 _10028_ (.A(net461),
    .B(net237),
    .Y(_05016_));
 sky130_fd_sc_hd__o22a_1 _10029_ (.A1(\tms1x00.ins_pla_ors[9][9] ),
    .A2(net238),
    .B1(_05015_),
    .B2(net365),
    .X(_01505_));
 sky130_fd_sc_hd__mux2_1 _10030_ (.A0(\tms1x00.ins_pla_ors[9][10] ),
    .A1(net972),
    .S(net238),
    .X(_05017_));
 sky130_fd_sc_hd__or2_1 _10031_ (.A(net519),
    .B(_05017_),
    .X(_01506_));
 sky130_fd_sc_hd__mux2_1 _10032_ (.A0(\tms1x00.ins_pla_ors[9][11] ),
    .A1(net968),
    .S(net238),
    .X(_05018_));
 sky130_fd_sc_hd__or2_1 _10033_ (.A(net519),
    .B(_05018_),
    .X(_01507_));
 sky130_fd_sc_hd__mux2_1 _10034_ (.A0(\tms1x00.ins_pla_ors[9][12] ),
    .A1(net965),
    .S(net238),
    .X(_05019_));
 sky130_fd_sc_hd__or2_1 _10035_ (.A(net519),
    .B(_05019_),
    .X(_01508_));
 sky130_fd_sc_hd__mux2_1 _10036_ (.A0(\tms1x00.ins_pla_ors[9][13] ),
    .A1(net960),
    .S(net238),
    .X(_05020_));
 sky130_fd_sc_hd__or2_1 _10037_ (.A(net519),
    .B(_05020_),
    .X(_01509_));
 sky130_fd_sc_hd__mux2_1 _10038_ (.A0(\tms1x00.ins_pla_ors[9][14] ),
    .A1(net953),
    .S(net238),
    .X(_05021_));
 sky130_fd_sc_hd__or2_1 _10039_ (.A(net519),
    .B(_05021_),
    .X(_01510_));
 sky130_fd_sc_hd__a22o_1 _10040_ (.A1(\tms1x00.ins_pla_ors[9][15] ),
    .A2(net237),
    .B1(_05016_),
    .B2(_03530_),
    .X(_01511_));
 sky130_fd_sc_hd__a22o_1 _10041_ (.A1(\tms1x00.ins_pla_ors[9][16] ),
    .A2(net237),
    .B1(_05016_),
    .B2(_03440_),
    .X(_01512_));
 sky130_fd_sc_hd__mux2_1 _10042_ (.A0(\tms1x00.ins_pla_ors[9][17] ),
    .A1(net940),
    .S(net239),
    .X(_05022_));
 sky130_fd_sc_hd__or2_1 _10043_ (.A(net538),
    .B(_05022_),
    .X(_01513_));
 sky130_fd_sc_hd__a22o_1 _10044_ (.A1(\tms1x00.ins_pla_ors[9][18] ),
    .A2(net237),
    .B1(_05016_),
    .B2(_03444_),
    .X(_01514_));
 sky130_fd_sc_hd__mux2_1 _10045_ (.A0(\tms1x00.ins_pla_ors[9][19] ),
    .A1(net937),
    .S(net238),
    .X(_05023_));
 sky130_fd_sc_hd__or2_1 _10046_ (.A(net520),
    .B(_05023_),
    .X(_01515_));
 sky130_fd_sc_hd__mux2_1 _10047_ (.A0(\tms1x00.ins_pla_ors[9][20] ),
    .A1(net1078),
    .S(net239),
    .X(_05024_));
 sky130_fd_sc_hd__or2_1 _10048_ (.A(net537),
    .B(_05024_),
    .X(_01516_));
 sky130_fd_sc_hd__mux2_1 _10049_ (.A0(\tms1x00.ins_pla_ors[9][21] ),
    .A1(net1077),
    .S(net238),
    .X(_05025_));
 sky130_fd_sc_hd__or2_1 _10050_ (.A(net520),
    .B(_05025_),
    .X(_01517_));
 sky130_fd_sc_hd__mux2_1 _10051_ (.A0(\tms1x00.ins_pla_ors[9][22] ),
    .A1(net1075),
    .S(net238),
    .X(_05026_));
 sky130_fd_sc_hd__or2_1 _10052_ (.A(net537),
    .B(_05026_),
    .X(_01518_));
 sky130_fd_sc_hd__mux2_1 _10053_ (.A0(\tms1x00.ins_pla_ors[9][23] ),
    .A1(net1074),
    .S(net239),
    .X(_05027_));
 sky130_fd_sc_hd__or2_1 _10054_ (.A(net537),
    .B(_05027_),
    .X(_01519_));
 sky130_fd_sc_hd__mux2_1 _10055_ (.A0(\tms1x00.ins_pla_ors[9][24] ),
    .A1(net1073),
    .S(net239),
    .X(_05028_));
 sky130_fd_sc_hd__or2_1 _10056_ (.A(net539),
    .B(_05028_),
    .X(_01520_));
 sky130_fd_sc_hd__mux2_1 _10057_ (.A0(\tms1x00.ins_pla_ors[9][25] ),
    .A1(net105),
    .S(net239),
    .X(_05029_));
 sky130_fd_sc_hd__or2_1 _10058_ (.A(net537),
    .B(_05029_),
    .X(_01521_));
 sky130_fd_sc_hd__a22o_1 _10059_ (.A1(\tms1x00.ins_pla_ors[9][26] ),
    .A2(net237),
    .B1(_05016_),
    .B2(_03447_),
    .X(_01522_));
 sky130_fd_sc_hd__o22a_1 _10060_ (.A1(\tms1x00.ins_pla_ors[9][28] ),
    .A2(net239),
    .B1(_05015_),
    .B2(_03449_),
    .X(_01523_));
 sky130_fd_sc_hd__or3_4 _10061_ (.A(net855),
    .B(net361),
    .C(net710),
    .X(_05030_));
 sky130_fd_sc_hd__mux2_1 _10062_ (.A0(net978),
    .A1(\tms1x00.O_pla_ands[27][0] ),
    .S(_05030_),
    .X(_01524_));
 sky130_fd_sc_hd__mux2_1 _10063_ (.A0(net927),
    .A1(\tms1x00.O_pla_ands[27][1] ),
    .S(_05030_),
    .X(_01525_));
 sky130_fd_sc_hd__mux2_1 _10064_ (.A0(net1063),
    .A1(\tms1x00.O_pla_ands[27][2] ),
    .S(_05030_),
    .X(_01526_));
 sky130_fd_sc_hd__mux2_1 _10065_ (.A0(net1054),
    .A1(\tms1x00.O_pla_ands[27][3] ),
    .S(_05030_),
    .X(_01527_));
 sky130_fd_sc_hd__mux2_1 _10066_ (.A0(net1046),
    .A1(\tms1x00.O_pla_ands[27][4] ),
    .S(_05030_),
    .X(_01528_));
 sky130_fd_sc_hd__mux2_1 _10067_ (.A0(net1038),
    .A1(\tms1x00.O_pla_ands[27][5] ),
    .S(_05030_),
    .X(_01529_));
 sky130_fd_sc_hd__mux2_1 _10068_ (.A0(net1030),
    .A1(\tms1x00.O_pla_ands[27][6] ),
    .S(_05030_),
    .X(_01530_));
 sky130_fd_sc_hd__mux2_1 _10069_ (.A0(net1024),
    .A1(\tms1x00.O_pla_ands[27][7] ),
    .S(_05030_),
    .X(_01531_));
 sky130_fd_sc_hd__mux2_1 _10070_ (.A0(net1016),
    .A1(\tms1x00.O_pla_ands[27][8] ),
    .S(_05030_),
    .X(_01532_));
 sky130_fd_sc_hd__mux2_1 _10071_ (.A0(net1007),
    .A1(\tms1x00.O_pla_ands[27][9] ),
    .S(_05030_),
    .X(_01533_));
 sky130_fd_sc_hd__or3_4 _10072_ (.A(net804),
    .B(net361),
    .C(net710),
    .X(_05031_));
 sky130_fd_sc_hd__mux2_1 _10073_ (.A0(net978),
    .A1(\tms1x00.O_pla_ands[28][0] ),
    .S(_05031_),
    .X(_01534_));
 sky130_fd_sc_hd__mux2_1 _10074_ (.A0(net927),
    .A1(\tms1x00.O_pla_ands[28][1] ),
    .S(_05031_),
    .X(_01535_));
 sky130_fd_sc_hd__mux2_1 _10075_ (.A0(net1063),
    .A1(\tms1x00.O_pla_ands[28][2] ),
    .S(_05031_),
    .X(_01536_));
 sky130_fd_sc_hd__mux2_1 _10076_ (.A0(net1054),
    .A1(\tms1x00.O_pla_ands[28][3] ),
    .S(_05031_),
    .X(_01537_));
 sky130_fd_sc_hd__mux2_1 _10077_ (.A0(net1046),
    .A1(\tms1x00.O_pla_ands[28][4] ),
    .S(_05031_),
    .X(_01538_));
 sky130_fd_sc_hd__mux2_1 _10078_ (.A0(net1038),
    .A1(\tms1x00.O_pla_ands[28][5] ),
    .S(_05031_),
    .X(_01539_));
 sky130_fd_sc_hd__mux2_1 _10079_ (.A0(net1030),
    .A1(\tms1x00.O_pla_ands[28][6] ),
    .S(_05031_),
    .X(_01540_));
 sky130_fd_sc_hd__mux2_1 _10080_ (.A0(net1024),
    .A1(\tms1x00.O_pla_ands[28][7] ),
    .S(_05031_),
    .X(_01541_));
 sky130_fd_sc_hd__mux2_1 _10081_ (.A0(net1016),
    .A1(\tms1x00.O_pla_ands[28][8] ),
    .S(_05031_),
    .X(_01542_));
 sky130_fd_sc_hd__mux2_1 _10082_ (.A0(net1007),
    .A1(\tms1x00.O_pla_ands[28][9] ),
    .S(_05031_),
    .X(_01543_));
 sky130_fd_sc_hd__mux2_1 _10083_ (.A0(\tms1x00.ins_pla_ors[9][3] ),
    .A1(_03534_),
    .S(_05016_),
    .X(_01544_));
 sky130_fd_sc_hd__mux2_1 _10084_ (.A0(\tms1x00.ins_pla_ors[9][27] ),
    .A1(_03636_),
    .S(_05016_),
    .X(_01545_));
 sky130_fd_sc_hd__mux2_1 _10085_ (.A0(\tms1x00.ins_pla_ors[9][29] ),
    .A1(_03452_),
    .S(_05016_),
    .X(_01546_));
 sky130_fd_sc_hd__and3_4 _10086_ (.A(net849),
    .B(net359),
    .C(net708),
    .X(_05032_));
 sky130_fd_sc_hd__or3_4 _10087_ (.A(net834),
    .B(net357),
    .C(net707),
    .X(_05033_));
 sky130_fd_sc_hd__a21o_1 _10088_ (.A1(net977),
    .A2(_05032_),
    .B1(net532),
    .X(_05034_));
 sky130_fd_sc_hd__a21o_1 _10089_ (.A1(\tms1x00.O_pla_ands[0][0] ),
    .A2(_05033_),
    .B1(_05034_),
    .X(_01547_));
 sky130_fd_sc_hd__or2_1 _10090_ (.A(\tms1x00.O_pla_ands[0][1] ),
    .B(_05032_),
    .X(_05035_));
 sky130_fd_sc_hd__o211a_1 _10091_ (.A1(net929),
    .A2(_05033_),
    .B1(_05035_),
    .C1(net476),
    .X(_01548_));
 sky130_fd_sc_hd__a21o_1 _10092_ (.A1(net1071),
    .A2(_05032_),
    .B1(net532),
    .X(_05036_));
 sky130_fd_sc_hd__a21o_1 _10093_ (.A1(\tms1x00.O_pla_ands[0][2] ),
    .A2(_05033_),
    .B1(_05036_),
    .X(_01549_));
 sky130_fd_sc_hd__or2_1 _10094_ (.A(\tms1x00.O_pla_ands[0][3] ),
    .B(_05032_),
    .X(_05037_));
 sky130_fd_sc_hd__o211a_1 _10095_ (.A1(net1057),
    .A2(_05033_),
    .B1(_05037_),
    .C1(net476),
    .X(_01550_));
 sky130_fd_sc_hd__a21o_1 _10096_ (.A1(net1048),
    .A2(_05032_),
    .B1(net532),
    .X(_05038_));
 sky130_fd_sc_hd__a21o_1 _10097_ (.A1(\tms1x00.O_pla_ands[0][4] ),
    .A2(_05033_),
    .B1(_05038_),
    .X(_01551_));
 sky130_fd_sc_hd__or2_1 _10098_ (.A(\tms1x00.O_pla_ands[0][5] ),
    .B(_05032_),
    .X(_05039_));
 sky130_fd_sc_hd__o211a_1 _10099_ (.A1(net1040),
    .A2(_05033_),
    .B1(_05039_),
    .C1(net476),
    .X(_01552_));
 sky130_fd_sc_hd__a21o_1 _10100_ (.A1(net1031),
    .A2(_05032_),
    .B1(net532),
    .X(_05040_));
 sky130_fd_sc_hd__a21o_1 _10101_ (.A1(\tms1x00.O_pla_ands[0][6] ),
    .A2(_05033_),
    .B1(_05040_),
    .X(_01553_));
 sky130_fd_sc_hd__or2_1 _10102_ (.A(\tms1x00.O_pla_ands[0][7] ),
    .B(_05032_),
    .X(_05041_));
 sky130_fd_sc_hd__o211a_1 _10103_ (.A1(net1025),
    .A2(_05033_),
    .B1(_05041_),
    .C1(net476),
    .X(_01554_));
 sky130_fd_sc_hd__or2_1 _10104_ (.A(\tms1x00.O_pla_ands[0][8] ),
    .B(_05032_),
    .X(_05042_));
 sky130_fd_sc_hd__o211a_1 _10105_ (.A1(net1017),
    .A2(_05033_),
    .B1(_05042_),
    .C1(net476),
    .X(_01555_));
 sky130_fd_sc_hd__a21o_1 _10106_ (.A1(net1009),
    .A2(_05032_),
    .B1(net532),
    .X(_05043_));
 sky130_fd_sc_hd__a21o_1 _10107_ (.A1(\tms1x00.O_pla_ands[0][9] ),
    .A2(_05033_),
    .B1(_05043_),
    .X(_01556_));
 sky130_fd_sc_hd__or3_4 _10108_ (.A(net830),
    .B(net361),
    .C(_03472_),
    .X(_05044_));
 sky130_fd_sc_hd__mux2_1 _10109_ (.A0(net978),
    .A1(\tms1x00.O_pla_ands[24][0] ),
    .S(_05044_),
    .X(_01557_));
 sky130_fd_sc_hd__mux2_1 _10110_ (.A0(net927),
    .A1(\tms1x00.O_pla_ands[24][1] ),
    .S(_05044_),
    .X(_01558_));
 sky130_fd_sc_hd__mux2_1 _10111_ (.A0(net1063),
    .A1(\tms1x00.O_pla_ands[24][2] ),
    .S(_05044_),
    .X(_01559_));
 sky130_fd_sc_hd__mux2_1 _10112_ (.A0(net1054),
    .A1(\tms1x00.O_pla_ands[24][3] ),
    .S(_05044_),
    .X(_01560_));
 sky130_fd_sc_hd__mux2_1 _10113_ (.A0(net1046),
    .A1(\tms1x00.O_pla_ands[24][4] ),
    .S(_05044_),
    .X(_01561_));
 sky130_fd_sc_hd__mux2_1 _10114_ (.A0(net1038),
    .A1(\tms1x00.O_pla_ands[24][5] ),
    .S(_05044_),
    .X(_01562_));
 sky130_fd_sc_hd__mux2_1 _10115_ (.A0(net1030),
    .A1(\tms1x00.O_pla_ands[24][6] ),
    .S(_05044_),
    .X(_01563_));
 sky130_fd_sc_hd__mux2_1 _10116_ (.A0(net1026),
    .A1(\tms1x00.O_pla_ands[24][7] ),
    .S(_05044_),
    .X(_01564_));
 sky130_fd_sc_hd__mux2_1 _10117_ (.A0(net1016),
    .A1(\tms1x00.O_pla_ands[24][8] ),
    .S(_05044_),
    .X(_01565_));
 sky130_fd_sc_hd__mux2_1 _10118_ (.A0(net1007),
    .A1(\tms1x00.O_pla_ands[24][9] ),
    .S(_05044_),
    .X(_01566_));
 sky130_fd_sc_hd__or3_2 _10119_ (.A(net771),
    .B(net348),
    .C(net710),
    .X(_05045_));
 sky130_fd_sc_hd__mux2_1 _10120_ (.A0(net979),
    .A1(\tms1x00.ins_pla_ands[31][0] ),
    .S(net236),
    .X(_01567_));
 sky130_fd_sc_hd__mux2_1 _10121_ (.A0(net930),
    .A1(\tms1x00.ins_pla_ands[31][1] ),
    .S(net235),
    .X(_01568_));
 sky130_fd_sc_hd__mux2_1 _10122_ (.A0(net1066),
    .A1(\tms1x00.ins_pla_ands[31][2] ),
    .S(net236),
    .X(_01569_));
 sky130_fd_sc_hd__mux2_1 _10123_ (.A0(net1058),
    .A1(\tms1x00.ins_pla_ands[31][3] ),
    .S(net235),
    .X(_01570_));
 sky130_fd_sc_hd__mux2_1 _10124_ (.A0(net1049),
    .A1(\tms1x00.ins_pla_ands[31][4] ),
    .S(net235),
    .X(_01571_));
 sky130_fd_sc_hd__mux2_1 _10125_ (.A0(net1041),
    .A1(\tms1x00.ins_pla_ands[31][5] ),
    .S(net236),
    .X(_01572_));
 sky130_fd_sc_hd__mux2_1 _10126_ (.A0(net1033),
    .A1(\tms1x00.ins_pla_ands[31][6] ),
    .S(net236),
    .X(_01573_));
 sky130_fd_sc_hd__mux2_1 _10127_ (.A0(net1026),
    .A1(\tms1x00.ins_pla_ands[31][7] ),
    .S(net235),
    .X(_01574_));
 sky130_fd_sc_hd__mux2_1 _10128_ (.A0(net1014),
    .A1(\tms1x00.ins_pla_ands[31][8] ),
    .S(net235),
    .X(_01575_));
 sky130_fd_sc_hd__mux2_1 _10129_ (.A0(net1010),
    .A1(\tms1x00.ins_pla_ands[31][9] ),
    .S(net235),
    .X(_01576_));
 sky130_fd_sc_hd__mux2_1 _10130_ (.A0(net972),
    .A1(\tms1x00.ins_pla_ands[31][10] ),
    .S(net236),
    .X(_01577_));
 sky130_fd_sc_hd__mux2_1 _10131_ (.A0(net968),
    .A1(\tms1x00.ins_pla_ands[31][11] ),
    .S(net235),
    .X(_01578_));
 sky130_fd_sc_hd__mux2_1 _10132_ (.A0(net963),
    .A1(\tms1x00.ins_pla_ands[31][12] ),
    .S(net235),
    .X(_01579_));
 sky130_fd_sc_hd__mux2_1 _10133_ (.A0(net960),
    .A1(\tms1x00.ins_pla_ands[31][13] ),
    .S(net235),
    .X(_01580_));
 sky130_fd_sc_hd__mux2_1 _10134_ (.A0(net953),
    .A1(\tms1x00.ins_pla_ands[31][14] ),
    .S(net236),
    .X(_01581_));
 sky130_fd_sc_hd__mux2_1 _10135_ (.A0(net944),
    .A1(\tms1x00.ins_pla_ands[31][15] ),
    .S(net235),
    .X(_01582_));
 sky130_fd_sc_hd__and3_4 _10136_ (.A(net768),
    .B(net360),
    .C(net708),
    .X(_05046_));
 sky130_fd_sc_hd__or3_4 _10137_ (.A(net752),
    .B(net357),
    .C(net706),
    .X(_05047_));
 sky130_fd_sc_hd__or2_1 _10138_ (.A(\tms1x00.O_pla_ands[1][0] ),
    .B(_05046_),
    .X(_05048_));
 sky130_fd_sc_hd__o211a_1 _10139_ (.A1(net978),
    .A2(_05047_),
    .B1(_05048_),
    .C1(net477),
    .X(_01583_));
 sky130_fd_sc_hd__a21o_1 _10140_ (.A1(net929),
    .A2(_05046_),
    .B1(net532),
    .X(_05049_));
 sky130_fd_sc_hd__a21o_1 _10141_ (.A1(\tms1x00.O_pla_ands[1][1] ),
    .A2(_05047_),
    .B1(_05049_),
    .X(_01584_));
 sky130_fd_sc_hd__a21o_1 _10142_ (.A1(net1071),
    .A2(_05046_),
    .B1(net532),
    .X(_05050_));
 sky130_fd_sc_hd__a21o_1 _10143_ (.A1(\tms1x00.O_pla_ands[1][2] ),
    .A2(_05047_),
    .B1(_05050_),
    .X(_01585_));
 sky130_fd_sc_hd__or2_1 _10144_ (.A(\tms1x00.O_pla_ands[1][3] ),
    .B(_05046_),
    .X(_05051_));
 sky130_fd_sc_hd__o211a_1 _10145_ (.A1(net1057),
    .A2(_05047_),
    .B1(_05051_),
    .C1(net476),
    .X(_01586_));
 sky130_fd_sc_hd__a21o_1 _10146_ (.A1(net1048),
    .A2(_05046_),
    .B1(net533),
    .X(_05052_));
 sky130_fd_sc_hd__a21o_1 _10147_ (.A1(\tms1x00.O_pla_ands[1][4] ),
    .A2(_05047_),
    .B1(_05052_),
    .X(_01587_));
 sky130_fd_sc_hd__or2_1 _10148_ (.A(\tms1x00.O_pla_ands[1][5] ),
    .B(_05046_),
    .X(_05053_));
 sky130_fd_sc_hd__o211a_1 _10149_ (.A1(net1040),
    .A2(_05047_),
    .B1(_05053_),
    .C1(net477),
    .X(_01588_));
 sky130_fd_sc_hd__a21o_1 _10150_ (.A1(net1031),
    .A2(_05046_),
    .B1(net533),
    .X(_05054_));
 sky130_fd_sc_hd__a21o_1 _10151_ (.A1(\tms1x00.O_pla_ands[1][6] ),
    .A2(_05047_),
    .B1(_05054_),
    .X(_01589_));
 sky130_fd_sc_hd__or2_1 _10152_ (.A(\tms1x00.O_pla_ands[1][7] ),
    .B(_05046_),
    .X(_05055_));
 sky130_fd_sc_hd__o211a_1 _10153_ (.A1(net1025),
    .A2(_05047_),
    .B1(_05055_),
    .C1(net477),
    .X(_01590_));
 sky130_fd_sc_hd__or2_1 _10154_ (.A(\tms1x00.O_pla_ands[1][8] ),
    .B(_05046_),
    .X(_05056_));
 sky130_fd_sc_hd__o211a_1 _10155_ (.A1(net1023),
    .A2(_05047_),
    .B1(_05056_),
    .C1(net476),
    .X(_01591_));
 sky130_fd_sc_hd__a21o_1 _10156_ (.A1(net1010),
    .A2(_05046_),
    .B1(net532),
    .X(_05057_));
 sky130_fd_sc_hd__a21o_1 _10157_ (.A1(\tms1x00.O_pla_ands[1][9] ),
    .A2(_05047_),
    .B1(_05057_),
    .X(_01592_));
 sky130_fd_sc_hd__and3_4 _10158_ (.A(net876),
    .B(net359),
    .C(net709),
    .X(_05058_));
 sky130_fd_sc_hd__or3_4 _10159_ (.A(net868),
    .B(_03357_),
    .C(net706),
    .X(_05059_));
 sky130_fd_sc_hd__or2_1 _10160_ (.A(\tms1x00.O_pla_ands[3][0] ),
    .B(_05058_),
    .X(_05060_));
 sky130_fd_sc_hd__o211a_1 _10161_ (.A1(net981),
    .A2(_05059_),
    .B1(_05060_),
    .C1(net497),
    .X(_01593_));
 sky130_fd_sc_hd__a21o_1 _10162_ (.A1(net933),
    .A2(_05058_),
    .B1(net563),
    .X(_05061_));
 sky130_fd_sc_hd__a21o_1 _10163_ (.A1(\tms1x00.O_pla_ands[3][1] ),
    .A2(_05059_),
    .B1(_05061_),
    .X(_01594_));
 sky130_fd_sc_hd__or2_1 _10164_ (.A(\tms1x00.O_pla_ands[3][2] ),
    .B(_05058_),
    .X(_05062_));
 sky130_fd_sc_hd__o211a_1 _10165_ (.A1(net1069),
    .A2(_05059_),
    .B1(_05062_),
    .C1(net495),
    .X(_01595_));
 sky130_fd_sc_hd__a21o_1 _10166_ (.A1(net1061),
    .A2(_05058_),
    .B1(net563),
    .X(_05063_));
 sky130_fd_sc_hd__a21o_1 _10167_ (.A1(\tms1x00.O_pla_ands[3][3] ),
    .A2(_05059_),
    .B1(_05063_),
    .X(_01596_));
 sky130_fd_sc_hd__a21o_1 _10168_ (.A1(net1051),
    .A2(_05058_),
    .B1(net560),
    .X(_05064_));
 sky130_fd_sc_hd__a21o_1 _10169_ (.A1(\tms1x00.O_pla_ands[3][4] ),
    .A2(_05059_),
    .B1(_05064_),
    .X(_01597_));
 sky130_fd_sc_hd__or2_1 _10170_ (.A(\tms1x00.O_pla_ands[3][5] ),
    .B(_05058_),
    .X(_05065_));
 sky130_fd_sc_hd__o211a_1 _10171_ (.A1(net1043),
    .A2(_05059_),
    .B1(_05065_),
    .C1(net495),
    .X(_01598_));
 sky130_fd_sc_hd__a21o_1 _10172_ (.A1(net1036),
    .A2(_05058_),
    .B1(net559),
    .X(_05066_));
 sky130_fd_sc_hd__a21o_1 _10173_ (.A1(\tms1x00.O_pla_ands[3][6] ),
    .A2(_05059_),
    .B1(_05066_),
    .X(_01599_));
 sky130_fd_sc_hd__or2_1 _10174_ (.A(\tms1x00.O_pla_ands[3][7] ),
    .B(_05058_),
    .X(_05067_));
 sky130_fd_sc_hd__o211a_1 _10175_ (.A1(net1028),
    .A2(_05059_),
    .B1(_05067_),
    .C1(net497),
    .X(_01600_));
 sky130_fd_sc_hd__or2_1 _10176_ (.A(\tms1x00.O_pla_ands[3][8] ),
    .B(_05058_),
    .X(_05068_));
 sky130_fd_sc_hd__o211a_1 _10177_ (.A1(net1023),
    .A2(_05059_),
    .B1(_05068_),
    .C1(net495),
    .X(_01601_));
 sky130_fd_sc_hd__a21o_1 _10178_ (.A1(net1012),
    .A2(_05058_),
    .B1(net559),
    .X(_05069_));
 sky130_fd_sc_hd__a21o_1 _10179_ (.A1(\tms1x00.O_pla_ands[3][9] ),
    .A2(_05059_),
    .B1(_05069_),
    .X(_01602_));
 sky130_fd_sc_hd__or3_4 _10180_ (.A(net885),
    .B(_03351_),
    .C(_03353_),
    .X(_05070_));
 sky130_fd_sc_hd__mux2_1 _10181_ (.A0(net978),
    .A1(\tms1x00.O_pla_ands[21][0] ),
    .S(_05070_),
    .X(_01603_));
 sky130_fd_sc_hd__mux2_1 _10182_ (.A0(net929),
    .A1(\tms1x00.O_pla_ands[21][1] ),
    .S(_05070_),
    .X(_01604_));
 sky130_fd_sc_hd__mux2_1 _10183_ (.A0(net1064),
    .A1(\tms1x00.O_pla_ands[21][2] ),
    .S(_05070_),
    .X(_01605_));
 sky130_fd_sc_hd__mux2_1 _10184_ (.A0(net1057),
    .A1(\tms1x00.O_pla_ands[21][3] ),
    .S(_05070_),
    .X(_01606_));
 sky130_fd_sc_hd__mux2_1 _10185_ (.A0(net1048),
    .A1(\tms1x00.O_pla_ands[21][4] ),
    .S(_05070_),
    .X(_01607_));
 sky130_fd_sc_hd__mux2_1 _10186_ (.A0(net1041),
    .A1(\tms1x00.O_pla_ands[21][5] ),
    .S(_05070_),
    .X(_01608_));
 sky130_fd_sc_hd__mux2_1 _10187_ (.A0(net1032),
    .A1(\tms1x00.O_pla_ands[21][6] ),
    .S(_05070_),
    .X(_01609_));
 sky130_fd_sc_hd__mux2_1 _10188_ (.A0(net1026),
    .A1(\tms1x00.O_pla_ands[21][7] ),
    .S(_05070_),
    .X(_01610_));
 sky130_fd_sc_hd__mux2_1 _10189_ (.A0(net1018),
    .A1(\tms1x00.O_pla_ands[21][8] ),
    .S(_05070_),
    .X(_01611_));
 sky130_fd_sc_hd__mux2_1 _10190_ (.A0(net1008),
    .A1(\tms1x00.O_pla_ands[21][9] ),
    .S(_05070_),
    .X(_01612_));
 sky130_fd_sc_hd__a31o_1 _10191_ (.A1(net648),
    .A2(_04568_),
    .A3(net242),
    .B1(net128),
    .X(_05071_));
 sky130_fd_sc_hd__o311a_1 _10192_ (.A1(net651),
    .A2(_04569_),
    .A3(net240),
    .B1(_05071_),
    .C1(net634),
    .X(_01613_));
 sky130_fd_sc_hd__dfxtp_1 _10193_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(_00037_),
    .Q(\tms1x00.O_pla_ands[18][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10194_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_00038_),
    .Q(\tms1x00.O_pla_ands[18][1] ));
 sky130_fd_sc_hd__dfxtp_1 _10195_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(_00039_),
    .Q(\tms1x00.O_pla_ands[18][2] ));
 sky130_fd_sc_hd__dfxtp_1 _10196_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(_00040_),
    .Q(\tms1x00.O_pla_ands[18][3] ));
 sky130_fd_sc_hd__dfxtp_1 _10197_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_00041_),
    .Q(\tms1x00.O_pla_ands[18][4] ));
 sky130_fd_sc_hd__dfxtp_1 _10198_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(_00042_),
    .Q(\tms1x00.O_pla_ands[18][5] ));
 sky130_fd_sc_hd__dfxtp_1 _10199_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_00043_),
    .Q(\tms1x00.O_pla_ands[18][6] ));
 sky130_fd_sc_hd__dfxtp_1 _10200_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_00044_),
    .Q(\tms1x00.O_pla_ands[18][7] ));
 sky130_fd_sc_hd__dfxtp_1 _10201_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_00045_),
    .Q(\tms1x00.O_pla_ands[18][8] ));
 sky130_fd_sc_hd__dfxtp_1 _10202_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_00046_),
    .Q(\tms1x00.O_pla_ands[18][9] ));
 sky130_fd_sc_hd__dfxtp_1 _10203_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_00047_),
    .Q(\tms1x00.O_pla_ands[20][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10204_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_00048_),
    .Q(\tms1x00.O_pla_ands[20][1] ));
 sky130_fd_sc_hd__dfxtp_1 _10205_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(_00049_),
    .Q(\tms1x00.O_pla_ands[20][2] ));
 sky130_fd_sc_hd__dfxtp_1 _10206_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_00050_),
    .Q(\tms1x00.O_pla_ands[20][3] ));
 sky130_fd_sc_hd__dfxtp_1 _10207_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_00051_),
    .Q(\tms1x00.O_pla_ands[20][4] ));
 sky130_fd_sc_hd__dfxtp_1 _10208_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(_00052_),
    .Q(\tms1x00.O_pla_ands[20][5] ));
 sky130_fd_sc_hd__dfxtp_1 _10209_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_00053_),
    .Q(\tms1x00.O_pla_ands[20][6] ));
 sky130_fd_sc_hd__dfxtp_1 _10210_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_00054_),
    .Q(\tms1x00.O_pla_ands[20][7] ));
 sky130_fd_sc_hd__dfxtp_1 _10211_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(_00055_),
    .Q(\tms1x00.O_pla_ands[20][8] ));
 sky130_fd_sc_hd__dfxtp_1 _10212_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_00056_),
    .Q(\tms1x00.O_pla_ands[20][9] ));
 sky130_fd_sc_hd__dfxtp_4 _10213_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_00001_),
    .Q(net145));
 sky130_fd_sc_hd__dfxtp_2 _10214_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_00004_),
    .Q(\tms1x00.wb_step ));
 sky130_fd_sc_hd__dfxtp_1 _10215_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_00003_),
    .Q(wb_rst_override));
 sky130_fd_sc_hd__dfxtp_4 _10216_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_00002_),
    .Q(\tms1x00.pla_override ));
 sky130_fd_sc_hd__dfxtp_1 _10217_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_00000_),
    .Q(chip_sel_override));
 sky130_fd_sc_hd__dfxtp_1 _10218_ (.CLK(clknet_leaf_99_wb_clk_i),
    .D(_00057_),
    .Q(net153));
 sky130_fd_sc_hd__dfxtp_1 _10219_ (.CLK(clknet_leaf_99_wb_clk_i),
    .D(_00058_),
    .Q(net154));
 sky130_fd_sc_hd__dfxtp_1 _10220_ (.CLK(clknet_leaf_81_wb_clk_i),
    .D(_00059_),
    .Q(net155));
 sky130_fd_sc_hd__dfxtp_2 _10221_ (.CLK(clknet_leaf_81_wb_clk_i),
    .D(_00060_),
    .Q(net156));
 sky130_fd_sc_hd__dfxtp_2 _10222_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_00005_),
    .Q(\wbs_o_buff[0] ));
 sky130_fd_sc_hd__dfxtp_2 _10223_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_00016_),
    .Q(\wbs_o_buff[1] ));
 sky130_fd_sc_hd__dfxtp_2 _10224_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_00027_),
    .Q(\wbs_o_buff[2] ));
 sky130_fd_sc_hd__dfxtp_2 _10225_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_00030_),
    .Q(\wbs_o_buff[3] ));
 sky130_fd_sc_hd__dfxtp_2 _10226_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_00031_),
    .Q(\wbs_o_buff[4] ));
 sky130_fd_sc_hd__dfxtp_2 _10227_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_00032_),
    .Q(\wbs_o_buff[5] ));
 sky130_fd_sc_hd__dfxtp_2 _10228_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_00033_),
    .Q(\wbs_o_buff[6] ));
 sky130_fd_sc_hd__dfxtp_2 _10229_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_00034_),
    .Q(\wbs_o_buff[7] ));
 sky130_fd_sc_hd__dfxtp_2 _10230_ (.CLK(clknet_leaf_56_wb_clk_i),
    .D(_00035_),
    .Q(\wbs_o_buff[8] ));
 sky130_fd_sc_hd__dfxtp_2 _10231_ (.CLK(clknet_leaf_89_wb_clk_i),
    .D(_00036_),
    .Q(\wbs_o_buff[9] ));
 sky130_fd_sc_hd__dfxtp_2 _10232_ (.CLK(clknet_leaf_126_wb_clk_i),
    .D(_00006_),
    .Q(\wbs_o_buff[10] ));
 sky130_fd_sc_hd__dfxtp_2 _10233_ (.CLK(clknet_leaf_126_wb_clk_i),
    .D(_00007_),
    .Q(\wbs_o_buff[11] ));
 sky130_fd_sc_hd__dfxtp_2 _10234_ (.CLK(clknet_leaf_89_wb_clk_i),
    .D(_00008_),
    .Q(\wbs_o_buff[12] ));
 sky130_fd_sc_hd__dfxtp_2 _10235_ (.CLK(clknet_leaf_88_wb_clk_i),
    .D(_00009_),
    .Q(\wbs_o_buff[13] ));
 sky130_fd_sc_hd__dfxtp_2 _10236_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_00010_),
    .Q(\wbs_o_buff[14] ));
 sky130_fd_sc_hd__dfxtp_2 _10237_ (.CLK(clknet_leaf_126_wb_clk_i),
    .D(_00011_),
    .Q(\wbs_o_buff[15] ));
 sky130_fd_sc_hd__dfxtp_2 _10238_ (.CLK(clknet_leaf_91_wb_clk_i),
    .D(_00012_),
    .Q(\wbs_o_buff[16] ));
 sky130_fd_sc_hd__dfxtp_2 _10239_ (.CLK(clknet_leaf_87_wb_clk_i),
    .D(_00013_),
    .Q(\wbs_o_buff[17] ));
 sky130_fd_sc_hd__dfxtp_2 _10240_ (.CLK(clknet_leaf_87_wb_clk_i),
    .D(_00014_),
    .Q(\wbs_o_buff[18] ));
 sky130_fd_sc_hd__dfxtp_2 _10241_ (.CLK(clknet_leaf_83_wb_clk_i),
    .D(_00015_),
    .Q(\wbs_o_buff[19] ));
 sky130_fd_sc_hd__dfxtp_1 _10242_ (.CLK(clknet_leaf_114_wb_clk_i),
    .D(_00017_),
    .Q(\wbs_o_buff[20] ));
 sky130_fd_sc_hd__dfxtp_1 _10243_ (.CLK(clknet_leaf_113_wb_clk_i),
    .D(_00018_),
    .Q(\wbs_o_buff[21] ));
 sky130_fd_sc_hd__dfxtp_1 _10244_ (.CLK(clknet_leaf_114_wb_clk_i),
    .D(_00019_),
    .Q(\wbs_o_buff[22] ));
 sky130_fd_sc_hd__dfxtp_1 _10245_ (.CLK(clknet_leaf_113_wb_clk_i),
    .D(_00020_),
    .Q(\wbs_o_buff[23] ));
 sky130_fd_sc_hd__dfxtp_2 _10246_ (.CLK(clknet_leaf_93_wb_clk_i),
    .D(_00021_),
    .Q(\wbs_o_buff[24] ));
 sky130_fd_sc_hd__dfxtp_1 _10247_ (.CLK(clknet_leaf_113_wb_clk_i),
    .D(_00022_),
    .Q(\wbs_o_buff[25] ));
 sky130_fd_sc_hd__dfxtp_1 _10248_ (.CLK(clknet_leaf_114_wb_clk_i),
    .D(_00023_),
    .Q(\wbs_o_buff[26] ));
 sky130_fd_sc_hd__dfxtp_1 _10249_ (.CLK(clknet_leaf_113_wb_clk_i),
    .D(_00024_),
    .Q(\wbs_o_buff[27] ));
 sky130_fd_sc_hd__dfxtp_1 _10250_ (.CLK(clknet_leaf_110_wb_clk_i),
    .D(_00025_),
    .Q(\wbs_o_buff[28] ));
 sky130_fd_sc_hd__dfxtp_1 _10251_ (.CLK(clknet_leaf_114_wb_clk_i),
    .D(_00026_),
    .Q(\wbs_o_buff[29] ));
 sky130_fd_sc_hd__dfxtp_1 _10252_ (.CLK(clknet_leaf_114_wb_clk_i),
    .D(_00028_),
    .Q(\wbs_o_buff[30] ));
 sky130_fd_sc_hd__dfxtp_1 _10253_ (.CLK(clknet_leaf_114_wb_clk_i),
    .D(_00029_),
    .Q(\wbs_o_buff[31] ));
 sky130_fd_sc_hd__dfxtp_1 _10254_ (.CLK(clknet_leaf_137_wb_clk_i),
    .D(net1133),
    .Q(net179));
 sky130_fd_sc_hd__dfxtp_1 _10255_ (.CLK(clknet_leaf_137_wb_clk_i),
    .D(valid),
    .Q(feedback_delay));
 sky130_fd_sc_hd__dfxtp_1 _10256_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(_00061_),
    .Q(\tms1x00.O_pla_ands[19][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10257_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_00062_),
    .Q(\tms1x00.O_pla_ands[19][1] ));
 sky130_fd_sc_hd__dfxtp_1 _10258_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(_00063_),
    .Q(\tms1x00.O_pla_ands[19][2] ));
 sky130_fd_sc_hd__dfxtp_1 _10259_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(_00064_),
    .Q(\tms1x00.O_pla_ands[19][3] ));
 sky130_fd_sc_hd__dfxtp_1 _10260_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(_00065_),
    .Q(\tms1x00.O_pla_ands[19][4] ));
 sky130_fd_sc_hd__dfxtp_1 _10261_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_00066_),
    .Q(\tms1x00.O_pla_ands[19][5] ));
 sky130_fd_sc_hd__dfxtp_1 _10262_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_00067_),
    .Q(\tms1x00.O_pla_ands[19][6] ));
 sky130_fd_sc_hd__dfxtp_1 _10263_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_00068_),
    .Q(\tms1x00.O_pla_ands[19][7] ));
 sky130_fd_sc_hd__dfxtp_1 _10264_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_00069_),
    .Q(\tms1x00.O_pla_ands[19][8] ));
 sky130_fd_sc_hd__dfxtp_1 _10265_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(_00070_),
    .Q(\tms1x00.O_pla_ands[19][9] ));
 sky130_fd_sc_hd__dfxtp_1 _10266_ (.CLK(clknet_leaf_124_wb_clk_i),
    .D(_00071_),
    .Q(\tms1x00.ins_pla_ors[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _10267_ (.CLK(clknet_leaf_124_wb_clk_i),
    .D(_00072_),
    .Q(\tms1x00.ins_pla_ors[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _10268_ (.CLK(clknet_leaf_123_wb_clk_i),
    .D(_00073_),
    .Q(\tms1x00.ins_pla_ors[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _10269_ (.CLK(clknet_leaf_90_wb_clk_i),
    .D(_00074_),
    .Q(\tms1x00.ins_pla_ors[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 _10270_ (.CLK(clknet_leaf_125_wb_clk_i),
    .D(_00075_),
    .Q(\tms1x00.ins_pla_ors[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 _10271_ (.CLK(clknet_leaf_126_wb_clk_i),
    .D(_00076_),
    .Q(\tms1x00.ins_pla_ors[12][8] ));
 sky130_fd_sc_hd__dfxtp_1 _10272_ (.CLK(clknet_leaf_133_wb_clk_i),
    .D(_00077_),
    .Q(\tms1x00.ins_pla_ors[12][14] ));
 sky130_fd_sc_hd__dfxtp_1 _10273_ (.CLK(clknet_leaf_122_wb_clk_i),
    .D(_00078_),
    .Q(\tms1x00.ins_pla_ors[12][16] ));
 sky130_fd_sc_hd__dfxtp_1 _10274_ (.CLK(clknet_leaf_122_wb_clk_i),
    .D(_00079_),
    .Q(\tms1x00.ins_pla_ors[12][17] ));
 sky130_fd_sc_hd__dfxtp_1 _10275_ (.CLK(clknet_leaf_122_wb_clk_i),
    .D(_00080_),
    .Q(\tms1x00.ins_pla_ors[12][18] ));
 sky130_fd_sc_hd__dfxtp_1 _10276_ (.CLK(clknet_leaf_133_wb_clk_i),
    .D(_00081_),
    .Q(\tms1x00.ins_pla_ors[12][21] ));
 sky130_fd_sc_hd__dfxtp_1 _10277_ (.CLK(clknet_leaf_117_wb_clk_i),
    .D(_00082_),
    .Q(\tms1x00.ins_pla_ors[12][26] ));
 sky130_fd_sc_hd__dfxtp_1 _10278_ (.CLK(clknet_leaf_113_wb_clk_i),
    .D(_00083_),
    .Q(\tms1x00.ins_pla_ors[12][28] ));
 sky130_fd_sc_hd__dfxtp_1 _10279_ (.CLK(clknet_leaf_120_wb_clk_i),
    .D(_00084_),
    .Q(\tms1x00.ins_pla_ors[12][29] ));
 sky130_fd_sc_hd__dfxtp_2 _10280_ (.CLK(clknet_leaf_130_wb_clk_i),
    .D(_00085_),
    .Q(\tms1x00.ins_pla_ors[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10281_ (.CLK(clknet_leaf_127_wb_clk_i),
    .D(_00086_),
    .Q(\tms1x00.ins_pla_ors[14][1] ));
 sky130_fd_sc_hd__dfxtp_2 _10282_ (.CLK(clknet_leaf_130_wb_clk_i),
    .D(_00087_),
    .Q(\tms1x00.ins_pla_ors[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _10283_ (.CLK(clknet_leaf_125_wb_clk_i),
    .D(_00088_),
    .Q(\tms1x00.ins_pla_ors[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 _10284_ (.CLK(clknet_leaf_124_wb_clk_i),
    .D(_00089_),
    .Q(\tms1x00.ins_pla_ors[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 _10285_ (.CLK(clknet_leaf_129_wb_clk_i),
    .D(_00090_),
    .Q(\tms1x00.ins_pla_ors[14][7] ));
 sky130_fd_sc_hd__dfxtp_1 _10286_ (.CLK(clknet_leaf_129_wb_clk_i),
    .D(_00091_),
    .Q(\tms1x00.ins_pla_ors[14][8] ));
 sky130_fd_sc_hd__dfxtp_1 _10287_ (.CLK(clknet_leaf_129_wb_clk_i),
    .D(_00092_),
    .Q(\tms1x00.ins_pla_ors[14][9] ));
 sky130_fd_sc_hd__dfxtp_1 _10288_ (.CLK(clknet_leaf_133_wb_clk_i),
    .D(_00093_),
    .Q(\tms1x00.ins_pla_ors[14][10] ));
 sky130_fd_sc_hd__dfxtp_2 _10289_ (.CLK(clknet_leaf_129_wb_clk_i),
    .D(_00094_),
    .Q(\tms1x00.ins_pla_ors[14][11] ));
 sky130_fd_sc_hd__dfxtp_1 _10290_ (.CLK(clknet_leaf_134_wb_clk_i),
    .D(_00095_),
    .Q(\tms1x00.ins_pla_ors[14][14] ));
 sky130_fd_sc_hd__dfxtp_1 _10291_ (.CLK(clknet_leaf_116_wb_clk_i),
    .D(_00096_),
    .Q(\tms1x00.ins_pla_ors[14][15] ));
 sky130_fd_sc_hd__dfxtp_1 _10292_ (.CLK(clknet_leaf_120_wb_clk_i),
    .D(_00097_),
    .Q(\tms1x00.ins_pla_ors[14][17] ));
 sky130_fd_sc_hd__dfxtp_2 _10293_ (.CLK(clknet_leaf_115_wb_clk_i),
    .D(_00098_),
    .Q(\tms1x00.ins_pla_ors[14][18] ));
 sky130_fd_sc_hd__dfxtp_1 _10294_ (.CLK(clknet_leaf_128_wb_clk_i),
    .D(_00099_),
    .Q(\tms1x00.ins_pla_ors[14][19] ));
 sky130_fd_sc_hd__dfxtp_1 _10295_ (.CLK(clknet_leaf_114_wb_clk_i),
    .D(_00100_),
    .Q(\tms1x00.ins_pla_ors[14][20] ));
 sky130_fd_sc_hd__dfxtp_1 _10296_ (.CLK(clknet_leaf_135_wb_clk_i),
    .D(_00101_),
    .Q(\tms1x00.ins_pla_ors[14][21] ));
 sky130_fd_sc_hd__dfxtp_1 _10297_ (.CLK(clknet_leaf_124_wb_clk_i),
    .D(_00102_),
    .Q(\tms1x00.ins_pla_ors[14][24] ));
 sky130_fd_sc_hd__dfxtp_1 _10298_ (.CLK(clknet_leaf_116_wb_clk_i),
    .D(_00103_),
    .Q(\tms1x00.ins_pla_ors[14][26] ));
 sky130_fd_sc_hd__dfxtp_1 _10299_ (.CLK(clknet_leaf_120_wb_clk_i),
    .D(_00104_),
    .Q(\tms1x00.ins_pla_ors[14][28] ));
 sky130_fd_sc_hd__dfxtp_1 _10300_ (.CLK(clknet_leaf_130_wb_clk_i),
    .D(_00105_),
    .Q(\tms1x00.ins_pla_ands[26][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10301_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_00106_),
    .Q(\tms1x00.ins_pla_ands[26][2] ));
 sky130_fd_sc_hd__dfxtp_1 _10302_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_00107_),
    .Q(\tms1x00.ins_pla_ands[26][4] ));
 sky130_fd_sc_hd__dfxtp_1 _10303_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_00108_),
    .Q(\tms1x00.ins_pla_ands[26][6] ));
 sky130_fd_sc_hd__dfxtp_1 _10304_ (.CLK(clknet_leaf_139_wb_clk_i),
    .D(_00109_),
    .Q(\tms1x00.ins_pla_ands[26][8] ));
 sky130_fd_sc_hd__dfxtp_1 _10305_ (.CLK(clknet_leaf_138_wb_clk_i),
    .D(_00110_),
    .Q(\tms1x00.ins_pla_ands[26][9] ));
 sky130_fd_sc_hd__dfxtp_1 _10306_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_00111_),
    .Q(\tms1x00.ins_pla_ands[26][10] ));
 sky130_fd_sc_hd__dfxtp_1 _10307_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_00112_),
    .Q(\tms1x00.ins_pla_ands[26][11] ));
 sky130_fd_sc_hd__dfxtp_1 _10308_ (.CLK(clknet_leaf_131_wb_clk_i),
    .D(_00113_),
    .Q(\tms1x00.ins_pla_ands[26][12] ));
 sky130_fd_sc_hd__dfxtp_1 _10309_ (.CLK(clknet_leaf_139_wb_clk_i),
    .D(_00114_),
    .Q(\tms1x00.ins_pla_ands[26][13] ));
 sky130_fd_sc_hd__dfxtp_1 _10310_ (.CLK(clknet_leaf_131_wb_clk_i),
    .D(_00115_),
    .Q(\tms1x00.ins_pla_ors[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10311_ (.CLK(clknet_leaf_127_wb_clk_i),
    .D(_00116_),
    .Q(\tms1x00.ins_pla_ors[15][1] ));
 sky130_fd_sc_hd__dfxtp_2 _10312_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_00117_),
    .Q(\tms1x00.ins_pla_ors[15][2] ));
 sky130_fd_sc_hd__dfxtp_2 _10313_ (.CLK(clknet_leaf_129_wb_clk_i),
    .D(_00118_),
    .Q(\tms1x00.ins_pla_ors[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _10314_ (.CLK(clknet_leaf_129_wb_clk_i),
    .D(_00119_),
    .Q(\tms1x00.ins_pla_ors[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 _10315_ (.CLK(clknet_leaf_125_wb_clk_i),
    .D(_00120_),
    .Q(\tms1x00.ins_pla_ors[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 _10316_ (.CLK(clknet_leaf_118_wb_clk_i),
    .D(_00121_),
    .Q(\tms1x00.ins_pla_ors[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 _10317_ (.CLK(clknet_leaf_129_wb_clk_i),
    .D(_00122_),
    .Q(\tms1x00.ins_pla_ors[15][8] ));
 sky130_fd_sc_hd__dfxtp_2 _10318_ (.CLK(clknet_leaf_129_wb_clk_i),
    .D(_00123_),
    .Q(\tms1x00.ins_pla_ors[15][9] ));
 sky130_fd_sc_hd__dfxtp_1 _10319_ (.CLK(clknet_leaf_133_wb_clk_i),
    .D(_00124_),
    .Q(\tms1x00.ins_pla_ors[15][10] ));
 sky130_fd_sc_hd__dfxtp_1 _10320_ (.CLK(clknet_leaf_129_wb_clk_i),
    .D(_00125_),
    .Q(\tms1x00.ins_pla_ors[15][11] ));
 sky130_fd_sc_hd__dfxtp_1 _10321_ (.CLK(clknet_leaf_129_wb_clk_i),
    .D(_00126_),
    .Q(\tms1x00.ins_pla_ors[15][12] ));
 sky130_fd_sc_hd__dfxtp_1 _10322_ (.CLK(clknet_leaf_131_wb_clk_i),
    .D(_00127_),
    .Q(\tms1x00.ins_pla_ors[15][13] ));
 sky130_fd_sc_hd__dfxtp_1 _10323_ (.CLK(clknet_leaf_134_wb_clk_i),
    .D(_00128_),
    .Q(\tms1x00.ins_pla_ors[15][14] ));
 sky130_fd_sc_hd__dfxtp_1 _10324_ (.CLK(clknet_leaf_116_wb_clk_i),
    .D(_00129_),
    .Q(\tms1x00.ins_pla_ors[15][15] ));
 sky130_fd_sc_hd__dfxtp_2 _10325_ (.CLK(clknet_leaf_115_wb_clk_i),
    .D(_00130_),
    .Q(\tms1x00.ins_pla_ors[15][16] ));
 sky130_fd_sc_hd__dfxtp_2 _10326_ (.CLK(clknet_leaf_120_wb_clk_i),
    .D(_00131_),
    .Q(\tms1x00.ins_pla_ors[15][17] ));
 sky130_fd_sc_hd__dfxtp_2 _10327_ (.CLK(clknet_leaf_115_wb_clk_i),
    .D(_00132_),
    .Q(\tms1x00.ins_pla_ors[15][18] ));
 sky130_fd_sc_hd__dfxtp_1 _10328_ (.CLK(clknet_leaf_128_wb_clk_i),
    .D(_00133_),
    .Q(\tms1x00.ins_pla_ors[15][19] ));
 sky130_fd_sc_hd__dfxtp_1 _10329_ (.CLK(clknet_leaf_115_wb_clk_i),
    .D(_00134_),
    .Q(\tms1x00.ins_pla_ors[15][20] ));
 sky130_fd_sc_hd__dfxtp_1 _10330_ (.CLK(clknet_leaf_133_wb_clk_i),
    .D(_00135_),
    .Q(\tms1x00.ins_pla_ors[15][21] ));
 sky130_fd_sc_hd__dfxtp_1 _10331_ (.CLK(clknet_leaf_115_wb_clk_i),
    .D(_00136_),
    .Q(\tms1x00.ins_pla_ors[15][22] ));
 sky130_fd_sc_hd__dfxtp_1 _10332_ (.CLK(clknet_leaf_119_wb_clk_i),
    .D(_00137_),
    .Q(\tms1x00.ins_pla_ors[15][23] ));
 sky130_fd_sc_hd__dfxtp_1 _10333_ (.CLK(clknet_leaf_118_wb_clk_i),
    .D(_00138_),
    .Q(\tms1x00.ins_pla_ors[15][25] ));
 sky130_fd_sc_hd__dfxtp_1 _10334_ (.CLK(clknet_leaf_116_wb_clk_i),
    .D(_00139_),
    .Q(\tms1x00.ins_pla_ors[15][26] ));
 sky130_fd_sc_hd__dfxtp_1 _10335_ (.CLK(clknet_leaf_119_wb_clk_i),
    .D(_00140_),
    .Q(\tms1x00.ins_pla_ors[15][27] ));
 sky130_fd_sc_hd__dfxtp_1 _10336_ (.CLK(clknet_leaf_113_wb_clk_i),
    .D(_00141_),
    .Q(\tms1x00.ins_pla_ors[15][28] ));
 sky130_fd_sc_hd__dfxtp_1 _10337_ (.CLK(clknet_leaf_93_wb_clk_i),
    .D(_00142_),
    .Q(\tms1x00.ins_pla_ors[15][29] ));
 sky130_fd_sc_hd__dfxtp_1 _10338_ (.CLK(clknet_leaf_99_wb_clk_i),
    .D(_00143_),
    .Q(\tms1x00.ins_pla_ors[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10339_ (.CLK(clknet_leaf_93_wb_clk_i),
    .D(_00144_),
    .Q(\tms1x00.ins_pla_ors[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _10340_ (.CLK(clknet_leaf_96_wb_clk_i),
    .D(_00145_),
    .Q(\tms1x00.ins_pla_ors[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _10341_ (.CLK(clknet_leaf_92_wb_clk_i),
    .D(_00146_),
    .Q(\tms1x00.ins_pla_ors[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _10342_ (.CLK(clknet_leaf_91_wb_clk_i),
    .D(_00147_),
    .Q(\tms1x00.ins_pla_ors[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _10343_ (.CLK(clknet_leaf_96_wb_clk_i),
    .D(_00148_),
    .Q(\tms1x00.ins_pla_ors[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _10344_ (.CLK(clknet_leaf_100_wb_clk_i),
    .D(_00149_),
    .Q(\tms1x00.ins_pla_ors[4][9] ));
 sky130_fd_sc_hd__dfxtp_1 _10345_ (.CLK(clknet_leaf_99_wb_clk_i),
    .D(_00150_),
    .Q(\tms1x00.ins_pla_ors[4][10] ));
 sky130_fd_sc_hd__dfxtp_1 _10346_ (.CLK(clknet_leaf_110_wb_clk_i),
    .D(_00151_),
    .Q(\tms1x00.ins_pla_ors[4][12] ));
 sky130_fd_sc_hd__dfxtp_1 _10347_ (.CLK(clknet_leaf_92_wb_clk_i),
    .D(_00152_),
    .Q(\tms1x00.ins_pla_ors[4][13] ));
 sky130_fd_sc_hd__dfxtp_1 _10348_ (.CLK(clknet_leaf_112_wb_clk_i),
    .D(_00153_),
    .Q(\tms1x00.ins_pla_ors[4][15] ));
 sky130_fd_sc_hd__dfxtp_1 _10349_ (.CLK(clknet_leaf_101_wb_clk_i),
    .D(_00154_),
    .Q(\tms1x00.ins_pla_ors[4][19] ));
 sky130_fd_sc_hd__dfxtp_2 _10350_ (.CLK(clknet_leaf_106_wb_clk_i),
    .D(_00155_),
    .Q(\tms1x00.ins_pla_ors[4][20] ));
 sky130_fd_sc_hd__dfxtp_2 _10351_ (.CLK(clknet_leaf_109_wb_clk_i),
    .D(_00156_),
    .Q(\tms1x00.ins_pla_ors[4][21] ));
 sky130_fd_sc_hd__dfxtp_1 _10352_ (.CLK(clknet_leaf_110_wb_clk_i),
    .D(_00157_),
    .Q(\tms1x00.ins_pla_ors[4][22] ));
 sky130_fd_sc_hd__dfxtp_2 _10353_ (.CLK(clknet_leaf_100_wb_clk_i),
    .D(_00158_),
    .Q(\tms1x00.ins_pla_ors[4][23] ));
 sky130_fd_sc_hd__dfxtp_1 _10354_ (.CLK(clknet_leaf_127_wb_clk_i),
    .D(_00159_),
    .Q(\tms1x00.ins_pla_ors[15][7] ));
 sky130_fd_sc_hd__dfxtp_1 _10355_ (.CLK(clknet_leaf_124_wb_clk_i),
    .D(_00160_),
    .Q(\tms1x00.ins_pla_ors[15][24] ));
 sky130_fd_sc_hd__dfxtp_2 _10356_ (.CLK(clknet_leaf_131_wb_clk_i),
    .D(_00161_),
    .Q(\tms1x00.ins_pla_ors[8][12] ));
 sky130_fd_sc_hd__dfxtp_1 _10357_ (.CLK(clknet_leaf_131_wb_clk_i),
    .D(_00162_),
    .Q(\tms1x00.ins_pla_ors[8][13] ));
 sky130_fd_sc_hd__dfxtp_1 _10358_ (.CLK(clknet_leaf_116_wb_clk_i),
    .D(_00163_),
    .Q(\tms1x00.ins_pla_ors[8][15] ));
 sky130_fd_sc_hd__dfxtp_1 _10359_ (.CLK(clknet_leaf_133_wb_clk_i),
    .D(_00164_),
    .Q(\tms1x00.ins_pla_ors[8][19] ));
 sky130_fd_sc_hd__dfxtp_2 _10360_ (.CLK(clknet_leaf_117_wb_clk_i),
    .D(_00165_),
    .Q(\tms1x00.ins_pla_ors[8][22] ));
 sky130_fd_sc_hd__dfxtp_1 _10361_ (.CLK(clknet_leaf_120_wb_clk_i),
    .D(_00166_),
    .Q(\tms1x00.ins_pla_ors[8][27] ));
 sky130_fd_sc_hd__dfxtp_1 _10362_ (.CLK(clknet_leaf_117_wb_clk_i),
    .D(_00167_),
    .Q(\tms1x00.ins_pla_ors[8][28] ));
 sky130_fd_sc_hd__dfxtp_2 _10363_ (.CLK(clknet_leaf_120_wb_clk_i),
    .D(_00168_),
    .Q(\tms1x00.ins_pla_ors[8][29] ));
 sky130_fd_sc_hd__dfxtp_1 _10364_ (.CLK(clknet_leaf_124_wb_clk_i),
    .D(_00169_),
    .Q(\tms1x00.ins_pla_ors[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10365_ (.CLK(clknet_leaf_127_wb_clk_i),
    .D(_00170_),
    .Q(\tms1x00.ins_pla_ors[13][8] ));
 sky130_fd_sc_hd__dfxtp_1 _10366_ (.CLK(clknet_leaf_124_wb_clk_i),
    .D(_00171_),
    .Q(\tms1x00.ins_pla_ors[13][9] ));
 sky130_fd_sc_hd__dfxtp_1 _10367_ (.CLK(clknet_leaf_128_wb_clk_i),
    .D(_00172_),
    .Q(\tms1x00.ins_pla_ors[13][11] ));
 sky130_fd_sc_hd__dfxtp_1 _10368_ (.CLK(clknet_leaf_131_wb_clk_i),
    .D(_00173_),
    .Q(\tms1x00.ins_pla_ors[13][14] ));
 sky130_fd_sc_hd__dfxtp_1 _10369_ (.CLK(clknet_leaf_123_wb_clk_i),
    .D(_00174_),
    .Q(\tms1x00.ins_pla_ors[13][15] ));
 sky130_fd_sc_hd__dfxtp_1 _10370_ (.CLK(clknet_leaf_122_wb_clk_i),
    .D(_00175_),
    .Q(\tms1x00.ins_pla_ors[13][16] ));
 sky130_fd_sc_hd__dfxtp_1 _10371_ (.CLK(clknet_leaf_123_wb_clk_i),
    .D(_00176_),
    .Q(\tms1x00.ins_pla_ors[13][18] ));
 sky130_fd_sc_hd__dfxtp_1 _10372_ (.CLK(clknet_leaf_120_wb_clk_i),
    .D(_00177_),
    .Q(\tms1x00.ins_pla_ors[13][20] ));
 sky130_fd_sc_hd__dfxtp_1 _10373_ (.CLK(clknet_leaf_134_wb_clk_i),
    .D(_00178_),
    .Q(\tms1x00.ins_pla_ors[13][21] ));
 sky130_fd_sc_hd__dfxtp_1 _10374_ (.CLK(clknet_leaf_123_wb_clk_i),
    .D(_00179_),
    .Q(\tms1x00.ins_pla_ors[13][25] ));
 sky130_fd_sc_hd__dfxtp_1 _10375_ (.CLK(clknet_leaf_117_wb_clk_i),
    .D(_00180_),
    .Q(\tms1x00.ins_pla_ors[13][26] ));
 sky130_fd_sc_hd__dfxtp_1 _10376_ (.CLK(clknet_leaf_119_wb_clk_i),
    .D(_00181_),
    .Q(\tms1x00.ins_pla_ors[13][27] ));
 sky130_fd_sc_hd__dfxtp_1 _10377_ (.CLK(clknet_leaf_113_wb_clk_i),
    .D(_00182_),
    .Q(\tms1x00.ins_pla_ors[13][28] ));
 sky130_fd_sc_hd__dfxtp_1 _10378_ (.CLK(clknet_leaf_120_wb_clk_i),
    .D(_00183_),
    .Q(\tms1x00.ins_pla_ors[13][29] ));
 sky130_fd_sc_hd__dfxtp_1 _10379_ (.CLK(clknet_leaf_129_wb_clk_i),
    .D(_00184_),
    .Q(\tms1x00.ins_pla_ors[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10380_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_00185_),
    .Q(\tms1x00.ins_pla_ors[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _10381_ (.CLK(clknet_leaf_123_wb_clk_i),
    .D(_00186_),
    .Q(\tms1x00.ins_pla_ors[11][3] ));
 sky130_fd_sc_hd__dfxtp_2 _10382_ (.CLK(clknet_leaf_126_wb_clk_i),
    .D(_00187_),
    .Q(\tms1x00.ins_pla_ors[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 _10383_ (.CLK(clknet_leaf_90_wb_clk_i),
    .D(_00188_),
    .Q(\tms1x00.ins_pla_ors[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 _10384_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_00189_),
    .Q(\tms1x00.ins_pla_ors[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 _10385_ (.CLK(clknet_leaf_136_wb_clk_i),
    .D(_00190_),
    .Q(\tms1x00.ins_pla_ors[11][13] ));
 sky130_fd_sc_hd__dfxtp_1 _10386_ (.CLK(clknet_leaf_136_wb_clk_i),
    .D(_00191_),
    .Q(\tms1x00.ins_pla_ors[11][14] ));
 sky130_fd_sc_hd__dfxtp_1 _10387_ (.CLK(clknet_leaf_132_wb_clk_i),
    .D(_00192_),
    .Q(\tms1x00.ins_pla_ors[11][15] ));
 sky130_fd_sc_hd__dfxtp_1 _10388_ (.CLK(clknet_leaf_122_wb_clk_i),
    .D(_00193_),
    .Q(\tms1x00.ins_pla_ors[11][16] ));
 sky130_fd_sc_hd__dfxtp_1 _10389_ (.CLK(clknet_leaf_121_wb_clk_i),
    .D(_00194_),
    .Q(\tms1x00.ins_pla_ors[11][17] ));
 sky130_fd_sc_hd__dfxtp_1 _10390_ (.CLK(clknet_leaf_121_wb_clk_i),
    .D(_00195_),
    .Q(\tms1x00.ins_pla_ors[11][18] ));
 sky130_fd_sc_hd__dfxtp_1 _10391_ (.CLK(clknet_leaf_132_wb_clk_i),
    .D(_00196_),
    .Q(\tms1x00.ins_pla_ors[11][19] ));
 sky130_fd_sc_hd__dfxtp_2 _10392_ (.CLK(clknet_leaf_134_wb_clk_i),
    .D(_00197_),
    .Q(\tms1x00.ins_pla_ors[11][21] ));
 sky130_fd_sc_hd__dfxtp_1 _10393_ (.CLK(clknet_leaf_116_wb_clk_i),
    .D(_00198_),
    .Q(\tms1x00.ins_pla_ors[11][22] ));
 sky130_fd_sc_hd__dfxtp_1 _10394_ (.CLK(clknet_leaf_118_wb_clk_i),
    .D(_00199_),
    .Q(\tms1x00.ins_pla_ors[11][25] ));
 sky130_fd_sc_hd__dfxtp_1 _10395_ (.CLK(clknet_leaf_116_wb_clk_i),
    .D(_00200_),
    .Q(\tms1x00.ins_pla_ors[11][26] ));
 sky130_fd_sc_hd__dfxtp_1 _10396_ (.CLK(clknet_leaf_99_wb_clk_i),
    .D(_00201_),
    .Q(\tms1x00.ins_pla_ors[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10397_ (.CLK(clknet_leaf_95_wb_clk_i),
    .D(_00202_),
    .Q(\tms1x00.ins_pla_ors[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _10398_ (.CLK(clknet_leaf_97_wb_clk_i),
    .D(_00203_),
    .Q(\tms1x00.ins_pla_ors[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _10399_ (.CLK(clknet_leaf_101_wb_clk_i),
    .D(_00204_),
    .Q(\tms1x00.ins_pla_ors[3][5] ));
 sky130_fd_sc_hd__dfxtp_2 _10400_ (.CLK(clknet_leaf_102_wb_clk_i),
    .D(_00205_),
    .Q(\tms1x00.ins_pla_ors[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _10401_ (.CLK(clknet_leaf_91_wb_clk_i),
    .D(_00206_),
    .Q(\tms1x00.ins_pla_ors[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _10402_ (.CLK(clknet_leaf_100_wb_clk_i),
    .D(_00207_),
    .Q(\tms1x00.ins_pla_ors[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _10403_ (.CLK(clknet_leaf_100_wb_clk_i),
    .D(_00208_),
    .Q(\tms1x00.ins_pla_ors[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _10404_ (.CLK(clknet_leaf_91_wb_clk_i),
    .D(_00209_),
    .Q(\tms1x00.ins_pla_ors[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _10405_ (.CLK(clknet_leaf_98_wb_clk_i),
    .D(_00210_),
    .Q(\tms1x00.ins_pla_ors[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _10406_ (.CLK(clknet_leaf_110_wb_clk_i),
    .D(_00211_),
    .Q(\tms1x00.ins_pla_ors[3][15] ));
 sky130_fd_sc_hd__dfxtp_2 _10407_ (.CLK(clknet_leaf_100_wb_clk_i),
    .D(_00212_),
    .Q(\tms1x00.ins_pla_ors[3][16] ));
 sky130_fd_sc_hd__dfxtp_1 _10408_ (.CLK(clknet_leaf_103_wb_clk_i),
    .D(_00213_),
    .Q(\tms1x00.ins_pla_ors[3][17] ));
 sky130_fd_sc_hd__dfxtp_2 _10409_ (.CLK(clknet_leaf_107_wb_clk_i),
    .D(_00214_),
    .Q(\tms1x00.ins_pla_ors[3][18] ));
 sky130_fd_sc_hd__dfxtp_2 _10410_ (.CLK(clknet_leaf_102_wb_clk_i),
    .D(_00215_),
    .Q(\tms1x00.ins_pla_ors[3][19] ));
 sky130_fd_sc_hd__dfxtp_2 _10411_ (.CLK(clknet_leaf_107_wb_clk_i),
    .D(_00216_),
    .Q(\tms1x00.ins_pla_ors[3][20] ));
 sky130_fd_sc_hd__dfxtp_1 _10412_ (.CLK(clknet_leaf_111_wb_clk_i),
    .D(_00217_),
    .Q(\tms1x00.ins_pla_ors[3][22] ));
 sky130_fd_sc_hd__dfxtp_2 _10413_ (.CLK(clknet_leaf_102_wb_clk_i),
    .D(_00218_),
    .Q(\tms1x00.ins_pla_ors[3][23] ));
 sky130_fd_sc_hd__dfxtp_1 _10414_ (.CLK(clknet_leaf_108_wb_clk_i),
    .D(_00219_),
    .Q(\tms1x00.ins_pla_ors[3][26] ));
 sky130_fd_sc_hd__dfxtp_1 _10415_ (.CLK(clknet_leaf_106_wb_clk_i),
    .D(_00220_),
    .Q(\tms1x00.ins_pla_ors[3][27] ));
 sky130_fd_sc_hd__dfxtp_1 _10416_ (.CLK(clknet_leaf_111_wb_clk_i),
    .D(_00221_),
    .Q(\tms1x00.ins_pla_ors[3][28] ));
 sky130_fd_sc_hd__dfxtp_1 _10417_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_00222_),
    .Q(\tms1x00.ins_pla_ands[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10418_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_00223_),
    .Q(\tms1x00.ins_pla_ands[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _10419_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_00224_),
    .Q(\tms1x00.ins_pla_ands[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _10420_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_00225_),
    .Q(\tms1x00.ins_pla_ands[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _10421_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_00226_),
    .Q(\tms1x00.ins_pla_ands[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _10422_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_00227_),
    .Q(\tms1x00.ins_pla_ands[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _10423_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_00228_),
    .Q(\tms1x00.ins_pla_ands[6][8] ));
 sky130_fd_sc_hd__dfxtp_1 _10424_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_00229_),
    .Q(\tms1x00.ins_pla_ands[6][9] ));
 sky130_fd_sc_hd__dfxtp_1 _10425_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_00230_),
    .Q(\tms1x00.ins_pla_ands[6][10] ));
 sky130_fd_sc_hd__dfxtp_1 _10426_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_00231_),
    .Q(\tms1x00.ins_pla_ands[6][11] ));
 sky130_fd_sc_hd__dfxtp_1 _10427_ (.CLK(clknet_leaf_58_wb_clk_i),
    .D(_00232_),
    .Q(\tms1x00.ins_pla_ands[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10428_ (.CLK(clknet_leaf_56_wb_clk_i),
    .D(_00233_),
    .Q(\tms1x00.ins_pla_ands[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _10429_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(_00234_),
    .Q(\tms1x00.ins_pla_ands[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _10430_ (.CLK(clknet_leaf_56_wb_clk_i),
    .D(_00235_),
    .Q(\tms1x00.ins_pla_ands[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _10431_ (.CLK(clknet_leaf_58_wb_clk_i),
    .D(_00236_),
    .Q(\tms1x00.ins_pla_ands[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _10432_ (.CLK(clknet_leaf_58_wb_clk_i),
    .D(_00237_),
    .Q(\tms1x00.ins_pla_ands[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _10433_ (.CLK(clknet_leaf_58_wb_clk_i),
    .D(_00238_),
    .Q(\tms1x00.ins_pla_ands[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _10434_ (.CLK(clknet_leaf_58_wb_clk_i),
    .D(_00239_),
    .Q(\tms1x00.ins_pla_ands[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _10435_ (.CLK(clknet_leaf_130_wb_clk_i),
    .D(_00240_),
    .Q(\tms1x00.ins_pla_ands[29][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10436_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_00241_),
    .Q(\tms1x00.ins_pla_ands[29][1] ));
 sky130_fd_sc_hd__dfxtp_1 _10437_ (.CLK(clknet_leaf_139_wb_clk_i),
    .D(_00242_),
    .Q(\tms1x00.ins_pla_ands[29][2] ));
 sky130_fd_sc_hd__dfxtp_1 _10438_ (.CLK(clknet_leaf_141_wb_clk_i),
    .D(_00243_),
    .Q(\tms1x00.ins_pla_ands[29][3] ));
 sky130_fd_sc_hd__dfxtp_1 _10439_ (.CLK(clknet_leaf_140_wb_clk_i),
    .D(_00244_),
    .Q(\tms1x00.ins_pla_ands[29][4] ));
 sky130_fd_sc_hd__dfxtp_1 _10440_ (.CLK(clknet_leaf_140_wb_clk_i),
    .D(_00245_),
    .Q(\tms1x00.ins_pla_ands[29][5] ));
 sky130_fd_sc_hd__dfxtp_1 _10441_ (.CLK(clknet_leaf_141_wb_clk_i),
    .D(_00246_),
    .Q(\tms1x00.ins_pla_ands[29][6] ));
 sky130_fd_sc_hd__dfxtp_1 _10442_ (.CLK(clknet_leaf_141_wb_clk_i),
    .D(_00247_),
    .Q(\tms1x00.ins_pla_ands[29][7] ));
 sky130_fd_sc_hd__dfxtp_1 _10443_ (.CLK(clknet_leaf_139_wb_clk_i),
    .D(_00248_),
    .Q(\tms1x00.ins_pla_ands[29][9] ));
 sky130_fd_sc_hd__dfxtp_1 _10444_ (.CLK(clknet_leaf_130_wb_clk_i),
    .D(_00249_),
    .Q(\tms1x00.ins_pla_ands[29][11] ));
 sky130_fd_sc_hd__dfxtp_1 _10445_ (.CLK(clknet_leaf_138_wb_clk_i),
    .D(_00250_),
    .Q(\tms1x00.ins_pla_ands[29][12] ));
 sky130_fd_sc_hd__dfxtp_1 _10446_ (.CLK(clknet_leaf_138_wb_clk_i),
    .D(_00251_),
    .Q(\tms1x00.ins_pla_ands[29][15] ));
 sky130_fd_sc_hd__dfxtp_1 _10447_ (.CLK(clknet_leaf_139_wb_clk_i),
    .D(_00252_),
    .Q(\tms1x00.ins_pla_ands[27][8] ));
 sky130_fd_sc_hd__dfxtp_1 _10448_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_00253_),
    .Q(\tms1x00.ins_pla_ands[27][11] ));
 sky130_fd_sc_hd__dfxtp_1 _10449_ (.CLK(clknet_leaf_136_wb_clk_i),
    .D(_00254_),
    .Q(\tms1x00.ins_pla_ands[27][13] ));
 sky130_fd_sc_hd__dfxtp_1 _10450_ (.CLK(clknet_leaf_138_wb_clk_i),
    .D(_00255_),
    .Q(\tms1x00.ins_pla_ands[27][14] ));
 sky130_fd_sc_hd__dfxtp_1 _10451_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_00256_),
    .Q(\tms1x00.ins_pla_ands[23][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10452_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_00257_),
    .Q(\tms1x00.ins_pla_ands[23][1] ));
 sky130_fd_sc_hd__dfxtp_1 _10453_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_00258_),
    .Q(\tms1x00.ins_pla_ands[23][10] ));
 sky130_fd_sc_hd__dfxtp_1 _10454_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_00259_),
    .Q(\tms1x00.ins_pla_ands[23][11] ));
 sky130_fd_sc_hd__dfxtp_1 _10455_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_00260_),
    .Q(\tms1x00.ins_pla_ands[22][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10456_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_00261_),
    .Q(\tms1x00.ins_pla_ands[22][1] ));
 sky130_fd_sc_hd__dfxtp_1 _10457_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_00262_),
    .Q(\tms1x00.ins_pla_ands[22][2] ));
 sky130_fd_sc_hd__dfxtp_1 _10458_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_00263_),
    .Q(\tms1x00.ins_pla_ands[22][3] ));
 sky130_fd_sc_hd__dfxtp_1 _10459_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_00264_),
    .Q(\tms1x00.ins_pla_ands[22][4] ));
 sky130_fd_sc_hd__dfxtp_1 _10460_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_00265_),
    .Q(\tms1x00.ins_pla_ands[22][5] ));
 sky130_fd_sc_hd__dfxtp_1 _10461_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_00266_),
    .Q(\tms1x00.ins_pla_ands[22][11] ));
 sky130_fd_sc_hd__dfxtp_1 _10462_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_00267_),
    .Q(\tms1x00.ins_pla_ands[19][2] ));
 sky130_fd_sc_hd__dfxtp_1 _10463_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_00268_),
    .Q(\tms1x00.ins_pla_ands[19][3] ));
 sky130_fd_sc_hd__dfxtp_1 _10464_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_00269_),
    .Q(\tms1x00.ins_pla_ands[19][4] ));
 sky130_fd_sc_hd__dfxtp_1 _10465_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_00270_),
    .Q(\tms1x00.ins_pla_ands[19][5] ));
 sky130_fd_sc_hd__dfxtp_1 _10466_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_00271_),
    .Q(\tms1x00.ins_pla_ands[19][6] ));
 sky130_fd_sc_hd__dfxtp_1 _10467_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_00272_),
    .Q(\tms1x00.ins_pla_ands[19][7] ));
 sky130_fd_sc_hd__dfxtp_1 _10468_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_00273_),
    .Q(\tms1x00.ins_pla_ands[19][8] ));
 sky130_fd_sc_hd__dfxtp_1 _10469_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_00274_),
    .Q(\tms1x00.ins_pla_ands[19][9] ));
 sky130_fd_sc_hd__dfxtp_1 _10470_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_00275_),
    .Q(\tms1x00.ins_pla_ands[19][12] ));
 sky130_fd_sc_hd__dfxtp_1 _10471_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_00276_),
    .Q(\tms1x00.ins_pla_ands[19][13] ));
 sky130_fd_sc_hd__dfxtp_1 _10472_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_00277_),
    .Q(\tms1x00.ins_pla_ands[19][14] ));
 sky130_fd_sc_hd__dfxtp_1 _10473_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_00278_),
    .Q(\tms1x00.ins_pla_ands[19][15] ));
 sky130_fd_sc_hd__dfxtp_1 _10474_ (.CLK(clknet_leaf_134_wb_clk_i),
    .D(_00279_),
    .Q(\tms1x00.ins_pla_ors[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10475_ (.CLK(clknet_leaf_128_wb_clk_i),
    .D(_00280_),
    .Q(\tms1x00.ins_pla_ors[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _10476_ (.CLK(clknet_leaf_90_wb_clk_i),
    .D(_00281_),
    .Q(\tms1x00.ins_pla_ors[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _10477_ (.CLK(clknet_leaf_134_wb_clk_i),
    .D(_00282_),
    .Q(\tms1x00.ins_pla_ors[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _10478_ (.CLK(clknet_leaf_125_wb_clk_i),
    .D(_00283_),
    .Q(\tms1x00.ins_pla_ors[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _10479_ (.CLK(clknet_leaf_126_wb_clk_i),
    .D(_00284_),
    .Q(\tms1x00.ins_pla_ors[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _10480_ (.CLK(clknet_leaf_115_wb_clk_i),
    .D(_00285_),
    .Q(\tms1x00.ins_pla_ors[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 _10481_ (.CLK(clknet_leaf_126_wb_clk_i),
    .D(_00286_),
    .Q(\tms1x00.ins_pla_ors[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 _10482_ (.CLK(clknet_leaf_90_wb_clk_i),
    .D(_00287_),
    .Q(\tms1x00.ins_pla_ors[8][8] ));
 sky130_fd_sc_hd__dfxtp_1 _10483_ (.CLK(clknet_leaf_133_wb_clk_i),
    .D(_00288_),
    .Q(\tms1x00.ins_pla_ors[8][9] ));
 sky130_fd_sc_hd__dfxtp_1 _10484_ (.CLK(clknet_leaf_132_wb_clk_i),
    .D(_00289_),
    .Q(\tms1x00.ins_pla_ors[8][10] ));
 sky130_fd_sc_hd__dfxtp_1 _10485_ (.CLK(clknet_leaf_128_wb_clk_i),
    .D(_00290_),
    .Q(\tms1x00.ins_pla_ors[8][11] ));
 sky130_fd_sc_hd__dfxtp_1 _10486_ (.CLK(clknet_leaf_133_wb_clk_i),
    .D(_00291_),
    .Q(\tms1x00.ins_pla_ors[8][14] ));
 sky130_fd_sc_hd__dfxtp_2 _10487_ (.CLK(clknet_leaf_114_wb_clk_i),
    .D(_00292_),
    .Q(\tms1x00.ins_pla_ors[8][16] ));
 sky130_fd_sc_hd__dfxtp_2 _10488_ (.CLK(clknet_leaf_114_wb_clk_i),
    .D(_00293_),
    .Q(\tms1x00.ins_pla_ors[8][17] ));
 sky130_fd_sc_hd__dfxtp_1 _10489_ (.CLK(clknet_leaf_122_wb_clk_i),
    .D(_00294_),
    .Q(\tms1x00.ins_pla_ors[8][18] ));
 sky130_fd_sc_hd__dfxtp_1 _10490_ (.CLK(clknet_leaf_114_wb_clk_i),
    .D(_00295_),
    .Q(\tms1x00.ins_pla_ors[8][20] ));
 sky130_fd_sc_hd__dfxtp_1 _10491_ (.CLK(clknet_leaf_134_wb_clk_i),
    .D(_00296_),
    .Q(\tms1x00.ins_pla_ors[8][21] ));
 sky130_fd_sc_hd__dfxtp_2 _10492_ (.CLK(clknet_leaf_115_wb_clk_i),
    .D(_00297_),
    .Q(\tms1x00.ins_pla_ors[8][23] ));
 sky130_fd_sc_hd__dfxtp_2 _10493_ (.CLK(clknet_leaf_115_wb_clk_i),
    .D(_00298_),
    .Q(\tms1x00.ins_pla_ors[8][24] ));
 sky130_fd_sc_hd__dfxtp_1 _10494_ (.CLK(clknet_leaf_116_wb_clk_i),
    .D(_00299_),
    .Q(\tms1x00.ins_pla_ors[8][25] ));
 sky130_fd_sc_hd__dfxtp_1 _10495_ (.CLK(clknet_leaf_116_wb_clk_i),
    .D(_00300_),
    .Q(\tms1x00.ins_pla_ors[8][26] ));
 sky130_fd_sc_hd__dfxtp_2 _10496_ (.CLK(clknet_leaf_105_wb_clk_i),
    .D(_00301_),
    .Q(\tms1x00.ins_pla_ors[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10497_ (.CLK(clknet_leaf_95_wb_clk_i),
    .D(_00302_),
    .Q(\tms1x00.ins_pla_ors[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _10498_ (.CLK(clknet_leaf_95_wb_clk_i),
    .D(_00303_),
    .Q(\tms1x00.ins_pla_ors[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _10499_ (.CLK(clknet_leaf_95_wb_clk_i),
    .D(_00304_),
    .Q(\tms1x00.ins_pla_ors[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _10500_ (.CLK(clknet_leaf_103_wb_clk_i),
    .D(_00305_),
    .Q(\tms1x00.ins_pla_ors[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _10501_ (.CLK(clknet_leaf_103_wb_clk_i),
    .D(_00306_),
    .Q(\tms1x00.ins_pla_ors[2][18] ));
 sky130_fd_sc_hd__dfxtp_2 _10502_ (.CLK(clknet_leaf_111_wb_clk_i),
    .D(_00307_),
    .Q(\tms1x00.ins_pla_ors[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _10503_ (.CLK(clknet_leaf_105_wb_clk_i),
    .D(_00308_),
    .Q(\tms1x00.ins_pla_ors[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _10504_ (.CLK(clknet_leaf_105_wb_clk_i),
    .D(_00309_),
    .Q(\tms1x00.ins_pla_ors[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _10505_ (.CLK(clknet_leaf_95_wb_clk_i),
    .D(_00310_),
    .Q(\tms1x00.ins_pla_ors[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _10506_ (.CLK(clknet_leaf_112_wb_clk_i),
    .D(_00311_),
    .Q(\tms1x00.ins_pla_ors[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _10507_ (.CLK(clknet_leaf_132_wb_clk_i),
    .D(_00312_),
    .Q(\tms1x00.ins_pla_ors[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10508_ (.CLK(clknet_leaf_89_wb_clk_i),
    .D(_00313_),
    .Q(\tms1x00.ins_pla_ors[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 _10509_ (.CLK(clknet_leaf_126_wb_clk_i),
    .D(_00314_),
    .Q(\tms1x00.ins_pla_ors[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 _10510_ (.CLK(clknet_leaf_126_wb_clk_i),
    .D(_00315_),
    .Q(\tms1x00.ins_pla_ors[12][9] ));
 sky130_fd_sc_hd__dfxtp_1 _10511_ (.CLK(clknet_leaf_124_wb_clk_i),
    .D(_00316_),
    .Q(\tms1x00.ins_pla_ors[12][10] ));
 sky130_fd_sc_hd__dfxtp_1 _10512_ (.CLK(clknet_leaf_124_wb_clk_i),
    .D(_00317_),
    .Q(\tms1x00.ins_pla_ors[12][11] ));
 sky130_fd_sc_hd__dfxtp_1 _10513_ (.CLK(clknet_leaf_132_wb_clk_i),
    .D(_00318_),
    .Q(\tms1x00.ins_pla_ors[12][12] ));
 sky130_fd_sc_hd__dfxtp_1 _10514_ (.CLK(clknet_leaf_128_wb_clk_i),
    .D(_00319_),
    .Q(\tms1x00.ins_pla_ors[12][13] ));
 sky130_fd_sc_hd__dfxtp_1 _10515_ (.CLK(clknet_leaf_118_wb_clk_i),
    .D(_00320_),
    .Q(\tms1x00.ins_pla_ors[12][15] ));
 sky130_fd_sc_hd__dfxtp_1 _10516_ (.CLK(clknet_leaf_128_wb_clk_i),
    .D(_00321_),
    .Q(\tms1x00.ins_pla_ors[12][19] ));
 sky130_fd_sc_hd__dfxtp_2 _10517_ (.CLK(clknet_leaf_113_wb_clk_i),
    .D(_00322_),
    .Q(\tms1x00.ins_pla_ors[12][20] ));
 sky130_fd_sc_hd__dfxtp_1 _10518_ (.CLK(clknet_leaf_113_wb_clk_i),
    .D(_00323_),
    .Q(\tms1x00.ins_pla_ors[12][22] ));
 sky130_fd_sc_hd__dfxtp_2 _10519_ (.CLK(clknet_leaf_113_wb_clk_i),
    .D(_00324_),
    .Q(\tms1x00.ins_pla_ors[12][23] ));
 sky130_fd_sc_hd__dfxtp_1 _10520_ (.CLK(clknet_leaf_122_wb_clk_i),
    .D(_00325_),
    .Q(\tms1x00.ins_pla_ors[12][24] ));
 sky130_fd_sc_hd__dfxtp_1 _10521_ (.CLK(clknet_leaf_123_wb_clk_i),
    .D(_00326_),
    .Q(\tms1x00.ins_pla_ors[12][25] ));
 sky130_fd_sc_hd__dfxtp_1 _10522_ (.CLK(clknet_leaf_118_wb_clk_i),
    .D(_00327_),
    .Q(\tms1x00.ins_pla_ors[12][27] ));
 sky130_fd_sc_hd__dfxtp_2 _10523_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_00328_),
    .Q(\tms1x00.ins_pla_ors[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _10524_ (.CLK(clknet_leaf_129_wb_clk_i),
    .D(_00329_),
    .Q(\tms1x00.ins_pla_ors[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 _10525_ (.CLK(clknet_leaf_128_wb_clk_i),
    .D(_00330_),
    .Q(\tms1x00.ins_pla_ors[14][12] ));
 sky130_fd_sc_hd__dfxtp_2 _10526_ (.CLK(clknet_leaf_134_wb_clk_i),
    .D(_00331_),
    .Q(\tms1x00.ins_pla_ors[14][13] ));
 sky130_fd_sc_hd__dfxtp_2 _10527_ (.CLK(clknet_leaf_122_wb_clk_i),
    .D(_00332_),
    .Q(\tms1x00.ins_pla_ors[14][16] ));
 sky130_fd_sc_hd__dfxtp_1 _10528_ (.CLK(clknet_leaf_116_wb_clk_i),
    .D(_00333_),
    .Q(\tms1x00.ins_pla_ors[14][22] ));
 sky130_fd_sc_hd__dfxtp_1 _10529_ (.CLK(clknet_leaf_117_wb_clk_i),
    .D(_00334_),
    .Q(\tms1x00.ins_pla_ors[14][23] ));
 sky130_fd_sc_hd__dfxtp_1 _10530_ (.CLK(clknet_leaf_118_wb_clk_i),
    .D(_00335_),
    .Q(\tms1x00.ins_pla_ors[14][25] ));
 sky130_fd_sc_hd__dfxtp_1 _10531_ (.CLK(clknet_leaf_120_wb_clk_i),
    .D(_00336_),
    .Q(\tms1x00.ins_pla_ors[14][27] ));
 sky130_fd_sc_hd__dfxtp_1 _10532_ (.CLK(clknet_leaf_120_wb_clk_i),
    .D(_00337_),
    .Q(\tms1x00.ins_pla_ors[14][29] ));
 sky130_fd_sc_hd__dfxtp_1 _10533_ (.CLK(clknet_leaf_97_wb_clk_i),
    .D(_00338_),
    .Q(\tms1x00.ins_pla_ors[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _10534_ (.CLK(clknet_leaf_97_wb_clk_i),
    .D(_00339_),
    .Q(\tms1x00.ins_pla_ors[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _10535_ (.CLK(clknet_leaf_97_wb_clk_i),
    .D(_00340_),
    .Q(\tms1x00.ins_pla_ors[2][5] ));
 sky130_fd_sc_hd__dfxtp_2 _10536_ (.CLK(clknet_leaf_100_wb_clk_i),
    .D(_00341_),
    .Q(\tms1x00.ins_pla_ors[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _10537_ (.CLK(clknet_leaf_96_wb_clk_i),
    .D(_00342_),
    .Q(\tms1x00.ins_pla_ors[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _10538_ (.CLK(clknet_leaf_98_wb_clk_i),
    .D(_00343_),
    .Q(\tms1x00.ins_pla_ors[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _10539_ (.CLK(clknet_leaf_95_wb_clk_i),
    .D(_00344_),
    .Q(\tms1x00.ins_pla_ors[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _10540_ (.CLK(clknet_leaf_104_wb_clk_i),
    .D(_00345_),
    .Q(\tms1x00.ins_pla_ors[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _10541_ (.CLK(clknet_leaf_104_wb_clk_i),
    .D(_00346_),
    .Q(\tms1x00.ins_pla_ors[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _10542_ (.CLK(clknet_leaf_98_wb_clk_i),
    .D(_00347_),
    .Q(\tms1x00.ins_pla_ors[2][13] ));
 sky130_fd_sc_hd__dfxtp_2 _10543_ (.CLK(clknet_leaf_107_wb_clk_i),
    .D(_00348_),
    .Q(\tms1x00.ins_pla_ors[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _10544_ (.CLK(clknet_leaf_109_wb_clk_i),
    .D(_00349_),
    .Q(\tms1x00.ins_pla_ors[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _10545_ (.CLK(clknet_leaf_102_wb_clk_i),
    .D(_00350_),
    .Q(\tms1x00.ins_pla_ors[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _10546_ (.CLK(clknet_leaf_106_wb_clk_i),
    .D(_00351_),
    .Q(\tms1x00.ins_pla_ors[2][19] ));
 sky130_fd_sc_hd__dfxtp_2 _10547_ (.CLK(clknet_leaf_107_wb_clk_i),
    .D(_00352_),
    .Q(\tms1x00.ins_pla_ors[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _10548_ (.CLK(clknet_leaf_109_wb_clk_i),
    .D(_00353_),
    .Q(\tms1x00.ins_pla_ors[2][21] ));
 sky130_fd_sc_hd__dfxtp_2 _10549_ (.CLK(clknet_leaf_110_wb_clk_i),
    .D(_00354_),
    .Q(\tms1x00.ins_pla_ors[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _10550_ (.CLK(clknet_leaf_102_wb_clk_i),
    .D(_00355_),
    .Q(\tms1x00.ins_pla_ors[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _10551_ (.CLK(clknet_leaf_101_wb_clk_i),
    .D(_00356_),
    .Q(\tms1x00.ins_pla_ors[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _10552_ (.CLK(clknet_leaf_110_wb_clk_i),
    .D(_00357_),
    .Q(\tms1x00.ins_pla_ors[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _10553_ (.CLK(clknet_leaf_104_wb_clk_i),
    .D(_00358_),
    .Q(\tms1x00.ins_pla_ors[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _10554_ (.CLK(clknet_leaf_81_wb_clk_i),
    .D(_00359_),
    .Q(\tms1x00.ins_pla_ors[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10555_ (.CLK(clknet_leaf_83_wb_clk_i),
    .D(_00360_),
    .Q(\tms1x00.ins_pla_ors[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _10556_ (.CLK(clknet_leaf_83_wb_clk_i),
    .D(_00361_),
    .Q(\tms1x00.ins_pla_ors[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _10557_ (.CLK(clknet_leaf_92_wb_clk_i),
    .D(_00362_),
    .Q(\tms1x00.ins_pla_ors[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _10558_ (.CLK(clknet_leaf_82_wb_clk_i),
    .D(_00363_),
    .Q(\tms1x00.ins_pla_ors[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _10559_ (.CLK(clknet_leaf_97_wb_clk_i),
    .D(_00364_),
    .Q(\tms1x00.ins_pla_ors[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _10560_ (.CLK(clknet_leaf_102_wb_clk_i),
    .D(_00365_),
    .Q(\tms1x00.ins_pla_ors[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _10561_ (.CLK(clknet_leaf_83_wb_clk_i),
    .D(_00366_),
    .Q(\tms1x00.ins_pla_ors[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _10562_ (.CLK(clknet_leaf_83_wb_clk_i),
    .D(_00367_),
    .Q(\tms1x00.ins_pla_ors[7][8] ));
 sky130_fd_sc_hd__dfxtp_1 _10563_ (.CLK(clknet_leaf_81_wb_clk_i),
    .D(_00368_),
    .Q(\tms1x00.ins_pla_ors[7][9] ));
 sky130_fd_sc_hd__dfxtp_1 _10564_ (.CLK(clknet_leaf_81_wb_clk_i),
    .D(_00369_),
    .Q(\tms1x00.ins_pla_ors[7][10] ));
 sky130_fd_sc_hd__dfxtp_1 _10565_ (.CLK(clknet_leaf_104_wb_clk_i),
    .D(_00370_),
    .Q(\tms1x00.ins_pla_ors[7][11] ));
 sky130_fd_sc_hd__dfxtp_1 _10566_ (.CLK(clknet_leaf_104_wb_clk_i),
    .D(_00371_),
    .Q(\tms1x00.ins_pla_ors[7][12] ));
 sky130_fd_sc_hd__dfxtp_1 _10567_ (.CLK(clknet_leaf_82_wb_clk_i),
    .D(_00372_),
    .Q(\tms1x00.ins_pla_ors[7][13] ));
 sky130_fd_sc_hd__dfxtp_1 _10568_ (.CLK(clknet_leaf_112_wb_clk_i),
    .D(_00373_),
    .Q(\tms1x00.ins_pla_ors[7][14] ));
 sky130_fd_sc_hd__dfxtp_2 _10569_ (.CLK(clknet_leaf_110_wb_clk_i),
    .D(_00374_),
    .Q(\tms1x00.ins_pla_ors[7][15] ));
 sky130_fd_sc_hd__dfxtp_1 _10570_ (.CLK(clknet_leaf_102_wb_clk_i),
    .D(_00375_),
    .Q(\tms1x00.ins_pla_ors[7][16] ));
 sky130_fd_sc_hd__dfxtp_1 _10571_ (.CLK(clknet_leaf_107_wb_clk_i),
    .D(_00376_),
    .Q(\tms1x00.ins_pla_ors[7][17] ));
 sky130_fd_sc_hd__dfxtp_1 _10572_ (.CLK(clknet_leaf_102_wb_clk_i),
    .D(_00377_),
    .Q(\tms1x00.ins_pla_ors[7][18] ));
 sky130_fd_sc_hd__dfxtp_2 _10573_ (.CLK(clknet_leaf_107_wb_clk_i),
    .D(_00378_),
    .Q(\tms1x00.ins_pla_ors[7][19] ));
 sky130_fd_sc_hd__dfxtp_1 _10574_ (.CLK(clknet_leaf_107_wb_clk_i),
    .D(_00379_),
    .Q(\tms1x00.ins_pla_ors[7][20] ));
 sky130_fd_sc_hd__dfxtp_1 _10575_ (.CLK(clknet_leaf_108_wb_clk_i),
    .D(_00380_),
    .Q(\tms1x00.ins_pla_ors[7][21] ));
 sky130_fd_sc_hd__dfxtp_2 _10576_ (.CLK(clknet_leaf_110_wb_clk_i),
    .D(_00381_),
    .Q(\tms1x00.ins_pla_ors[7][22] ));
 sky130_fd_sc_hd__dfxtp_2 _10577_ (.CLK(clknet_leaf_100_wb_clk_i),
    .D(_00382_),
    .Q(\tms1x00.ins_pla_ors[7][23] ));
 sky130_fd_sc_hd__dfxtp_1 _10578_ (.CLK(clknet_leaf_99_wb_clk_i),
    .D(_00383_),
    .Q(\tms1x00.ins_pla_ors[7][24] ));
 sky130_fd_sc_hd__dfxtp_1 _10579_ (.CLK(clknet_leaf_121_wb_clk_i),
    .D(_00384_),
    .Q(\tms1x00.ins_pla_ors[7][25] ));
 sky130_fd_sc_hd__dfxtp_1 _10580_ (.CLK(clknet_leaf_108_wb_clk_i),
    .D(_00385_),
    .Q(\tms1x00.ins_pla_ors[7][26] ));
 sky130_fd_sc_hd__dfxtp_1 _10581_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(_00386_),
    .Q(\tms1x00.ins_pla_ands[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10582_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(_00387_),
    .Q(\tms1x00.ins_pla_ands[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _10583_ (.CLK(clknet_leaf_56_wb_clk_i),
    .D(_00388_),
    .Q(\tms1x00.ins_pla_ands[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _10584_ (.CLK(clknet_leaf_56_wb_clk_i),
    .D(_00389_),
    .Q(\tms1x00.ins_pla_ands[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _10585_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(_00390_),
    .Q(\tms1x00.ins_pla_ands[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _10586_ (.CLK(clknet_leaf_56_wb_clk_i),
    .D(_00391_),
    .Q(\tms1x00.ins_pla_ands[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _10587_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(_00392_),
    .Q(\tms1x00.ins_pla_ands[5][8] ));
 sky130_fd_sc_hd__dfxtp_1 _10588_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(_00393_),
    .Q(\tms1x00.ins_pla_ands[5][9] ));
 sky130_fd_sc_hd__dfxtp_1 _10589_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(_00394_),
    .Q(\tms1x00.ins_pla_ands[5][10] ));
 sky130_fd_sc_hd__dfxtp_1 _10590_ (.CLK(clknet_leaf_56_wb_clk_i),
    .D(_00395_),
    .Q(\tms1x00.ins_pla_ands[5][11] ));
 sky130_fd_sc_hd__dfxtp_1 _10591_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(_00396_),
    .Q(\tms1x00.ins_pla_ands[4][0] ));
 sky130_fd_sc_hd__dfxtp_2 _10592_ (.CLK(clknet_leaf_88_wb_clk_i),
    .D(_00397_),
    .Q(\tms1x00.ins_pla_ands[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _10593_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(_00398_),
    .Q(\tms1x00.ins_pla_ands[4][5] ));
 sky130_fd_sc_hd__dfxtp_2 _10594_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(_00399_),
    .Q(\tms1x00.ins_pla_ands[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _10595_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(_00400_),
    .Q(\tms1x00.ins_pla_ands[4][12] ));
 sky130_fd_sc_hd__dfxtp_1 _10596_ (.CLK(clknet_leaf_58_wb_clk_i),
    .D(_00401_),
    .Q(\tms1x00.ins_pla_ands[4][13] ));
 sky130_fd_sc_hd__dfxtp_1 _10597_ (.CLK(clknet_leaf_139_wb_clk_i),
    .D(_00402_),
    .Q(\tms1x00.ins_pla_ands[28][9] ));
 sky130_fd_sc_hd__dfxtp_1 _10598_ (.CLK(clknet_leaf_130_wb_clk_i),
    .D(_00403_),
    .Q(\tms1x00.ins_pla_ands[28][10] ));
 sky130_fd_sc_hd__dfxtp_1 _10599_ (.CLK(clknet_leaf_138_wb_clk_i),
    .D(_00404_),
    .Q(\tms1x00.ins_pla_ands[28][13] ));
 sky130_fd_sc_hd__dfxtp_1 _10600_ (.CLK(clknet_leaf_142_wb_clk_i),
    .D(_00405_),
    .Q(\tms1x00.ins_pla_ands[28][14] ));
 sky130_fd_sc_hd__dfxtp_1 _10601_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_00406_),
    .Q(\tms1x00.ins_pla_ands[24][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10602_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_00407_),
    .Q(\tms1x00.ins_pla_ands[24][1] ));
 sky130_fd_sc_hd__dfxtp_1 _10603_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_00408_),
    .Q(\tms1x00.ins_pla_ands[24][2] ));
 sky130_fd_sc_hd__dfxtp_1 _10604_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_00409_),
    .Q(\tms1x00.ins_pla_ands[24][3] ));
 sky130_fd_sc_hd__dfxtp_1 _10605_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_00410_),
    .Q(\tms1x00.ins_pla_ands[24][10] ));
 sky130_fd_sc_hd__dfxtp_1 _10606_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_00411_),
    .Q(\tms1x00.ins_pla_ands[24][11] ));
 sky130_fd_sc_hd__dfxtp_1 _10607_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_00412_),
    .Q(\tms1x00.ins_pla_ands[21][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10608_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_00413_),
    .Q(\tms1x00.ins_pla_ands[21][1] ));
 sky130_fd_sc_hd__dfxtp_1 _10609_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_00414_),
    .Q(\tms1x00.ins_pla_ands[21][11] ));
 sky130_fd_sc_hd__dfxtp_1 _10610_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_00415_),
    .Q(\tms1x00.ins_pla_ands[20][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10611_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_00416_),
    .Q(\tms1x00.ins_pla_ands[20][1] ));
 sky130_fd_sc_hd__dfxtp_1 _10612_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_00417_),
    .Q(\tms1x00.ins_pla_ands[20][2] ));
 sky130_fd_sc_hd__dfxtp_1 _10613_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_00418_),
    .Q(\tms1x00.ins_pla_ands[20][3] ));
 sky130_fd_sc_hd__dfxtp_1 _10614_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_00419_),
    .Q(\tms1x00.ins_pla_ands[20][10] ));
 sky130_fd_sc_hd__dfxtp_1 _10615_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_00420_),
    .Q(\tms1x00.ins_pla_ands[20][11] ));
 sky130_fd_sc_hd__dfxtp_1 _10616_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_00421_),
    .Q(\tms1x00.ins_pla_ands[19][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10617_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_00422_),
    .Q(\tms1x00.ins_pla_ands[19][1] ));
 sky130_fd_sc_hd__dfxtp_1 _10618_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_00423_),
    .Q(\tms1x00.ins_pla_ands[19][10] ));
 sky130_fd_sc_hd__dfxtp_1 _10619_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_00424_),
    .Q(\tms1x00.ins_pla_ands[19][11] ));
 sky130_fd_sc_hd__dfxtp_1 _10620_ (.CLK(clknet_leaf_130_wb_clk_i),
    .D(_00425_),
    .Q(\tms1x00.ins_pla_ors[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _10621_ (.CLK(clknet_leaf_126_wb_clk_i),
    .D(_00426_),
    .Q(\tms1x00.ins_pla_ors[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 _10622_ (.CLK(clknet_leaf_126_wb_clk_i),
    .D(_00427_),
    .Q(\tms1x00.ins_pla_ors[11][8] ));
 sky130_fd_sc_hd__dfxtp_1 _10623_ (.CLK(clknet_leaf_127_wb_clk_i),
    .D(_00428_),
    .Q(\tms1x00.ins_pla_ors[11][9] ));
 sky130_fd_sc_hd__dfxtp_1 _10624_ (.CLK(clknet_leaf_131_wb_clk_i),
    .D(_00429_),
    .Q(\tms1x00.ins_pla_ors[11][10] ));
 sky130_fd_sc_hd__dfxtp_1 _10625_ (.CLK(clknet_leaf_129_wb_clk_i),
    .D(_00430_),
    .Q(\tms1x00.ins_pla_ors[11][11] ));
 sky130_fd_sc_hd__dfxtp_1 _10626_ (.CLK(clknet_leaf_130_wb_clk_i),
    .D(_00431_),
    .Q(\tms1x00.ins_pla_ors[11][12] ));
 sky130_fd_sc_hd__dfxtp_1 _10627_ (.CLK(clknet_leaf_113_wb_clk_i),
    .D(_00432_),
    .Q(\tms1x00.ins_pla_ors[11][20] ));
 sky130_fd_sc_hd__dfxtp_1 _10628_ (.CLK(clknet_leaf_117_wb_clk_i),
    .D(_00433_),
    .Q(\tms1x00.ins_pla_ors[11][23] ));
 sky130_fd_sc_hd__dfxtp_1 _10629_ (.CLK(clknet_leaf_125_wb_clk_i),
    .D(_00434_),
    .Q(\tms1x00.ins_pla_ors[11][24] ));
 sky130_fd_sc_hd__dfxtp_1 _10630_ (.CLK(clknet_leaf_120_wb_clk_i),
    .D(_00435_),
    .Q(\tms1x00.ins_pla_ors[11][27] ));
 sky130_fd_sc_hd__dfxtp_2 _10631_ (.CLK(clknet_leaf_113_wb_clk_i),
    .D(_00436_),
    .Q(\tms1x00.ins_pla_ors[11][28] ));
 sky130_fd_sc_hd__dfxtp_2 _10632_ (.CLK(clknet_leaf_122_wb_clk_i),
    .D(_00437_),
    .Q(\tms1x00.ins_pla_ors[11][29] ));
 sky130_fd_sc_hd__dfxtp_1 _10633_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_00438_),
    .Q(\tms1x00.ins_pla_ands[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10634_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_00439_),
    .Q(\tms1x00.ins_pla_ands[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _10635_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_00440_),
    .Q(\tms1x00.ins_pla_ands[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _10636_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_00441_),
    .Q(\tms1x00.ins_pla_ands[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _10637_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_00442_),
    .Q(\tms1x00.ins_pla_ands[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _10638_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_00443_),
    .Q(\tms1x00.ins_pla_ands[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _10639_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_00444_),
    .Q(\tms1x00.ins_pla_ands[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _10640_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_00445_),
    .Q(\tms1x00.ins_pla_ands[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _10641_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_00446_),
    .Q(\tms1x00.ins_pla_ands[7][8] ));
 sky130_fd_sc_hd__dfxtp_1 _10642_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_00447_),
    .Q(\tms1x00.ins_pla_ands[7][9] ));
 sky130_fd_sc_hd__dfxtp_1 _10643_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_00448_),
    .Q(\tms1x00.ins_pla_ands[7][10] ));
 sky130_fd_sc_hd__dfxtp_1 _10644_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_00449_),
    .Q(\tms1x00.ins_pla_ands[7][11] ));
 sky130_fd_sc_hd__dfxtp_1 _10645_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_00450_),
    .Q(\tms1x00.ins_pla_ands[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10646_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_00451_),
    .Q(\tms1x00.ins_pla_ands[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _10647_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_00452_),
    .Q(\tms1x00.ins_pla_ands[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _10648_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_00453_),
    .Q(\tms1x00.ins_pla_ands[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 _10649_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_00454_),
    .Q(\tms1x00.ins_pla_ands[8][7] ));
 sky130_fd_sc_hd__dfxtp_2 _10650_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_00455_),
    .Q(\tms1x00.ins_pla_ands[8][8] ));
 sky130_fd_sc_hd__dfxtp_2 _10651_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_00456_),
    .Q(\tms1x00.ins_pla_ands[8][9] ));
 sky130_fd_sc_hd__dfxtp_1 _10652_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_00457_),
    .Q(\tms1x00.ins_pla_ands[8][10] ));
 sky130_fd_sc_hd__dfxtp_1 _10653_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(_00458_),
    .Q(\tms1x00.ins_pla_ands[8][11] ));
 sky130_fd_sc_hd__dfxtp_1 _10654_ (.CLK(clknet_leaf_99_wb_clk_i),
    .D(_00459_),
    .Q(\tms1x00.ins_pla_ors[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10655_ (.CLK(clknet_leaf_97_wb_clk_i),
    .D(_00460_),
    .Q(\tms1x00.ins_pla_ors[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _10656_ (.CLK(clknet_leaf_96_wb_clk_i),
    .D(_00461_),
    .Q(\tms1x00.ins_pla_ors[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _10657_ (.CLK(clknet_leaf_91_wb_clk_i),
    .D(_00462_),
    .Q(\tms1x00.ins_pla_ors[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _10658_ (.CLK(clknet_leaf_98_wb_clk_i),
    .D(_00463_),
    .Q(\tms1x00.ins_pla_ors[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _10659_ (.CLK(clknet_leaf_99_wb_clk_i),
    .D(_00464_),
    .Q(\tms1x00.ins_pla_ors[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _10660_ (.CLK(clknet_leaf_96_wb_clk_i),
    .D(_00465_),
    .Q(\tms1x00.ins_pla_ors[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _10661_ (.CLK(clknet_leaf_92_wb_clk_i),
    .D(_00466_),
    .Q(\tms1x00.ins_pla_ors[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _10662_ (.CLK(clknet_leaf_101_wb_clk_i),
    .D(_00467_),
    .Q(\tms1x00.ins_pla_ors[1][9] ));
 sky130_fd_sc_hd__dfxtp_2 _10663_ (.CLK(clknet_leaf_108_wb_clk_i),
    .D(_00468_),
    .Q(\tms1x00.ins_pla_ors[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _10664_ (.CLK(clknet_leaf_91_wb_clk_i),
    .D(_00469_),
    .Q(\tms1x00.ins_pla_ors[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _10665_ (.CLK(clknet_leaf_106_wb_clk_i),
    .D(_00470_),
    .Q(\tms1x00.ins_pla_ors[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _10666_ (.CLK(clknet_leaf_98_wb_clk_i),
    .D(_00471_),
    .Q(\tms1x00.ins_pla_ors[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _10667_ (.CLK(clknet_leaf_107_wb_clk_i),
    .D(_00472_),
    .Q(\tms1x00.ins_pla_ors[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _10668_ (.CLK(clknet_leaf_106_wb_clk_i),
    .D(_00473_),
    .Q(\tms1x00.ins_pla_ors[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _10669_ (.CLK(clknet_leaf_102_wb_clk_i),
    .D(_00474_),
    .Q(\tms1x00.ins_pla_ors[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _10670_ (.CLK(clknet_leaf_102_wb_clk_i),
    .D(_00475_),
    .Q(\tms1x00.ins_pla_ors[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _10671_ (.CLK(clknet_leaf_101_wb_clk_i),
    .D(_00476_),
    .Q(\tms1x00.ins_pla_ors[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _10672_ (.CLK(clknet_leaf_106_wb_clk_i),
    .D(_00477_),
    .Q(\tms1x00.ins_pla_ors[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _10673_ (.CLK(clknet_leaf_107_wb_clk_i),
    .D(_00478_),
    .Q(\tms1x00.ins_pla_ors[1][20] ));
 sky130_fd_sc_hd__dfxtp_2 _10674_ (.CLK(clknet_leaf_108_wb_clk_i),
    .D(_00479_),
    .Q(\tms1x00.ins_pla_ors[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _10675_ (.CLK(clknet_leaf_111_wb_clk_i),
    .D(_00480_),
    .Q(\tms1x00.ins_pla_ors[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _10676_ (.CLK(clknet_leaf_101_wb_clk_i),
    .D(_00481_),
    .Q(\tms1x00.ins_pla_ors[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _10677_ (.CLK(clknet_leaf_99_wb_clk_i),
    .D(_00482_),
    .Q(\tms1x00.ins_pla_ors[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _10678_ (.CLK(clknet_leaf_93_wb_clk_i),
    .D(_00483_),
    .Q(\tms1x00.ins_pla_ors[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _10679_ (.CLK(clknet_leaf_108_wb_clk_i),
    .D(_00484_),
    .Q(\tms1x00.ins_pla_ors[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _10680_ (.CLK(clknet_leaf_111_wb_clk_i),
    .D(_00485_),
    .Q(\tms1x00.ins_pla_ors[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _10681_ (.CLK(clknet_leaf_106_wb_clk_i),
    .D(_00486_),
    .Q(\tms1x00.ins_pla_ors[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _10682_ (.CLK(clknet_leaf_124_wb_clk_i),
    .D(_00487_),
    .Q(\tms1x00.ins_pla_ors[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _10683_ (.CLK(clknet_leaf_125_wb_clk_i),
    .D(_00488_),
    .Q(\tms1x00.ins_pla_ors[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _10684_ (.CLK(clknet_leaf_123_wb_clk_i),
    .D(_00489_),
    .Q(\tms1x00.ins_pla_ors[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _10685_ (.CLK(clknet_leaf_127_wb_clk_i),
    .D(_00490_),
    .Q(\tms1x00.ins_pla_ors[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 _10686_ (.CLK(clknet_leaf_125_wb_clk_i),
    .D(_00491_),
    .Q(\tms1x00.ins_pla_ors[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 _10687_ (.CLK(clknet_leaf_90_wb_clk_i),
    .D(_00492_),
    .Q(\tms1x00.ins_pla_ors[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 _10688_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_00493_),
    .Q(\tms1x00.ins_pla_ors[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 _10689_ (.CLK(clknet_leaf_118_wb_clk_i),
    .D(_00494_),
    .Q(\tms1x00.ins_pla_ors[13][10] ));
 sky130_fd_sc_hd__dfxtp_1 _10690_ (.CLK(clknet_leaf_128_wb_clk_i),
    .D(_00495_),
    .Q(\tms1x00.ins_pla_ors[13][12] ));
 sky130_fd_sc_hd__dfxtp_1 _10691_ (.CLK(clknet_leaf_128_wb_clk_i),
    .D(_00496_),
    .Q(\tms1x00.ins_pla_ors[13][13] ));
 sky130_fd_sc_hd__dfxtp_1 _10692_ (.CLK(clknet_leaf_121_wb_clk_i),
    .D(_00497_),
    .Q(\tms1x00.ins_pla_ors[13][17] ));
 sky130_fd_sc_hd__dfxtp_1 _10693_ (.CLK(clknet_leaf_128_wb_clk_i),
    .D(_00498_),
    .Q(\tms1x00.ins_pla_ors[13][19] ));
 sky130_fd_sc_hd__dfxtp_1 _10694_ (.CLK(clknet_leaf_115_wb_clk_i),
    .D(_00499_),
    .Q(\tms1x00.ins_pla_ors[13][22] ));
 sky130_fd_sc_hd__dfxtp_1 _10695_ (.CLK(clknet_leaf_119_wb_clk_i),
    .D(_00500_),
    .Q(\tms1x00.ins_pla_ors[13][23] ));
 sky130_fd_sc_hd__dfxtp_1 _10696_ (.CLK(clknet_leaf_122_wb_clk_i),
    .D(_00501_),
    .Q(\tms1x00.ins_pla_ors[13][24] ));
 sky130_fd_sc_hd__dfxtp_1 _10697_ (.CLK(clknet_leaf_81_wb_clk_i),
    .D(_00502_),
    .Q(\tms1x00.ins_pla_ors[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10698_ (.CLK(clknet_leaf_83_wb_clk_i),
    .D(_00503_),
    .Q(\tms1x00.ins_pla_ors[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _10699_ (.CLK(clknet_leaf_83_wb_clk_i),
    .D(_00504_),
    .Q(\tms1x00.ins_pla_ors[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _10700_ (.CLK(clknet_leaf_93_wb_clk_i),
    .D(_00505_),
    .Q(\tms1x00.ins_pla_ors[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _10701_ (.CLK(clknet_leaf_82_wb_clk_i),
    .D(_00506_),
    .Q(\tms1x00.ins_pla_ors[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _10702_ (.CLK(clknet_leaf_101_wb_clk_i),
    .D(_00507_),
    .Q(\tms1x00.ins_pla_ors[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _10703_ (.CLK(clknet_leaf_102_wb_clk_i),
    .D(_00508_),
    .Q(\tms1x00.ins_pla_ors[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _10704_ (.CLK(clknet_leaf_99_wb_clk_i),
    .D(_00509_),
    .Q(\tms1x00.ins_pla_ors[6][9] ));
 sky130_fd_sc_hd__dfxtp_1 _10705_ (.CLK(clknet_leaf_99_wb_clk_i),
    .D(_00510_),
    .Q(\tms1x00.ins_pla_ors[6][10] ));
 sky130_fd_sc_hd__dfxtp_1 _10706_ (.CLK(clknet_leaf_104_wb_clk_i),
    .D(_00511_),
    .Q(\tms1x00.ins_pla_ors[6][11] ));
 sky130_fd_sc_hd__dfxtp_1 _10707_ (.CLK(clknet_leaf_81_wb_clk_i),
    .D(_00512_),
    .Q(\tms1x00.ins_pla_ors[6][13] ));
 sky130_fd_sc_hd__dfxtp_2 _10708_ (.CLK(clknet_leaf_107_wb_clk_i),
    .D(_00513_),
    .Q(\tms1x00.ins_pla_ors[6][14] ));
 sky130_fd_sc_hd__dfxtp_1 _10709_ (.CLK(clknet_leaf_106_wb_clk_i),
    .D(_00514_),
    .Q(\tms1x00.ins_pla_ors[6][15] ));
 sky130_fd_sc_hd__dfxtp_1 _10710_ (.CLK(clknet_leaf_108_wb_clk_i),
    .D(_00515_),
    .Q(\tms1x00.ins_pla_ors[6][17] ));
 sky130_fd_sc_hd__dfxtp_2 _10711_ (.CLK(clknet_leaf_107_wb_clk_i),
    .D(_00516_),
    .Q(\tms1x00.ins_pla_ors[6][19] ));
 sky130_fd_sc_hd__dfxtp_1 _10712_ (.CLK(clknet_leaf_108_wb_clk_i),
    .D(_00517_),
    .Q(\tms1x00.ins_pla_ors[6][20] ));
 sky130_fd_sc_hd__dfxtp_1 _10713_ (.CLK(clknet_leaf_108_wb_clk_i),
    .D(_00518_),
    .Q(\tms1x00.ins_pla_ors[6][21] ));
 sky130_fd_sc_hd__dfxtp_1 _10714_ (.CLK(clknet_leaf_110_wb_clk_i),
    .D(_00519_),
    .Q(\tms1x00.ins_pla_ors[6][22] ));
 sky130_fd_sc_hd__dfxtp_1 _10715_ (.CLK(clknet_leaf_101_wb_clk_i),
    .D(_00520_),
    .Q(\tms1x00.ins_pla_ors[6][23] ));
 sky130_fd_sc_hd__dfxtp_1 _10716_ (.CLK(clknet_leaf_99_wb_clk_i),
    .D(_00521_),
    .Q(\tms1x00.ins_pla_ors[6][24] ));
 sky130_fd_sc_hd__dfxtp_1 _10717_ (.CLK(clknet_leaf_128_wb_clk_i),
    .D(_00522_),
    .Q(\tms1x00.ins_pla_ors[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10718_ (.CLK(clknet_leaf_131_wb_clk_i),
    .D(_00523_),
    .Q(\tms1x00.ins_pla_ors[10][2] ));
 sky130_fd_sc_hd__dfxtp_2 _10719_ (.CLK(clknet_leaf_134_wb_clk_i),
    .D(_00524_),
    .Q(\tms1x00.ins_pla_ors[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 _10720_ (.CLK(clknet_leaf_123_wb_clk_i),
    .D(_00525_),
    .Q(\tms1x00.ins_pla_ors[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 _10721_ (.CLK(clknet_leaf_127_wb_clk_i),
    .D(_00526_),
    .Q(\tms1x00.ins_pla_ors[10][8] ));
 sky130_fd_sc_hd__dfxtp_1 _10722_ (.CLK(clknet_leaf_127_wb_clk_i),
    .D(_00527_),
    .Q(\tms1x00.ins_pla_ors[10][9] ));
 sky130_fd_sc_hd__dfxtp_1 _10723_ (.CLK(clknet_leaf_131_wb_clk_i),
    .D(_00528_),
    .Q(\tms1x00.ins_pla_ors[10][10] ));
 sky130_fd_sc_hd__dfxtp_1 _10724_ (.CLK(clknet_leaf_127_wb_clk_i),
    .D(_00529_),
    .Q(\tms1x00.ins_pla_ors[10][11] ));
 sky130_fd_sc_hd__dfxtp_1 _10725_ (.CLK(clknet_leaf_128_wb_clk_i),
    .D(_00530_),
    .Q(\tms1x00.ins_pla_ors[10][12] ));
 sky130_fd_sc_hd__dfxtp_1 _10726_ (.CLK(clknet_leaf_131_wb_clk_i),
    .D(_00531_),
    .Q(\tms1x00.ins_pla_ors[10][13] ));
 sky130_fd_sc_hd__dfxtp_1 _10727_ (.CLK(clknet_leaf_131_wb_clk_i),
    .D(_00532_),
    .Q(\tms1x00.ins_pla_ors[10][14] ));
 sky130_fd_sc_hd__dfxtp_1 _10728_ (.CLK(clknet_leaf_132_wb_clk_i),
    .D(_00533_),
    .Q(\tms1x00.ins_pla_ors[10][15] ));
 sky130_fd_sc_hd__dfxtp_1 _10729_ (.CLK(clknet_leaf_122_wb_clk_i),
    .D(_00534_),
    .Q(\tms1x00.ins_pla_ors[10][16] ));
 sky130_fd_sc_hd__dfxtp_1 _10730_ (.CLK(clknet_leaf_122_wb_clk_i),
    .D(_00535_),
    .Q(\tms1x00.ins_pla_ors[10][18] ));
 sky130_fd_sc_hd__dfxtp_1 _10731_ (.CLK(clknet_leaf_115_wb_clk_i),
    .D(_00536_),
    .Q(\tms1x00.ins_pla_ors[10][20] ));
 sky130_fd_sc_hd__dfxtp_1 _10732_ (.CLK(clknet_leaf_134_wb_clk_i),
    .D(_00537_),
    .Q(\tms1x00.ins_pla_ors[10][21] ));
 sky130_fd_sc_hd__dfxtp_1 _10733_ (.CLK(clknet_leaf_117_wb_clk_i),
    .D(_00538_),
    .Q(\tms1x00.ins_pla_ors[10][22] ));
 sky130_fd_sc_hd__dfxtp_1 _10734_ (.CLK(clknet_leaf_117_wb_clk_i),
    .D(_00539_),
    .Q(\tms1x00.ins_pla_ors[10][23] ));
 sky130_fd_sc_hd__dfxtp_1 _10735_ (.CLK(clknet_leaf_118_wb_clk_i),
    .D(_00540_),
    .Q(\tms1x00.ins_pla_ors[10][25] ));
 sky130_fd_sc_hd__dfxtp_1 _10736_ (.CLK(clknet_leaf_120_wb_clk_i),
    .D(_00541_),
    .Q(\tms1x00.ins_pla_ors[10][27] ));
 sky130_fd_sc_hd__dfxtp_2 _10737_ (.CLK(clknet_leaf_122_wb_clk_i),
    .D(_00542_),
    .Q(\tms1x00.ins_pla_ors[10][29] ));
 sky130_fd_sc_hd__dfxtp_1 _10738_ (.CLK(clknet_leaf_139_wb_clk_i),
    .D(_00543_),
    .Q(\tms1x00.ins_pla_ands[29][8] ));
 sky130_fd_sc_hd__dfxtp_1 _10739_ (.CLK(clknet_leaf_130_wb_clk_i),
    .D(_00544_),
    .Q(\tms1x00.ins_pla_ands[29][10] ));
 sky130_fd_sc_hd__dfxtp_1 _10740_ (.CLK(clknet_leaf_138_wb_clk_i),
    .D(_00545_),
    .Q(\tms1x00.ins_pla_ands[29][13] ));
 sky130_fd_sc_hd__dfxtp_1 _10741_ (.CLK(clknet_leaf_138_wb_clk_i),
    .D(_00546_),
    .Q(\tms1x00.ins_pla_ands[29][14] ));
 sky130_fd_sc_hd__dfxtp_2 _10742_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_00547_),
    .Q(\tms1x00.ins_pla_ands[25][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10743_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_00548_),
    .Q(\tms1x00.ins_pla_ands[25][1] ));
 sky130_fd_sc_hd__dfxtp_1 _10744_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_00549_),
    .Q(\tms1x00.ins_pla_ands[25][10] ));
 sky130_fd_sc_hd__dfxtp_1 _10745_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_00550_),
    .Q(\tms1x00.ins_pla_ands[25][11] ));
 sky130_fd_sc_hd__dfxtp_1 _10746_ (.CLK(clknet_leaf_99_wb_clk_i),
    .D(_00551_),
    .Q(\tms1x00.ins_pla_ors[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10747_ (.CLK(clknet_leaf_95_wb_clk_i),
    .D(_00552_),
    .Q(\tms1x00.ins_pla_ors[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _10748_ (.CLK(clknet_leaf_96_wb_clk_i),
    .D(_00553_),
    .Q(\tms1x00.ins_pla_ors[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _10749_ (.CLK(clknet_leaf_83_wb_clk_i),
    .D(_00554_),
    .Q(\tms1x00.ins_pla_ors[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _10750_ (.CLK(clknet_leaf_83_wb_clk_i),
    .D(_00555_),
    .Q(\tms1x00.ins_pla_ors[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _10751_ (.CLK(clknet_leaf_83_wb_clk_i),
    .D(_00556_),
    .Q(\tms1x00.ins_pla_ors[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _10752_ (.CLK(clknet_leaf_94_wb_clk_i),
    .D(_00557_),
    .Q(\tms1x00.ins_pla_ors[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _10753_ (.CLK(clknet_leaf_100_wb_clk_i),
    .D(_00558_),
    .Q(\tms1x00.ins_pla_ors[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _10754_ (.CLK(clknet_leaf_83_wb_clk_i),
    .D(_00559_),
    .Q(\tms1x00.ins_pla_ors[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _10755_ (.CLK(clknet_leaf_81_wb_clk_i),
    .D(_00560_),
    .Q(\tms1x00.ins_pla_ors[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _10756_ (.CLK(clknet_leaf_107_wb_clk_i),
    .D(_00561_),
    .Q(\tms1x00.ins_pla_ors[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _10757_ (.CLK(clknet_leaf_104_wb_clk_i),
    .D(_00562_),
    .Q(\tms1x00.ins_pla_ors[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _10758_ (.CLK(clknet_leaf_103_wb_clk_i),
    .D(_00563_),
    .Q(\tms1x00.ins_pla_ors[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _10759_ (.CLK(clknet_leaf_103_wb_clk_i),
    .D(_00564_),
    .Q(\tms1x00.ins_pla_ors[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _10760_ (.CLK(clknet_leaf_100_wb_clk_i),
    .D(_00565_),
    .Q(\tms1x00.ins_pla_ors[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _10761_ (.CLK(clknet_leaf_106_wb_clk_i),
    .D(_00566_),
    .Q(\tms1x00.ins_pla_ors[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _10762_ (.CLK(clknet_leaf_107_wb_clk_i),
    .D(_00567_),
    .Q(\tms1x00.ins_pla_ors[0][20] ));
 sky130_fd_sc_hd__dfxtp_2 _10763_ (.CLK(clknet_leaf_108_wb_clk_i),
    .D(_00568_),
    .Q(\tms1x00.ins_pla_ors[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _10764_ (.CLK(clknet_leaf_110_wb_clk_i),
    .D(_00569_),
    .Q(\tms1x00.ins_pla_ors[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _10765_ (.CLK(clknet_leaf_99_wb_clk_i),
    .D(_00570_),
    .Q(\tms1x00.ins_pla_ors[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _10766_ (.CLK(clknet_leaf_111_wb_clk_i),
    .D(_00571_),
    .Q(\tms1x00.ins_pla_ors[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _10767_ (.CLK(clknet_leaf_112_wb_clk_i),
    .D(_00572_),
    .Q(\tms1x00.ins_pla_ors[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _10768_ (.CLK(clknet_leaf_111_wb_clk_i),
    .D(_00573_),
    .Q(\tms1x00.ins_pla_ors[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _10769_ (.CLK(clknet_leaf_110_wb_clk_i),
    .D(_00574_),
    .Q(\tms1x00.ins_pla_ors[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _10770_ (.CLK(clknet_leaf_97_wb_clk_i),
    .D(_00575_),
    .Q(\tms1x00.ins_pla_ors[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _10771_ (.CLK(clknet_leaf_91_wb_clk_i),
    .D(_00576_),
    .Q(\tms1x00.ins_pla_ors[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _10772_ (.CLK(clknet_leaf_93_wb_clk_i),
    .D(_00577_),
    .Q(\tms1x00.ins_pla_ors[5][6] ));
 sky130_fd_sc_hd__dfxtp_2 _10773_ (.CLK(clknet_leaf_102_wb_clk_i),
    .D(_00578_),
    .Q(\tms1x00.ins_pla_ors[5][9] ));
 sky130_fd_sc_hd__dfxtp_2 _10774_ (.CLK(clknet_leaf_92_wb_clk_i),
    .D(_00579_),
    .Q(\tms1x00.ins_pla_ors[5][10] ));
 sky130_fd_sc_hd__dfxtp_1 _10775_ (.CLK(clknet_leaf_104_wb_clk_i),
    .D(_00580_),
    .Q(\tms1x00.ins_pla_ors[5][11] ));
 sky130_fd_sc_hd__dfxtp_1 _10776_ (.CLK(clknet_leaf_105_wb_clk_i),
    .D(_00581_),
    .Q(\tms1x00.ins_pla_ors[5][12] ));
 sky130_fd_sc_hd__dfxtp_1 _10777_ (.CLK(clknet_leaf_90_wb_clk_i),
    .D(_00582_),
    .Q(\tms1x00.ins_pla_ors[5][13] ));
 sky130_fd_sc_hd__dfxtp_2 _10778_ (.CLK(clknet_leaf_107_wb_clk_i),
    .D(_00583_),
    .Q(\tms1x00.ins_pla_ors[5][14] ));
 sky130_fd_sc_hd__dfxtp_1 _10779_ (.CLK(clknet_leaf_106_wb_clk_i),
    .D(_00584_),
    .Q(\tms1x00.ins_pla_ors[5][15] ));
 sky130_fd_sc_hd__dfxtp_2 _10780_ (.CLK(clknet_leaf_103_wb_clk_i),
    .D(_00585_),
    .Q(\tms1x00.ins_pla_ors[5][17] ));
 sky130_fd_sc_hd__dfxtp_1 _10781_ (.CLK(clknet_leaf_121_wb_clk_i),
    .D(_00586_),
    .Q(\tms1x00.ins_pla_ors[5][18] ));
 sky130_fd_sc_hd__dfxtp_2 _10782_ (.CLK(clknet_leaf_107_wb_clk_i),
    .D(_00587_),
    .Q(\tms1x00.ins_pla_ors[5][19] ));
 sky130_fd_sc_hd__dfxtp_2 _10783_ (.CLK(clknet_leaf_104_wb_clk_i),
    .D(_00588_),
    .Q(\tms1x00.ins_pla_ors[5][20] ));
 sky130_fd_sc_hd__dfxtp_1 _10784_ (.CLK(clknet_leaf_111_wb_clk_i),
    .D(_00589_),
    .Q(\tms1x00.ins_pla_ors[5][22] ));
 sky130_fd_sc_hd__dfxtp_2 _10785_ (.CLK(clknet_leaf_101_wb_clk_i),
    .D(_00590_),
    .Q(\tms1x00.ins_pla_ors[5][23] ));
 sky130_fd_sc_hd__dfxtp_1 _10786_ (.CLK(clknet_leaf_121_wb_clk_i),
    .D(_00591_),
    .Q(\tms1x00.ins_pla_ors[5][25] ));
 sky130_fd_sc_hd__dfxtp_1 _10787_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(_00592_),
    .Q(\tms1x00.ins_pla_ands[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _10788_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(_00593_),
    .Q(\tms1x00.ins_pla_ands[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _10789_ (.CLK(clknet_leaf_54_wb_clk_i),
    .D(_00594_),
    .Q(\tms1x00.ins_pla_ands[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _10790_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(_00595_),
    .Q(\tms1x00.ins_pla_ands[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _10791_ (.CLK(clknet_leaf_54_wb_clk_i),
    .D(_00596_),
    .Q(\tms1x00.ins_pla_ands[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _10792_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(_00597_),
    .Q(\tms1x00.ins_pla_ands[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _10793_ (.CLK(clknet_leaf_54_wb_clk_i),
    .D(_00598_),
    .Q(\tms1x00.ins_pla_ands[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _10794_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(_00599_),
    .Q(\tms1x00.ins_pla_ands[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _10795_ (.CLK(clknet_leaf_127_wb_clk_i),
    .D(_00600_),
    .Q(\tms1x00.ins_pla_ors[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _10796_ (.CLK(clknet_leaf_119_wb_clk_i),
    .D(_00601_),
    .Q(\tms1x00.ins_pla_ors[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _10797_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_00602_),
    .Q(\tms1x00.ins_pla_ors[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 _10798_ (.CLK(clknet_leaf_127_wb_clk_i),
    .D(_00603_),
    .Q(\tms1x00.ins_pla_ors[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 _10799_ (.CLK(clknet_leaf_121_wb_clk_i),
    .D(_00604_),
    .Q(\tms1x00.ins_pla_ors[10][17] ));
 sky130_fd_sc_hd__dfxtp_1 _10800_ (.CLK(clknet_leaf_132_wb_clk_i),
    .D(_00605_),
    .Q(\tms1x00.ins_pla_ors[10][19] ));
 sky130_fd_sc_hd__dfxtp_1 _10801_ (.CLK(clknet_leaf_124_wb_clk_i),
    .D(_00606_),
    .Q(\tms1x00.ins_pla_ors[10][24] ));
 sky130_fd_sc_hd__dfxtp_1 _10802_ (.CLK(clknet_leaf_116_wb_clk_i),
    .D(_00607_),
    .Q(\tms1x00.ins_pla_ors[10][26] ));
 sky130_fd_sc_hd__dfxtp_2 _10803_ (.CLK(clknet_leaf_113_wb_clk_i),
    .D(_00608_),
    .Q(\tms1x00.ins_pla_ors[10][28] ));
 sky130_fd_sc_hd__dfxtp_1 _10804_ (.CLK(clknet_leaf_95_wb_clk_i),
    .D(_00609_),
    .Q(\tms1x00.ins_pla_ors[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _10805_ (.CLK(clknet_leaf_97_wb_clk_i),
    .D(_00610_),
    .Q(\tms1x00.ins_pla_ors[0][6] ));
 sky130_fd_sc_hd__dfxtp_2 _10806_ (.CLK(clknet_leaf_106_wb_clk_i),
    .D(_00611_),
    .Q(\tms1x00.ins_pla_ors[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _10807_ (.CLK(clknet_leaf_112_wb_clk_i),
    .D(_00612_),
    .Q(\tms1x00.ins_pla_ors[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _10808_ (.CLK(clknet_leaf_100_wb_clk_i),
    .D(_00613_),
    .Q(\tms1x00.ins_pla_ors[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _10809_ (.CLK(clknet_leaf_94_wb_clk_i),
    .D(_00614_),
    .Q(\tms1x00.ins_pla_ors[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _10810_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_00615_),
    .Q(\tms1x00.ins_pla_ands[23][2] ));
 sky130_fd_sc_hd__dfxtp_1 _10811_ (.CLK(clknet_leaf_129_wb_clk_i),
    .D(_00616_),
    .Q(\tms1x00.ins_pla_ands[23][3] ));
 sky130_fd_sc_hd__dfxtp_1 _10812_ (.CLK(clknet_leaf_129_wb_clk_i),
    .D(_00617_),
    .Q(\tms1x00.ins_pla_ands[23][4] ));
 sky130_fd_sc_hd__dfxtp_1 _10813_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_00618_),
    .Q(\tms1x00.ins_pla_ands[23][5] ));
 sky130_fd_sc_hd__dfxtp_1 _10814_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_00619_),
    .Q(\tms1x00.ins_pla_ands[23][6] ));
 sky130_fd_sc_hd__dfxtp_1 _10815_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_00620_),
    .Q(\tms1x00.ins_pla_ands[23][7] ));
 sky130_fd_sc_hd__dfxtp_1 _10816_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_00621_),
    .Q(\tms1x00.ins_pla_ands[23][8] ));
 sky130_fd_sc_hd__dfxtp_1 _10817_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_00622_),
    .Q(\tms1x00.ins_pla_ands[23][9] ));
 sky130_fd_sc_hd__dfxtp_1 _10818_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_00623_),
    .Q(\tms1x00.ins_pla_ands[23][12] ));
 sky130_fd_sc_hd__dfxtp_1 _10819_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_00624_),
    .Q(\tms1x00.ins_pla_ands[23][13] ));
 sky130_fd_sc_hd__dfxtp_1 _10820_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_00625_),
    .Q(\tms1x00.ins_pla_ands[23][14] ));
 sky130_fd_sc_hd__dfxtp_1 _10821_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_00626_),
    .Q(\tms1x00.ins_pla_ands[23][15] ));
 sky130_fd_sc_hd__dfxtp_1 _10822_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_00627_),
    .Q(\tms1x00.ins_pla_ands[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _10823_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_00628_),
    .Q(\tms1x00.ins_pla_ands[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _10824_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_00629_),
    .Q(\tms1x00.ins_pla_ands[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 _10825_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_00630_),
    .Q(\tms1x00.ins_pla_ands[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 _10826_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_00631_),
    .Q(\tms1x00.ins_pla_ands[14][8] ));
 sky130_fd_sc_hd__dfxtp_1 _10827_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_00632_),
    .Q(\tms1x00.ins_pla_ands[14][9] ));
 sky130_fd_sc_hd__dfxtp_1 _10828_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_00633_),
    .Q(\tms1x00.ins_pla_ands[14][10] ));
 sky130_fd_sc_hd__dfxtp_1 _10829_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_00634_),
    .Q(\tms1x00.ins_pla_ands[14][11] ));
 sky130_fd_sc_hd__dfxtp_1 _10830_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_00635_),
    .Q(\tms1x00.ins_pla_ands[14][12] ));
 sky130_fd_sc_hd__dfxtp_1 _10831_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_00636_),
    .Q(\tms1x00.ins_pla_ands[14][13] ));
 sky130_fd_sc_hd__dfxtp_1 _10832_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_00637_),
    .Q(\tms1x00.ins_pla_ands[14][14] ));
 sky130_fd_sc_hd__dfxtp_1 _10833_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_00638_),
    .Q(\tms1x00.ins_pla_ands[14][15] ));
 sky130_fd_sc_hd__dfxtp_1 _10834_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(_00639_),
    .Q(\tms1x00.ins_pla_ands[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _10835_ (.CLK(clknet_leaf_88_wb_clk_i),
    .D(_00640_),
    .Q(\tms1x00.ins_pla_ands[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _10836_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(_00641_),
    .Q(\tms1x00.ins_pla_ands[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _10837_ (.CLK(clknet_leaf_88_wb_clk_i),
    .D(_00642_),
    .Q(\tms1x00.ins_pla_ands[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _10838_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(_00643_),
    .Q(\tms1x00.ins_pla_ands[4][8] ));
 sky130_fd_sc_hd__dfxtp_1 _10839_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(_00644_),
    .Q(\tms1x00.ins_pla_ands[4][9] ));
 sky130_fd_sc_hd__dfxtp_1 _10840_ (.CLK(clknet_leaf_88_wb_clk_i),
    .D(_00645_),
    .Q(\tms1x00.ins_pla_ands[4][10] ));
 sky130_fd_sc_hd__dfxtp_1 _10841_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(_00646_),
    .Q(\tms1x00.ins_pla_ands[4][11] ));
 sky130_fd_sc_hd__dfxtp_1 _10842_ (.CLK(clknet_leaf_62_wb_clk_i),
    .D(_00647_),
    .Q(\tms1x00.ins_pla_ands[4][14] ));
 sky130_fd_sc_hd__dfxtp_1 _10843_ (.CLK(clknet_leaf_62_wb_clk_i),
    .D(_00648_),
    .Q(\tms1x00.ins_pla_ands[4][15] ));
 sky130_fd_sc_hd__dfxtp_1 _10844_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_00649_),
    .Q(\tms1x00.ins_pla_ands[22][6] ));
 sky130_fd_sc_hd__dfxtp_1 _10845_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_00650_),
    .Q(\tms1x00.ins_pla_ands[22][7] ));
 sky130_fd_sc_hd__dfxtp_1 _10846_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_00651_),
    .Q(\tms1x00.ins_pla_ands[22][8] ));
 sky130_fd_sc_hd__dfxtp_1 _10847_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_00652_),
    .Q(\tms1x00.ins_pla_ands[22][9] ));
 sky130_fd_sc_hd__dfxtp_1 _10848_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_00653_),
    .Q(\tms1x00.ins_pla_ands[22][10] ));
 sky130_fd_sc_hd__dfxtp_1 _10849_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_00654_),
    .Q(\tms1x00.ins_pla_ands[22][12] ));
 sky130_fd_sc_hd__dfxtp_1 _10850_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_00655_),
    .Q(\tms1x00.ins_pla_ands[22][13] ));
 sky130_fd_sc_hd__dfxtp_1 _10851_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_00656_),
    .Q(\tms1x00.ins_pla_ands[22][14] ));
 sky130_fd_sc_hd__dfxtp_1 _10852_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_00657_),
    .Q(\tms1x00.ins_pla_ands[22][15] ));
 sky130_fd_sc_hd__dfxtp_1 _10853_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_00658_),
    .Q(\tms1x00.ins_pla_ands[13][8] ));
 sky130_fd_sc_hd__dfxtp_1 _10854_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_00659_),
    .Q(\tms1x00.ins_pla_ands[13][9] ));
 sky130_fd_sc_hd__dfxtp_1 _10855_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_00660_),
    .Q(\tms1x00.ins_pla_ands[13][10] ));
 sky130_fd_sc_hd__dfxtp_1 _10856_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_00661_),
    .Q(\tms1x00.ins_pla_ands[13][11] ));
 sky130_fd_sc_hd__dfxtp_1 _10857_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_00662_),
    .Q(\tms1x00.ins_pla_ands[13][12] ));
 sky130_fd_sc_hd__dfxtp_1 _10858_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_00663_),
    .Q(\tms1x00.ins_pla_ands[13][13] ));
 sky130_fd_sc_hd__dfxtp_1 _10859_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_00664_),
    .Q(\tms1x00.ins_pla_ands[13][14] ));
 sky130_fd_sc_hd__dfxtp_1 _10860_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_00665_),
    .Q(\tms1x00.ins_pla_ands[13][15] ));
 sky130_fd_sc_hd__dfxtp_1 _10861_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(_00666_),
    .Q(\tms1x00.ins_pla_ands[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10862_ (.CLK(clknet_leaf_56_wb_clk_i),
    .D(_00667_),
    .Q(\tms1x00.ins_pla_ands[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _10863_ (.CLK(clknet_leaf_58_wb_clk_i),
    .D(_00668_),
    .Q(\tms1x00.ins_pla_ands[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _10864_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(_00669_),
    .Q(\tms1x00.ins_pla_ands[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _10865_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_00670_),
    .Q(\tms1x00.ins_pla_ands[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _10866_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(_00671_),
    .Q(\tms1x00.ins_pla_ands[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _10867_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_00672_),
    .Q(\tms1x00.ins_pla_ands[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _10868_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_00673_),
    .Q(\tms1x00.ins_pla_ands[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _10869_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_00674_),
    .Q(\tms1x00.ins_pla_ands[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10870_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_00675_),
    .Q(\tms1x00.ins_pla_ands[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _10871_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_00676_),
    .Q(\tms1x00.ins_pla_ands[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 _10872_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_00677_),
    .Q(\tms1x00.ins_pla_ands[14][7] ));
 sky130_fd_sc_hd__dfxtp_1 _10873_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_00678_),
    .Q(\tms1x00.ins_pla_ands[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 _10874_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_00679_),
    .Q(\tms1x00.ins_pla_ands[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 _10875_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_00680_),
    .Q(\tms1x00.ins_pla_ands[21][2] ));
 sky130_fd_sc_hd__dfxtp_1 _10876_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_00681_),
    .Q(\tms1x00.ins_pla_ands[21][3] ));
 sky130_fd_sc_hd__dfxtp_1 _10877_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_00682_),
    .Q(\tms1x00.ins_pla_ands[21][4] ));
 sky130_fd_sc_hd__dfxtp_1 _10878_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_00683_),
    .Q(\tms1x00.ins_pla_ands[21][5] ));
 sky130_fd_sc_hd__dfxtp_1 _10879_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_00684_),
    .Q(\tms1x00.ins_pla_ands[21][6] ));
 sky130_fd_sc_hd__dfxtp_1 _10880_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_00685_),
    .Q(\tms1x00.ins_pla_ands[21][7] ));
 sky130_fd_sc_hd__dfxtp_1 _10881_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_00686_),
    .Q(\tms1x00.ins_pla_ands[21][8] ));
 sky130_fd_sc_hd__dfxtp_1 _10882_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_00687_),
    .Q(\tms1x00.ins_pla_ands[21][9] ));
 sky130_fd_sc_hd__dfxtp_1 _10883_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_00688_),
    .Q(\tms1x00.ins_pla_ands[21][10] ));
 sky130_fd_sc_hd__dfxtp_1 _10884_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_00689_),
    .Q(\tms1x00.ins_pla_ands[21][12] ));
 sky130_fd_sc_hd__dfxtp_1 _10885_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_00690_),
    .Q(\tms1x00.ins_pla_ands[21][13] ));
 sky130_fd_sc_hd__dfxtp_1 _10886_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_00691_),
    .Q(\tms1x00.ins_pla_ands[21][14] ));
 sky130_fd_sc_hd__dfxtp_1 _10887_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_00692_),
    .Q(\tms1x00.ins_pla_ands[21][15] ));
 sky130_fd_sc_hd__dfxtp_1 _10888_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_00693_),
    .Q(\tms1x00.ins_pla_ands[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10889_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_00694_),
    .Q(\tms1x00.ins_pla_ands[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _10890_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_00695_),
    .Q(\tms1x00.ins_pla_ands[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _10891_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_00696_),
    .Q(\tms1x00.ins_pla_ands[12][4] ));
 sky130_fd_sc_hd__dfxtp_2 _10892_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_00697_),
    .Q(\tms1x00.ins_pla_ands[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 _10893_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_00698_),
    .Q(\tms1x00.ins_pla_ands[12][8] ));
 sky130_fd_sc_hd__dfxtp_1 _10894_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_00699_),
    .Q(\tms1x00.ins_pla_ands[12][9] ));
 sky130_fd_sc_hd__dfxtp_1 _10895_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_00700_),
    .Q(\tms1x00.ins_pla_ands[12][10] ));
 sky130_fd_sc_hd__dfxtp_1 _10896_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_00701_),
    .Q(\tms1x00.ins_pla_ands[12][11] ));
 sky130_fd_sc_hd__dfxtp_1 _10897_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_00702_),
    .Q(\tms1x00.ins_pla_ands[12][12] ));
 sky130_fd_sc_hd__dfxtp_1 _10898_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_00703_),
    .Q(\tms1x00.ins_pla_ands[12][13] ));
 sky130_fd_sc_hd__dfxtp_2 _10899_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_00704_),
    .Q(\tms1x00.ins_pla_ands[12][14] ));
 sky130_fd_sc_hd__dfxtp_1 _10900_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_00705_),
    .Q(\tms1x00.ins_pla_ands[12][15] ));
 sky130_fd_sc_hd__dfxtp_1 _10901_ (.CLK(clknet_leaf_54_wb_clk_i),
    .D(_00706_),
    .Q(\tms1x00.ins_pla_ands[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _10902_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(_00707_),
    .Q(\tms1x00.ins_pla_ands[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _10903_ (.CLK(clknet_leaf_62_wb_clk_i),
    .D(_00708_),
    .Q(\tms1x00.ins_pla_ands[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _10904_ (.CLK(clknet_leaf_58_wb_clk_i),
    .D(_00709_),
    .Q(\tms1x00.ins_pla_ands[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _10905_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(_00710_),
    .Q(\tms1x00.ins_pla_ands[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _10906_ (.CLK(clknet_leaf_58_wb_clk_i),
    .D(_00711_),
    .Q(\tms1x00.ins_pla_ands[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _10907_ (.CLK(clknet_leaf_62_wb_clk_i),
    .D(_00712_),
    .Q(\tms1x00.ins_pla_ands[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _10908_ (.CLK(clknet_leaf_62_wb_clk_i),
    .D(_00713_),
    .Q(\tms1x00.ins_pla_ands[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _10909_ (.CLK(clknet_leaf_130_wb_clk_i),
    .D(_00714_),
    .Q(\tms1x00.ins_pla_ands[30][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10910_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_00715_),
    .Q(\tms1x00.ins_pla_ands[30][1] ));
 sky130_fd_sc_hd__dfxtp_1 _10911_ (.CLK(clknet_leaf_130_wb_clk_i),
    .D(_00716_),
    .Q(\tms1x00.ins_pla_ands[30][2] ));
 sky130_fd_sc_hd__dfxtp_1 _10912_ (.CLK(clknet_leaf_143_wb_clk_i),
    .D(_00717_),
    .Q(\tms1x00.ins_pla_ands[30][3] ));
 sky130_fd_sc_hd__dfxtp_1 _10913_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_00718_),
    .Q(\tms1x00.ins_pla_ands[30][4] ));
 sky130_fd_sc_hd__dfxtp_1 _10914_ (.CLK(clknet_leaf_138_wb_clk_i),
    .D(_00719_),
    .Q(\tms1x00.ins_pla_ands[30][5] ));
 sky130_fd_sc_hd__dfxtp_1 _10915_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_00720_),
    .Q(\tms1x00.ins_pla_ands[30][6] ));
 sky130_fd_sc_hd__dfxtp_1 _10916_ (.CLK(clknet_leaf_142_wb_clk_i),
    .D(_00721_),
    .Q(\tms1x00.ins_pla_ands[30][7] ));
 sky130_fd_sc_hd__dfxtp_1 _10917_ (.CLK(clknet_leaf_143_wb_clk_i),
    .D(_00722_),
    .Q(\tms1x00.ins_pla_ands[30][8] ));
 sky130_fd_sc_hd__dfxtp_1 _10918_ (.CLK(clknet_leaf_143_wb_clk_i),
    .D(_00723_),
    .Q(\tms1x00.ins_pla_ands[30][9] ));
 sky130_fd_sc_hd__dfxtp_1 _10919_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_00724_),
    .Q(\tms1x00.ins_pla_ands[30][10] ));
 sky130_fd_sc_hd__dfxtp_1 _10920_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_00725_),
    .Q(\tms1x00.ins_pla_ands[30][11] ));
 sky130_fd_sc_hd__dfxtp_1 _10921_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_00726_),
    .Q(\tms1x00.ins_pla_ands[30][12] ));
 sky130_fd_sc_hd__dfxtp_1 _10922_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_00727_),
    .Q(\tms1x00.ins_pla_ands[30][13] ));
 sky130_fd_sc_hd__dfxtp_1 _10923_ (.CLK(clknet_leaf_142_wb_clk_i),
    .D(_00728_),
    .Q(\tms1x00.ins_pla_ands[30][14] ));
 sky130_fd_sc_hd__dfxtp_1 _10924_ (.CLK(clknet_leaf_138_wb_clk_i),
    .D(_00729_),
    .Q(\tms1x00.ins_pla_ands[30][15] ));
 sky130_fd_sc_hd__dfxtp_1 _10925_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_00730_),
    .Q(\tms1x00.ins_pla_ands[20][4] ));
 sky130_fd_sc_hd__dfxtp_1 _10926_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_00731_),
    .Q(\tms1x00.ins_pla_ands[20][5] ));
 sky130_fd_sc_hd__dfxtp_1 _10927_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_00732_),
    .Q(\tms1x00.ins_pla_ands[20][6] ));
 sky130_fd_sc_hd__dfxtp_1 _10928_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_00733_),
    .Q(\tms1x00.ins_pla_ands[20][7] ));
 sky130_fd_sc_hd__dfxtp_1 _10929_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_00734_),
    .Q(\tms1x00.ins_pla_ands[20][8] ));
 sky130_fd_sc_hd__dfxtp_1 _10930_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_00735_),
    .Q(\tms1x00.ins_pla_ands[20][9] ));
 sky130_fd_sc_hd__dfxtp_1 _10931_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_00736_),
    .Q(\tms1x00.ins_pla_ands[20][12] ));
 sky130_fd_sc_hd__dfxtp_1 _10932_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_00737_),
    .Q(\tms1x00.ins_pla_ands[20][13] ));
 sky130_fd_sc_hd__dfxtp_1 _10933_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_00738_),
    .Q(\tms1x00.ins_pla_ands[20][14] ));
 sky130_fd_sc_hd__dfxtp_1 _10934_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_00739_),
    .Q(\tms1x00.ins_pla_ands[20][15] ));
 sky130_fd_sc_hd__dfxtp_1 _10935_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_00740_),
    .Q(\tms1x00.ins_pla_ands[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10936_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_00741_),
    .Q(\tms1x00.ins_pla_ands[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _10937_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_00742_),
    .Q(\tms1x00.ins_pla_ands[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _10938_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_00743_),
    .Q(\tms1x00.ins_pla_ands[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _10939_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_00744_),
    .Q(\tms1x00.ins_pla_ands[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 _10940_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_00745_),
    .Q(\tms1x00.ins_pla_ands[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 _10941_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_00746_),
    .Q(\tms1x00.ins_pla_ands[11][8] ));
 sky130_fd_sc_hd__dfxtp_1 _10942_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_00747_),
    .Q(\tms1x00.ins_pla_ands[11][9] ));
 sky130_fd_sc_hd__dfxtp_1 _10943_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_00748_),
    .Q(\tms1x00.ins_pla_ands[11][10] ));
 sky130_fd_sc_hd__dfxtp_1 _10944_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_00749_),
    .Q(\tms1x00.ins_pla_ands[11][11] ));
 sky130_fd_sc_hd__dfxtp_1 _10945_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_00750_),
    .Q(\tms1x00.ins_pla_ands[11][12] ));
 sky130_fd_sc_hd__dfxtp_1 _10946_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_00751_),
    .Q(\tms1x00.ins_pla_ands[11][13] ));
 sky130_fd_sc_hd__dfxtp_1 _10947_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_00752_),
    .Q(\tms1x00.ins_pla_ands[11][14] ));
 sky130_fd_sc_hd__dfxtp_1 _10948_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_00753_),
    .Q(\tms1x00.ins_pla_ands[11][15] ));
 sky130_fd_sc_hd__dfxtp_1 _10949_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(_00754_),
    .Q(\tms1x00.ins_pla_ands[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10950_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(_00755_),
    .Q(\tms1x00.ins_pla_ands[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _10951_ (.CLK(clknet_leaf_54_wb_clk_i),
    .D(_00756_),
    .Q(\tms1x00.ins_pla_ands[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _10952_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(_00757_),
    .Q(\tms1x00.ins_pla_ands[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _10953_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_00758_),
    .Q(\tms1x00.ins_pla_ands[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _10954_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_00759_),
    .Q(\tms1x00.ins_pla_ands[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _10955_ (.CLK(clknet_leaf_75_wb_clk_i),
    .D(_00760_),
    .Q(\tms1x00.O_pla_ors[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10956_ (.CLK(clknet_leaf_76_wb_clk_i),
    .D(_00761_),
    .Q(\tms1x00.O_pla_ors[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _10957_ (.CLK(clknet_leaf_61_wb_clk_i),
    .D(_00762_),
    .Q(\tms1x00.O_pla_ors[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _10958_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(_00763_),
    .Q(\tms1x00.O_pla_ors[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _10959_ (.CLK(clknet_leaf_61_wb_clk_i),
    .D(_00764_),
    .Q(\tms1x00.O_pla_ors[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _10960_ (.CLK(clknet_leaf_75_wb_clk_i),
    .D(_00765_),
    .Q(\tms1x00.O_pla_ors[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _10961_ (.CLK(clknet_leaf_79_wb_clk_i),
    .D(_00766_),
    .Q(\tms1x00.O_pla_ors[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _10962_ (.CLK(clknet_leaf_82_wb_clk_i),
    .D(_00767_),
    .Q(\tms1x00.O_pla_ors[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _10963_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(_00768_),
    .Q(\tms1x00.O_pla_ors[7][8] ));
 sky130_fd_sc_hd__dfxtp_1 _10964_ (.CLK(clknet_leaf_80_wb_clk_i),
    .D(_00769_),
    .Q(\tms1x00.O_pla_ors[7][9] ));
 sky130_fd_sc_hd__dfxtp_1 _10965_ (.CLK(clknet_leaf_80_wb_clk_i),
    .D(_00770_),
    .Q(\tms1x00.O_pla_ors[7][10] ));
 sky130_fd_sc_hd__dfxtp_1 _10966_ (.CLK(clknet_leaf_61_wb_clk_i),
    .D(_00771_),
    .Q(\tms1x00.O_pla_ors[7][11] ));
 sky130_fd_sc_hd__dfxtp_1 _10967_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(_00772_),
    .Q(\tms1x00.O_pla_ors[7][12] ));
 sky130_fd_sc_hd__dfxtp_1 _10968_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(_00773_),
    .Q(\tms1x00.O_pla_ors[7][13] ));
 sky130_fd_sc_hd__dfxtp_1 _10969_ (.CLK(clknet_leaf_82_wb_clk_i),
    .D(_00774_),
    .Q(\tms1x00.O_pla_ors[7][14] ));
 sky130_fd_sc_hd__dfxtp_1 _10970_ (.CLK(clknet_leaf_83_wb_clk_i),
    .D(_00775_),
    .Q(\tms1x00.O_pla_ors[7][15] ));
 sky130_fd_sc_hd__dfxtp_1 _10971_ (.CLK(clknet_leaf_82_wb_clk_i),
    .D(_00776_),
    .Q(\tms1x00.O_pla_ors[7][16] ));
 sky130_fd_sc_hd__dfxtp_1 _10972_ (.CLK(clknet_leaf_86_wb_clk_i),
    .D(_00777_),
    .Q(\tms1x00.O_pla_ors[7][17] ));
 sky130_fd_sc_hd__dfxtp_1 _10973_ (.CLK(clknet_leaf_75_wb_clk_i),
    .D(_00778_),
    .Q(\tms1x00.O_pla_ors[7][18] ));
 sky130_fd_sc_hd__dfxtp_1 _10974_ (.CLK(clknet_leaf_80_wb_clk_i),
    .D(_00779_),
    .Q(\tms1x00.O_pla_ors[7][19] ));
 sky130_fd_sc_hd__dfxtp_1 _10975_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_00780_),
    .Q(\tms1x00.ins_pla_ands[18][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10976_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_00781_),
    .Q(\tms1x00.ins_pla_ands[18][1] ));
 sky130_fd_sc_hd__dfxtp_1 _10977_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_00782_),
    .Q(\tms1x00.ins_pla_ands[18][2] ));
 sky130_fd_sc_hd__dfxtp_1 _10978_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_00783_),
    .Q(\tms1x00.ins_pla_ands[18][3] ));
 sky130_fd_sc_hd__dfxtp_1 _10979_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_00784_),
    .Q(\tms1x00.ins_pla_ands[18][4] ));
 sky130_fd_sc_hd__dfxtp_1 _10980_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_00785_),
    .Q(\tms1x00.ins_pla_ands[18][5] ));
 sky130_fd_sc_hd__dfxtp_1 _10981_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_00786_),
    .Q(\tms1x00.ins_pla_ands[18][6] ));
 sky130_fd_sc_hd__dfxtp_1 _10982_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_00787_),
    .Q(\tms1x00.ins_pla_ands[18][7] ));
 sky130_fd_sc_hd__dfxtp_1 _10983_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_00788_),
    .Q(\tms1x00.ins_pla_ands[18][10] ));
 sky130_fd_sc_hd__dfxtp_1 _10984_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_00789_),
    .Q(\tms1x00.ins_pla_ands[18][11] ));
 sky130_fd_sc_hd__dfxtp_1 _10985_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_00790_),
    .Q(\tms1x00.ins_pla_ands[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10986_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_00791_),
    .Q(\tms1x00.ins_pla_ands[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _10987_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_00792_),
    .Q(\tms1x00.ins_pla_ands[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _10988_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_00793_),
    .Q(\tms1x00.ins_pla_ands[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _10989_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_00794_),
    .Q(\tms1x00.ins_pla_ands[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 _10990_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_00795_),
    .Q(\tms1x00.ins_pla_ands[15][7] ));
 sky130_fd_sc_hd__dfxtp_1 _10991_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_00796_),
    .Q(\tms1x00.O_pla_ands[31][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10992_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_00797_),
    .Q(\tms1x00.O_pla_ands[31][1] ));
 sky130_fd_sc_hd__dfxtp_1 _10993_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_00798_),
    .Q(\tms1x00.O_pla_ands[31][2] ));
 sky130_fd_sc_hd__dfxtp_1 _10994_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_00799_),
    .Q(\tms1x00.O_pla_ands[31][3] ));
 sky130_fd_sc_hd__dfxtp_1 _10995_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_00800_),
    .Q(\tms1x00.O_pla_ands[31][4] ));
 sky130_fd_sc_hd__dfxtp_1 _10996_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_00801_),
    .Q(\tms1x00.O_pla_ands[31][5] ));
 sky130_fd_sc_hd__dfxtp_1 _10997_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_00802_),
    .Q(\tms1x00.O_pla_ands[31][6] ));
 sky130_fd_sc_hd__dfxtp_1 _10998_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_00803_),
    .Q(\tms1x00.O_pla_ands[31][7] ));
 sky130_fd_sc_hd__dfxtp_1 _10999_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_00804_),
    .Q(\tms1x00.O_pla_ands[31][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11000_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_00805_),
    .Q(\tms1x00.O_pla_ands[31][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11001_ (.CLK(clknet_leaf_54_wb_clk_i),
    .D(_00806_),
    .Q(\tms1x00.ins_pla_ands[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11002_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(_00807_),
    .Q(\tms1x00.ins_pla_ands[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11003_ (.CLK(clknet_leaf_54_wb_clk_i),
    .D(_00808_),
    .Q(\tms1x00.ins_pla_ands[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11004_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(_00809_),
    .Q(\tms1x00.ins_pla_ands[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11005_ (.CLK(clknet_leaf_54_wb_clk_i),
    .D(_00810_),
    .Q(\tms1x00.ins_pla_ands[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11006_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(_00811_),
    .Q(\tms1x00.ins_pla_ands[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11007_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(_00812_),
    .Q(\tms1x00.ins_pla_ands[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _11008_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(_00813_),
    .Q(\tms1x00.ins_pla_ands[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _11009_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(_00814_),
    .Q(\tms1x00.ins_pla_ands[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _11010_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(_00815_),
    .Q(\tms1x00.ins_pla_ands[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _11011_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_00816_),
    .Q(\tms1x00.ins_pla_ands[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11012_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_00817_),
    .Q(\tms1x00.ins_pla_ands[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11013_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_00818_),
    .Q(\tms1x00.ins_pla_ands[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11014_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_00819_),
    .Q(\tms1x00.ins_pla_ands[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11015_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_00820_),
    .Q(\tms1x00.ins_pla_ands[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11016_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_00821_),
    .Q(\tms1x00.ins_pla_ands[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11017_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_00822_),
    .Q(\tms1x00.ins_pla_ands[10][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11018_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_00823_),
    .Q(\tms1x00.ins_pla_ands[10][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11019_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_00824_),
    .Q(\tms1x00.ins_pla_ands[10][10] ));
 sky130_fd_sc_hd__dfxtp_1 _11020_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_00825_),
    .Q(\tms1x00.ins_pla_ands[10][11] ));
 sky130_fd_sc_hd__dfxtp_1 _11021_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_00826_),
    .Q(\tms1x00.ins_pla_ands[10][12] ));
 sky130_fd_sc_hd__dfxtp_1 _11022_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_00827_),
    .Q(\tms1x00.ins_pla_ands[10][13] ));
 sky130_fd_sc_hd__dfxtp_1 _11023_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_00828_),
    .Q(\tms1x00.ins_pla_ands[10][14] ));
 sky130_fd_sc_hd__dfxtp_1 _11024_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_00829_),
    .Q(\tms1x00.ins_pla_ands[10][15] ));
 sky130_fd_sc_hd__dfxtp_1 _11025_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(_00830_),
    .Q(\tms1x00.ins_pla_ands[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11026_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_00831_),
    .Q(\tms1x00.ins_pla_ands[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11027_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(_00832_),
    .Q(\tms1x00.ins_pla_ands[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11028_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(_00833_),
    .Q(\tms1x00.ins_pla_ands[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11029_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(_00834_),
    .Q(\tms1x00.ins_pla_ands[0][6] ));
 sky130_fd_sc_hd__dfxtp_2 _11030_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(_00835_),
    .Q(\tms1x00.ins_pla_ands[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11031_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_00836_),
    .Q(\tms1x00.ins_pla_ands[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _11032_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_00837_),
    .Q(\tms1x00.ins_pla_ands[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _11033_ (.CLK(clknet_leaf_77_wb_clk_i),
    .D(_00838_),
    .Q(\tms1x00.O_pla_ors[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11034_ (.CLK(clknet_leaf_76_wb_clk_i),
    .D(_00839_),
    .Q(\tms1x00.O_pla_ors[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11035_ (.CLK(clknet_leaf_61_wb_clk_i),
    .D(_00840_),
    .Q(\tms1x00.O_pla_ors[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11036_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(_00841_),
    .Q(\tms1x00.O_pla_ors[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11037_ (.CLK(clknet_leaf_60_wb_clk_i),
    .D(_00842_),
    .Q(\tms1x00.O_pla_ors[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11038_ (.CLK(clknet_leaf_75_wb_clk_i),
    .D(_00843_),
    .Q(\tms1x00.O_pla_ors[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11039_ (.CLK(clknet_leaf_79_wb_clk_i),
    .D(_00844_),
    .Q(\tms1x00.O_pla_ors[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11040_ (.CLK(clknet_leaf_84_wb_clk_i),
    .D(_00845_),
    .Q(\tms1x00.O_pla_ors[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11041_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(_00846_),
    .Q(\tms1x00.O_pla_ors[6][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11042_ (.CLK(clknet_leaf_79_wb_clk_i),
    .D(_00847_),
    .Q(\tms1x00.O_pla_ors[6][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11043_ (.CLK(clknet_leaf_82_wb_clk_i),
    .D(_00848_),
    .Q(\tms1x00.O_pla_ors[6][10] ));
 sky130_fd_sc_hd__dfxtp_1 _11044_ (.CLK(clknet_leaf_61_wb_clk_i),
    .D(_00849_),
    .Q(\tms1x00.O_pla_ors[6][11] ));
 sky130_fd_sc_hd__dfxtp_1 _11045_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(_00850_),
    .Q(\tms1x00.O_pla_ors[6][12] ));
 sky130_fd_sc_hd__dfxtp_1 _11046_ (.CLK(clknet_leaf_86_wb_clk_i),
    .D(_00851_),
    .Q(\tms1x00.O_pla_ors[6][13] ));
 sky130_fd_sc_hd__dfxtp_1 _11047_ (.CLK(clknet_leaf_83_wb_clk_i),
    .D(_00852_),
    .Q(\tms1x00.O_pla_ors[6][14] ));
 sky130_fd_sc_hd__dfxtp_1 _11048_ (.CLK(clknet_leaf_84_wb_clk_i),
    .D(_00853_),
    .Q(\tms1x00.O_pla_ors[6][15] ));
 sky130_fd_sc_hd__dfxtp_1 _11049_ (.CLK(clknet_leaf_82_wb_clk_i),
    .D(_00854_),
    .Q(\tms1x00.O_pla_ors[6][16] ));
 sky130_fd_sc_hd__dfxtp_1 _11050_ (.CLK(clknet_leaf_86_wb_clk_i),
    .D(_00855_),
    .Q(\tms1x00.O_pla_ors[6][17] ));
 sky130_fd_sc_hd__dfxtp_1 _11051_ (.CLK(clknet_leaf_75_wb_clk_i),
    .D(_00856_),
    .Q(\tms1x00.O_pla_ors[6][18] ));
 sky130_fd_sc_hd__dfxtp_1 _11052_ (.CLK(clknet_leaf_80_wb_clk_i),
    .D(_00857_),
    .Q(\tms1x00.O_pla_ors[6][19] ));
 sky130_fd_sc_hd__dfxtp_1 _11053_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_00858_),
    .Q(\tms1x00.ins_pla_ands[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11054_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_00859_),
    .Q(\tms1x00.ins_pla_ands[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11055_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_00860_),
    .Q(\tms1x00.ins_pla_ands[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11056_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_00861_),
    .Q(\tms1x00.ins_pla_ands[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11057_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_00862_),
    .Q(\tms1x00.ins_pla_ands[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11058_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_00863_),
    .Q(\tms1x00.ins_pla_ands[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11059_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_00864_),
    .Q(\tms1x00.ins_pla_ands[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11060_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_00865_),
    .Q(\tms1x00.ins_pla_ands[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11061_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(_00866_),
    .Q(\tms1x00.ins_pla_ands[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11062_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(_00867_),
    .Q(\tms1x00.ins_pla_ands[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11063_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(_00868_),
    .Q(\tms1x00.ins_pla_ands[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11064_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(_00869_),
    .Q(\tms1x00.ins_pla_ands[0][9] ));
 sky130_fd_sc_hd__dfxtp_2 _11065_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(_00870_),
    .Q(\tms1x00.ins_pla_ands[0][10] ));
 sky130_fd_sc_hd__dfxtp_2 _11066_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(_00871_),
    .Q(\tms1x00.ins_pla_ands[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _11067_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(_00872_),
    .Q(\tms1x00.ins_pla_ands[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _11068_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(_00873_),
    .Q(\tms1x00.ins_pla_ands[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _11069_ (.CLK(clknet_leaf_130_wb_clk_i),
    .D(_00874_),
    .Q(\tms1x00.ins_pla_ands[28][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11070_ (.CLK(clknet_leaf_140_wb_clk_i),
    .D(_00875_),
    .Q(\tms1x00.ins_pla_ands[28][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11071_ (.CLK(clknet_leaf_140_wb_clk_i),
    .D(_00876_),
    .Q(\tms1x00.ins_pla_ands[28][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11072_ (.CLK(clknet_leaf_140_wb_clk_i),
    .D(_00877_),
    .Q(\tms1x00.ins_pla_ands[28][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11073_ (.CLK(clknet_leaf_140_wb_clk_i),
    .D(_00878_),
    .Q(\tms1x00.ins_pla_ands[28][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11074_ (.CLK(clknet_leaf_140_wb_clk_i),
    .D(_00879_),
    .Q(\tms1x00.ins_pla_ands[28][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11075_ (.CLK(clknet_leaf_140_wb_clk_i),
    .D(_00880_),
    .Q(\tms1x00.ins_pla_ands[28][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11076_ (.CLK(clknet_leaf_141_wb_clk_i),
    .D(_00881_),
    .Q(\tms1x00.ins_pla_ands[28][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11077_ (.CLK(clknet_leaf_139_wb_clk_i),
    .D(_00882_),
    .Q(\tms1x00.ins_pla_ands[28][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11078_ (.CLK(clknet_leaf_130_wb_clk_i),
    .D(_00883_),
    .Q(\tms1x00.ins_pla_ands[28][11] ));
 sky130_fd_sc_hd__dfxtp_1 _11079_ (.CLK(clknet_leaf_142_wb_clk_i),
    .D(_00884_),
    .Q(\tms1x00.ins_pla_ands[28][12] ));
 sky130_fd_sc_hd__dfxtp_1 _11080_ (.CLK(clknet_leaf_142_wb_clk_i),
    .D(_00885_),
    .Q(\tms1x00.ins_pla_ands[28][15] ));
 sky130_fd_sc_hd__dfxtp_1 _11081_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_00886_),
    .Q(\tms1x00.ins_pla_ands[18][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11082_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_00887_),
    .Q(\tms1x00.ins_pla_ands[18][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11083_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_00888_),
    .Q(\tms1x00.ins_pla_ands[18][12] ));
 sky130_fd_sc_hd__dfxtp_1 _11084_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_00889_),
    .Q(\tms1x00.ins_pla_ands[18][13] ));
 sky130_fd_sc_hd__dfxtp_1 _11085_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_00890_),
    .Q(\tms1x00.ins_pla_ands[18][14] ));
 sky130_fd_sc_hd__dfxtp_1 _11086_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_00891_),
    .Q(\tms1x00.ins_pla_ands[18][15] ));
 sky130_fd_sc_hd__dfxtp_1 _11087_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_00892_),
    .Q(\tms1x00.ins_pla_ands[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11088_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_00893_),
    .Q(\tms1x00.ins_pla_ands[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11089_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_00894_),
    .Q(\tms1x00.ins_pla_ands[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11090_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_00895_),
    .Q(\tms1x00.ins_pla_ands[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11091_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(_00896_),
    .Q(\tms1x00.ins_pla_ands[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11092_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_00897_),
    .Q(\tms1x00.ins_pla_ands[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11093_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(_00898_),
    .Q(\tms1x00.ins_pla_ands[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11094_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_00899_),
    .Q(\tms1x00.ins_pla_ands[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11095_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_00900_),
    .Q(\tms1x00.ins_pla_ands[9][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11096_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_00901_),
    .Q(\tms1x00.ins_pla_ands[9][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11097_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(_00902_),
    .Q(\tms1x00.ins_pla_ands[9][10] ));
 sky130_fd_sc_hd__dfxtp_1 _11098_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_00903_),
    .Q(\tms1x00.ins_pla_ands[9][11] ));
 sky130_fd_sc_hd__dfxtp_1 _11099_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_00904_),
    .Q(\tms1x00.ins_pla_ands[9][12] ));
 sky130_fd_sc_hd__dfxtp_1 _11100_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(_00905_),
    .Q(\tms1x00.ins_pla_ands[9][13] ));
 sky130_fd_sc_hd__dfxtp_1 _11101_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(_00906_),
    .Q(\tms1x00.ins_pla_ands[9][14] ));
 sky130_fd_sc_hd__dfxtp_1 _11102_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(_00907_),
    .Q(\tms1x00.ins_pla_ands[9][15] ));
 sky130_fd_sc_hd__dfxtp_1 _11103_ (.CLK(clknet_leaf_74_wb_clk_i),
    .D(_00908_),
    .Q(\tms1x00.O_pla_ors[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11104_ (.CLK(clknet_leaf_76_wb_clk_i),
    .D(_00909_),
    .Q(\tms1x00.O_pla_ors[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11105_ (.CLK(clknet_leaf_69_wb_clk_i),
    .D(_00910_),
    .Q(\tms1x00.O_pla_ors[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11106_ (.CLK(clknet_leaf_70_wb_clk_i),
    .D(_00911_),
    .Q(\tms1x00.O_pla_ors[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11107_ (.CLK(clknet_leaf_85_wb_clk_i),
    .D(_00912_),
    .Q(\tms1x00.O_pla_ors[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11108_ (.CLK(clknet_leaf_75_wb_clk_i),
    .D(_00913_),
    .Q(\tms1x00.O_pla_ors[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11109_ (.CLK(clknet_leaf_79_wb_clk_i),
    .D(_00914_),
    .Q(\tms1x00.O_pla_ors[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11110_ (.CLK(clknet_leaf_84_wb_clk_i),
    .D(_00915_),
    .Q(\tms1x00.O_pla_ors[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11111_ (.CLK(clknet_leaf_69_wb_clk_i),
    .D(_00916_),
    .Q(\tms1x00.O_pla_ors[5][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11112_ (.CLK(clknet_leaf_79_wb_clk_i),
    .D(_00917_),
    .Q(\tms1x00.O_pla_ors[5][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11113_ (.CLK(clknet_leaf_80_wb_clk_i),
    .D(_00918_),
    .Q(\tms1x00.O_pla_ors[5][10] ));
 sky130_fd_sc_hd__dfxtp_1 _11114_ (.CLK(clknet_leaf_69_wb_clk_i),
    .D(_00919_),
    .Q(\tms1x00.O_pla_ors[5][11] ));
 sky130_fd_sc_hd__dfxtp_1 _11115_ (.CLK(clknet_leaf_85_wb_clk_i),
    .D(_00920_),
    .Q(\tms1x00.O_pla_ors[5][12] ));
 sky130_fd_sc_hd__dfxtp_1 _11116_ (.CLK(clknet_leaf_85_wb_clk_i),
    .D(_00921_),
    .Q(\tms1x00.O_pla_ors[5][13] ));
 sky130_fd_sc_hd__dfxtp_1 _11117_ (.CLK(clknet_leaf_84_wb_clk_i),
    .D(_00922_),
    .Q(\tms1x00.O_pla_ors[5][14] ));
 sky130_fd_sc_hd__dfxtp_1 _11118_ (.CLK(clknet_leaf_84_wb_clk_i),
    .D(_00923_),
    .Q(\tms1x00.O_pla_ors[5][15] ));
 sky130_fd_sc_hd__dfxtp_1 _11119_ (.CLK(clknet_leaf_80_wb_clk_i),
    .D(_00924_),
    .Q(\tms1x00.O_pla_ors[5][16] ));
 sky130_fd_sc_hd__dfxtp_1 _11120_ (.CLK(clknet_leaf_86_wb_clk_i),
    .D(_00925_),
    .Q(\tms1x00.O_pla_ors[5][17] ));
 sky130_fd_sc_hd__dfxtp_1 _11121_ (.CLK(clknet_leaf_75_wb_clk_i),
    .D(_00926_),
    .Q(\tms1x00.O_pla_ors[5][18] ));
 sky130_fd_sc_hd__dfxtp_1 _11122_ (.CLK(clknet_leaf_80_wb_clk_i),
    .D(_00927_),
    .Q(\tms1x00.O_pla_ors[5][19] ));
 sky130_fd_sc_hd__dfxtp_1 _11123_ (.CLK(clknet_leaf_130_wb_clk_i),
    .D(_00928_),
    .Q(\tms1x00.ins_pla_ands[27][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11124_ (.CLK(clknet_leaf_130_wb_clk_i),
    .D(_00929_),
    .Q(\tms1x00.ins_pla_ands[27][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11125_ (.CLK(clknet_leaf_140_wb_clk_i),
    .D(_00930_),
    .Q(\tms1x00.ins_pla_ands[27][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11126_ (.CLK(clknet_leaf_141_wb_clk_i),
    .D(_00931_),
    .Q(\tms1x00.ins_pla_ands[27][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11127_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_00932_),
    .Q(\tms1x00.ins_pla_ands[27][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11128_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_00933_),
    .Q(\tms1x00.ins_pla_ands[27][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11129_ (.CLK(clknet_leaf_141_wb_clk_i),
    .D(_00934_),
    .Q(\tms1x00.ins_pla_ands[27][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11130_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_00935_),
    .Q(\tms1x00.ins_pla_ands[27][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11131_ (.CLK(clknet_leaf_138_wb_clk_i),
    .D(_00936_),
    .Q(\tms1x00.ins_pla_ands[27][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11132_ (.CLK(clknet_leaf_140_wb_clk_i),
    .D(_00937_),
    .Q(\tms1x00.ins_pla_ands[27][10] ));
 sky130_fd_sc_hd__dfxtp_1 _11133_ (.CLK(clknet_leaf_136_wb_clk_i),
    .D(_00938_),
    .Q(\tms1x00.ins_pla_ands[27][12] ));
 sky130_fd_sc_hd__dfxtp_1 _11134_ (.CLK(clknet_leaf_141_wb_clk_i),
    .D(_00939_),
    .Q(\tms1x00.ins_pla_ands[27][15] ));
 sky130_fd_sc_hd__dfxtp_1 _11135_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_00940_),
    .Q(\tms1x00.ins_pla_ands[17][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11136_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_00941_),
    .Q(\tms1x00.ins_pla_ands[17][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11137_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_00942_),
    .Q(\tms1x00.ins_pla_ands[17][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11138_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_00943_),
    .Q(\tms1x00.ins_pla_ands[17][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11139_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_00944_),
    .Q(\tms1x00.ins_pla_ands[17][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11140_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_00945_),
    .Q(\tms1x00.ins_pla_ands[17][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11141_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_00946_),
    .Q(\tms1x00.ins_pla_ands[17][12] ));
 sky130_fd_sc_hd__dfxtp_1 _11142_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_00947_),
    .Q(\tms1x00.ins_pla_ands[17][13] ));
 sky130_fd_sc_hd__dfxtp_1 _11143_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_00948_),
    .Q(\tms1x00.ins_pla_ands[17][14] ));
 sky130_fd_sc_hd__dfxtp_1 _11144_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_00949_),
    .Q(\tms1x00.ins_pla_ands[17][15] ));
 sky130_fd_sc_hd__dfxtp_1 _11145_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_00950_),
    .Q(\tms1x00.ins_pla_ands[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11146_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_00951_),
    .Q(\tms1x00.ins_pla_ands[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11147_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_00952_),
    .Q(\tms1x00.ins_pla_ands[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11148_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_00953_),
    .Q(\tms1x00.ins_pla_ands[8][12] ));
 sky130_fd_sc_hd__dfxtp_1 _11149_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_00954_),
    .Q(\tms1x00.ins_pla_ands[8][13] ));
 sky130_fd_sc_hd__dfxtp_1 _11150_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_00955_),
    .Q(\tms1x00.ins_pla_ands[8][14] ));
 sky130_fd_sc_hd__dfxtp_1 _11151_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_00956_),
    .Q(\tms1x00.ins_pla_ands[8][15] ));
 sky130_fd_sc_hd__dfxtp_1 _11152_ (.CLK(clknet_leaf_77_wb_clk_i),
    .D(_00957_),
    .Q(\tms1x00.O_pla_ors[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11153_ (.CLK(clknet_leaf_76_wb_clk_i),
    .D(_00958_),
    .Q(\tms1x00.O_pla_ors[4][1] ));
 sky130_fd_sc_hd__dfxtp_2 _11154_ (.CLK(clknet_leaf_62_wb_clk_i),
    .D(_00959_),
    .Q(\tms1x00.O_pla_ors[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11155_ (.CLK(clknet_leaf_85_wb_clk_i),
    .D(_00960_),
    .Q(\tms1x00.O_pla_ors[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11156_ (.CLK(clknet_leaf_60_wb_clk_i),
    .D(_00961_),
    .Q(\tms1x00.O_pla_ors[4][4] ));
 sky130_fd_sc_hd__dfxtp_2 _11157_ (.CLK(clknet_leaf_60_wb_clk_i),
    .D(_00962_),
    .Q(\tms1x00.O_pla_ors[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11158_ (.CLK(clknet_leaf_78_wb_clk_i),
    .D(_00963_),
    .Q(\tms1x00.O_pla_ors[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11159_ (.CLK(clknet_leaf_84_wb_clk_i),
    .D(_00964_),
    .Q(\tms1x00.O_pla_ors[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11160_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(_00965_),
    .Q(\tms1x00.O_pla_ors[4][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11161_ (.CLK(clknet_leaf_78_wb_clk_i),
    .D(_00966_),
    .Q(\tms1x00.O_pla_ors[4][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11162_ (.CLK(clknet_leaf_78_wb_clk_i),
    .D(_00967_),
    .Q(\tms1x00.O_pla_ors[4][10] ));
 sky130_fd_sc_hd__dfxtp_2 _11163_ (.CLK(clknet_leaf_61_wb_clk_i),
    .D(_00968_),
    .Q(\tms1x00.O_pla_ors[4][11] ));
 sky130_fd_sc_hd__dfxtp_1 _11164_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(_00969_),
    .Q(\tms1x00.O_pla_ors[4][12] ));
 sky130_fd_sc_hd__dfxtp_1 _11165_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(_00970_),
    .Q(\tms1x00.O_pla_ors[4][13] ));
 sky130_fd_sc_hd__dfxtp_1 _11166_ (.CLK(clknet_leaf_84_wb_clk_i),
    .D(_00971_),
    .Q(\tms1x00.O_pla_ors[4][14] ));
 sky130_fd_sc_hd__dfxtp_1 _11167_ (.CLK(clknet_leaf_84_wb_clk_i),
    .D(_00972_),
    .Q(\tms1x00.O_pla_ors[4][15] ));
 sky130_fd_sc_hd__dfxtp_1 _11168_ (.CLK(clknet_leaf_80_wb_clk_i),
    .D(_00973_),
    .Q(\tms1x00.O_pla_ors[4][16] ));
 sky130_fd_sc_hd__dfxtp_1 _11169_ (.CLK(clknet_leaf_86_wb_clk_i),
    .D(_00974_),
    .Q(\tms1x00.O_pla_ors[4][17] ));
 sky130_fd_sc_hd__dfxtp_1 _11170_ (.CLK(clknet_leaf_77_wb_clk_i),
    .D(_00975_),
    .Q(\tms1x00.O_pla_ors[4][18] ));
 sky130_fd_sc_hd__dfxtp_2 _11171_ (.CLK(clknet_leaf_86_wb_clk_i),
    .D(_00976_),
    .Q(\tms1x00.O_pla_ors[4][19] ));
 sky130_fd_sc_hd__dfxtp_1 _11172_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_00977_),
    .Q(\tms1x00.ins_pla_ands[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11173_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_00978_),
    .Q(\tms1x00.ins_pla_ands[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11174_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_00979_),
    .Q(\tms1x00.ins_pla_ands[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11175_ (.CLK(clknet_leaf_130_wb_clk_i),
    .D(_00980_),
    .Q(\tms1x00.ins_pla_ands[26][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11176_ (.CLK(clknet_leaf_140_wb_clk_i),
    .D(_00981_),
    .Q(\tms1x00.ins_pla_ands[26][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11177_ (.CLK(clknet_leaf_140_wb_clk_i),
    .D(_00982_),
    .Q(\tms1x00.ins_pla_ands[26][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11178_ (.CLK(clknet_leaf_141_wb_clk_i),
    .D(_00983_),
    .Q(\tms1x00.ins_pla_ands[26][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11179_ (.CLK(clknet_leaf_141_wb_clk_i),
    .D(_00984_),
    .Q(\tms1x00.ins_pla_ands[26][14] ));
 sky130_fd_sc_hd__dfxtp_1 _11180_ (.CLK(clknet_leaf_141_wb_clk_i),
    .D(_00985_),
    .Q(\tms1x00.ins_pla_ands[26][15] ));
 sky130_fd_sc_hd__dfxtp_1 _11181_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_00986_),
    .Q(\tms1x00.ins_pla_ands[16][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11182_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_00987_),
    .Q(\tms1x00.ins_pla_ands[16][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11183_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_00988_),
    .Q(\tms1x00.ins_pla_ands[16][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11184_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_00989_),
    .Q(\tms1x00.ins_pla_ands[16][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11185_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(_00990_),
    .Q(\tms1x00.ins_pla_ands[7][12] ));
 sky130_fd_sc_hd__dfxtp_1 _11186_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(_00991_),
    .Q(\tms1x00.ins_pla_ands[7][13] ));
 sky130_fd_sc_hd__dfxtp_1 _11187_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_00992_),
    .Q(\tms1x00.ins_pla_ands[7][14] ));
 sky130_fd_sc_hd__dfxtp_1 _11188_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_00993_),
    .Q(\tms1x00.ins_pla_ands[7][15] ));
 sky130_fd_sc_hd__dfxtp_1 _11189_ (.CLK(clknet_leaf_77_wb_clk_i),
    .D(_00994_),
    .Q(\tms1x00.O_pla_ors[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11190_ (.CLK(clknet_leaf_77_wb_clk_i),
    .D(_00995_),
    .Q(\tms1x00.O_pla_ors[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11191_ (.CLK(clknet_leaf_60_wb_clk_i),
    .D(_00996_),
    .Q(\tms1x00.O_pla_ors[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11192_ (.CLK(clknet_leaf_60_wb_clk_i),
    .D(_00997_),
    .Q(\tms1x00.O_pla_ors[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11193_ (.CLK(clknet_leaf_60_wb_clk_i),
    .D(_00998_),
    .Q(\tms1x00.O_pla_ors[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11194_ (.CLK(clknet_leaf_77_wb_clk_i),
    .D(_00999_),
    .Q(\tms1x00.O_pla_ors[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11195_ (.CLK(clknet_leaf_79_wb_clk_i),
    .D(_01000_),
    .Q(\tms1x00.O_pla_ors[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11196_ (.CLK(clknet_leaf_84_wb_clk_i),
    .D(_01001_),
    .Q(\tms1x00.O_pla_ors[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11197_ (.CLK(clknet_leaf_60_wb_clk_i),
    .D(_01002_),
    .Q(\tms1x00.O_pla_ors[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11198_ (.CLK(clknet_leaf_79_wb_clk_i),
    .D(_01003_),
    .Q(\tms1x00.O_pla_ors[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11199_ (.CLK(clknet_leaf_79_wb_clk_i),
    .D(_01004_),
    .Q(\tms1x00.O_pla_ors[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _11200_ (.CLK(clknet_leaf_61_wb_clk_i),
    .D(_01005_),
    .Q(\tms1x00.O_pla_ors[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _11201_ (.CLK(clknet_leaf_60_wb_clk_i),
    .D(_01006_),
    .Q(\tms1x00.O_pla_ors[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _11202_ (.CLK(clknet_leaf_86_wb_clk_i),
    .D(_01007_),
    .Q(\tms1x00.O_pla_ors[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _11203_ (.CLK(clknet_leaf_84_wb_clk_i),
    .D(_01008_),
    .Q(\tms1x00.O_pla_ors[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _11204_ (.CLK(clknet_leaf_84_wb_clk_i),
    .D(_01009_),
    .Q(\tms1x00.O_pla_ors[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _11205_ (.CLK(clknet_leaf_84_wb_clk_i),
    .D(_01010_),
    .Q(\tms1x00.O_pla_ors[3][16] ));
 sky130_fd_sc_hd__dfxtp_1 _11206_ (.CLK(clknet_leaf_86_wb_clk_i),
    .D(_01011_),
    .Q(\tms1x00.O_pla_ors[3][17] ));
 sky130_fd_sc_hd__dfxtp_1 _11207_ (.CLK(clknet_leaf_77_wb_clk_i),
    .D(_01012_),
    .Q(\tms1x00.O_pla_ors[3][18] ));
 sky130_fd_sc_hd__dfxtp_1 _11208_ (.CLK(clknet_leaf_79_wb_clk_i),
    .D(_01013_),
    .Q(\tms1x00.O_pla_ors[3][19] ));
 sky130_fd_sc_hd__dfxtp_1 _11209_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_01014_),
    .Q(\tms1x00.ins_pla_ands[25][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11210_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_01015_),
    .Q(\tms1x00.ins_pla_ands[25][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11211_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_01016_),
    .Q(\tms1x00.ins_pla_ands[25][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11212_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_01017_),
    .Q(\tms1x00.ins_pla_ands[25][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11213_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_01018_),
    .Q(\tms1x00.ins_pla_ands[25][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11214_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_01019_),
    .Q(\tms1x00.ins_pla_ands[25][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11215_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_01020_),
    .Q(\tms1x00.ins_pla_ands[25][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11216_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_01021_),
    .Q(\tms1x00.ins_pla_ands[25][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11217_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_01022_),
    .Q(\tms1x00.ins_pla_ands[25][12] ));
 sky130_fd_sc_hd__dfxtp_1 _11218_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_01023_),
    .Q(\tms1x00.ins_pla_ands[25][13] ));
 sky130_fd_sc_hd__dfxtp_2 _11219_ (.CLK(clknet_leaf_143_wb_clk_i),
    .D(_01024_),
    .Q(\tms1x00.ins_pla_ands[25][14] ));
 sky130_fd_sc_hd__dfxtp_1 _11220_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_01025_),
    .Q(\tms1x00.ins_pla_ands[25][15] ));
 sky130_fd_sc_hd__dfxtp_1 _11221_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_01026_),
    .Q(\tms1x00.ins_pla_ands[16][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11222_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_01027_),
    .Q(\tms1x00.ins_pla_ands[16][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11223_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_01028_),
    .Q(\tms1x00.ins_pla_ands[16][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11224_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_01029_),
    .Q(\tms1x00.ins_pla_ands[16][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11225_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_01030_),
    .Q(\tms1x00.ins_pla_ands[16][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11226_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_01031_),
    .Q(\tms1x00.ins_pla_ands[16][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11227_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_01032_),
    .Q(\tms1x00.ins_pla_ands[16][10] ));
 sky130_fd_sc_hd__dfxtp_1 _11228_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_01033_),
    .Q(\tms1x00.ins_pla_ands[16][11] ));
 sky130_fd_sc_hd__dfxtp_1 _11229_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_01034_),
    .Q(\tms1x00.ins_pla_ands[16][12] ));
 sky130_fd_sc_hd__dfxtp_1 _11230_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_01035_),
    .Q(\tms1x00.ins_pla_ands[16][13] ));
 sky130_fd_sc_hd__dfxtp_1 _11231_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_01036_),
    .Q(\tms1x00.ins_pla_ands[16][14] ));
 sky130_fd_sc_hd__dfxtp_1 _11232_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_01037_),
    .Q(\tms1x00.ins_pla_ands[16][15] ));
 sky130_fd_sc_hd__dfxtp_1 _11233_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_01038_),
    .Q(\tms1x00.ins_pla_ands[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11234_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(_01039_),
    .Q(\tms1x00.ins_pla_ands[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11235_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(_01040_),
    .Q(\tms1x00.ins_pla_ands[6][12] ));
 sky130_fd_sc_hd__dfxtp_1 _11236_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(_01041_),
    .Q(\tms1x00.ins_pla_ands[6][13] ));
 sky130_fd_sc_hd__dfxtp_1 _11237_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(_01042_),
    .Q(\tms1x00.ins_pla_ands[6][14] ));
 sky130_fd_sc_hd__dfxtp_1 _11238_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_01043_),
    .Q(\tms1x00.ins_pla_ands[6][15] ));
 sky130_fd_sc_hd__dfxtp_1 _11239_ (.CLK(clknet_leaf_74_wb_clk_i),
    .D(_01044_),
    .Q(\tms1x00.O_pla_ors[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11240_ (.CLK(clknet_leaf_76_wb_clk_i),
    .D(_01045_),
    .Q(\tms1x00.O_pla_ors[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11241_ (.CLK(clknet_leaf_61_wb_clk_i),
    .D(_01046_),
    .Q(\tms1x00.O_pla_ors[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11242_ (.CLK(clknet_leaf_85_wb_clk_i),
    .D(_01047_),
    .Q(\tms1x00.O_pla_ors[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11243_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(_01048_),
    .Q(\tms1x00.O_pla_ors[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11244_ (.CLK(clknet_leaf_75_wb_clk_i),
    .D(_01049_),
    .Q(\tms1x00.O_pla_ors[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11245_ (.CLK(clknet_leaf_79_wb_clk_i),
    .D(_01050_),
    .Q(\tms1x00.O_pla_ors[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11246_ (.CLK(clknet_leaf_82_wb_clk_i),
    .D(_01051_),
    .Q(\tms1x00.O_pla_ors[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11247_ (.CLK(clknet_leaf_60_wb_clk_i),
    .D(_01052_),
    .Q(\tms1x00.O_pla_ors[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11248_ (.CLK(clknet_leaf_79_wb_clk_i),
    .D(_01053_),
    .Q(\tms1x00.O_pla_ors[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11249_ (.CLK(clknet_leaf_80_wb_clk_i),
    .D(_01054_),
    .Q(\tms1x00.O_pla_ors[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _11250_ (.CLK(clknet_leaf_69_wb_clk_i),
    .D(_01055_),
    .Q(\tms1x00.O_pla_ors[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _11251_ (.CLK(clknet_leaf_60_wb_clk_i),
    .D(_01056_),
    .Q(\tms1x00.O_pla_ors[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _11252_ (.CLK(clknet_leaf_86_wb_clk_i),
    .D(_01057_),
    .Q(\tms1x00.O_pla_ors[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _11253_ (.CLK(clknet_leaf_84_wb_clk_i),
    .D(_01058_),
    .Q(\tms1x00.O_pla_ors[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _11254_ (.CLK(clknet_leaf_84_wb_clk_i),
    .D(_01059_),
    .Q(\tms1x00.O_pla_ors[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _11255_ (.CLK(clknet_leaf_80_wb_clk_i),
    .D(_01060_),
    .Q(\tms1x00.O_pla_ors[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _11256_ (.CLK(clknet_leaf_86_wb_clk_i),
    .D(_01061_),
    .Q(\tms1x00.O_pla_ors[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _11257_ (.CLK(clknet_leaf_75_wb_clk_i),
    .D(_01062_),
    .Q(\tms1x00.O_pla_ors[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _11258_ (.CLK(clknet_leaf_80_wb_clk_i),
    .D(_01063_),
    .Q(\tms1x00.O_pla_ors[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _11259_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_01064_),
    .Q(\tms1x00.ins_pla_ands[24][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11260_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_01065_),
    .Q(\tms1x00.ins_pla_ands[24][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11261_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_01066_),
    .Q(\tms1x00.ins_pla_ands[24][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11262_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_01067_),
    .Q(\tms1x00.ins_pla_ands[24][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11263_ (.CLK(clknet_leaf_141_wb_clk_i),
    .D(_01068_),
    .Q(\tms1x00.ins_pla_ands[24][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11264_ (.CLK(clknet_leaf_141_wb_clk_i),
    .D(_01069_),
    .Q(\tms1x00.ins_pla_ands[24][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11265_ (.CLK(clknet_leaf_143_wb_clk_i),
    .D(_01070_),
    .Q(\tms1x00.ins_pla_ands[24][12] ));
 sky130_fd_sc_hd__dfxtp_1 _11266_ (.CLK(clknet_leaf_141_wb_clk_i),
    .D(_01071_),
    .Q(\tms1x00.ins_pla_ands[24][13] ));
 sky130_fd_sc_hd__dfxtp_1 _11267_ (.CLK(clknet_leaf_143_wb_clk_i),
    .D(_01072_),
    .Q(\tms1x00.ins_pla_ands[24][14] ));
 sky130_fd_sc_hd__dfxtp_1 _11268_ (.CLK(clknet_leaf_141_wb_clk_i),
    .D(_01073_),
    .Q(\tms1x00.ins_pla_ands[24][15] ));
 sky130_fd_sc_hd__dfxtp_1 _11269_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_01074_),
    .Q(\tms1x00.ins_pla_ands[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11270_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_01075_),
    .Q(\tms1x00.ins_pla_ands[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11271_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_01076_),
    .Q(\tms1x00.ins_pla_ands[15][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11272_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_01077_),
    .Q(\tms1x00.ins_pla_ands[15][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11273_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_01078_),
    .Q(\tms1x00.ins_pla_ands[15][10] ));
 sky130_fd_sc_hd__dfxtp_1 _11274_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_01079_),
    .Q(\tms1x00.ins_pla_ands[15][11] ));
 sky130_fd_sc_hd__dfxtp_1 _11275_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_01080_),
    .Q(\tms1x00.ins_pla_ands[15][12] ));
 sky130_fd_sc_hd__dfxtp_1 _11276_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_01081_),
    .Q(\tms1x00.ins_pla_ands[15][13] ));
 sky130_fd_sc_hd__dfxtp_1 _11277_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_01082_),
    .Q(\tms1x00.ins_pla_ands[15][14] ));
 sky130_fd_sc_hd__dfxtp_1 _11278_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_01083_),
    .Q(\tms1x00.ins_pla_ands[15][15] ));
 sky130_fd_sc_hd__dfxtp_1 _11279_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(_01084_),
    .Q(\tms1x00.ins_pla_ands[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11280_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(_01085_),
    .Q(\tms1x00.ins_pla_ands[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11281_ (.CLK(clknet_leaf_58_wb_clk_i),
    .D(_01086_),
    .Q(\tms1x00.ins_pla_ands[5][12] ));
 sky130_fd_sc_hd__dfxtp_1 _11282_ (.CLK(clknet_leaf_58_wb_clk_i),
    .D(_01087_),
    .Q(\tms1x00.ins_pla_ands[5][13] ));
 sky130_fd_sc_hd__dfxtp_1 _11283_ (.CLK(clknet_leaf_62_wb_clk_i),
    .D(_01088_),
    .Q(\tms1x00.ins_pla_ands[5][14] ));
 sky130_fd_sc_hd__dfxtp_1 _11284_ (.CLK(clknet_leaf_58_wb_clk_i),
    .D(_01089_),
    .Q(\tms1x00.ins_pla_ands[5][15] ));
 sky130_fd_sc_hd__dfxtp_1 _11285_ (.CLK(clknet_leaf_74_wb_clk_i),
    .D(_01090_),
    .Q(\tms1x00.O_pla_ors[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11286_ (.CLK(clknet_leaf_76_wb_clk_i),
    .D(_01091_),
    .Q(\tms1x00.O_pla_ors[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11287_ (.CLK(clknet_leaf_70_wb_clk_i),
    .D(_01092_),
    .Q(\tms1x00.O_pla_ors[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11288_ (.CLK(clknet_leaf_77_wb_clk_i),
    .D(_01093_),
    .Q(\tms1x00.O_pla_ors[1][3] ));
 sky130_fd_sc_hd__dfxtp_2 _11289_ (.CLK(clknet_leaf_77_wb_clk_i),
    .D(_01094_),
    .Q(\tms1x00.O_pla_ors[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11290_ (.CLK(clknet_leaf_75_wb_clk_i),
    .D(_01095_),
    .Q(\tms1x00.O_pla_ors[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11291_ (.CLK(clknet_leaf_75_wb_clk_i),
    .D(_01096_),
    .Q(\tms1x00.O_pla_ors[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11292_ (.CLK(clknet_leaf_78_wb_clk_i),
    .D(_01097_),
    .Q(\tms1x00.O_pla_ors[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11293_ (.CLK(clknet_leaf_77_wb_clk_i),
    .D(_01098_),
    .Q(\tms1x00.O_pla_ors[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11294_ (.CLK(clknet_leaf_79_wb_clk_i),
    .D(_01099_),
    .Q(\tms1x00.O_pla_ors[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11295_ (.CLK(clknet_leaf_77_wb_clk_i),
    .D(_01100_),
    .Q(\tms1x00.O_pla_ors[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _11296_ (.CLK(clknet_leaf_77_wb_clk_i),
    .D(_01101_),
    .Q(\tms1x00.O_pla_ors[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _11297_ (.CLK(clknet_leaf_77_wb_clk_i),
    .D(_01102_),
    .Q(\tms1x00.O_pla_ors[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _11298_ (.CLK(clknet_leaf_85_wb_clk_i),
    .D(_01103_),
    .Q(\tms1x00.O_pla_ors[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _11299_ (.CLK(clknet_leaf_78_wb_clk_i),
    .D(_01104_),
    .Q(\tms1x00.O_pla_ors[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _11300_ (.CLK(clknet_leaf_77_wb_clk_i),
    .D(_01105_),
    .Q(\tms1x00.O_pla_ors[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _11301_ (.CLK(clknet_leaf_78_wb_clk_i),
    .D(_01106_),
    .Q(\tms1x00.O_pla_ors[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _11302_ (.CLK(clknet_leaf_85_wb_clk_i),
    .D(_01107_),
    .Q(\tms1x00.O_pla_ors[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _11303_ (.CLK(clknet_leaf_76_wb_clk_i),
    .D(_01108_),
    .Q(\tms1x00.O_pla_ors[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _11304_ (.CLK(clknet_leaf_78_wb_clk_i),
    .D(_01109_),
    .Q(\tms1x00.O_pla_ors[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _11305_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_01110_),
    .Q(\tms1x00.ins_pla_ands[17][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11306_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_01111_),
    .Q(\tms1x00.ins_pla_ands[17][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11307_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_01112_),
    .Q(\tms1x00.ins_pla_ands[17][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11308_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_01113_),
    .Q(\tms1x00.ins_pla_ands[17][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11309_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_01114_),
    .Q(\tms1x00.ins_pla_ands[17][10] ));
 sky130_fd_sc_hd__dfxtp_1 _11310_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_01115_),
    .Q(\tms1x00.ins_pla_ands[17][11] ));
 sky130_fd_sc_hd__dfxtp_1 _11311_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_01116_),
    .Q(\tms1x00.ins_pla_ands[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11312_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_01117_),
    .Q(\tms1x00.ins_pla_ands[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11313_ (.CLK(clknet_leaf_74_wb_clk_i),
    .D(_01118_),
    .Q(\tms1x00.O_pla_ors[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11314_ (.CLK(clknet_leaf_76_wb_clk_i),
    .D(_01119_),
    .Q(\tms1x00.O_pla_ors[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11315_ (.CLK(clknet_leaf_70_wb_clk_i),
    .D(_01120_),
    .Q(\tms1x00.O_pla_ors[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11316_ (.CLK(clknet_leaf_70_wb_clk_i),
    .D(_01121_),
    .Q(\tms1x00.O_pla_ors[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11317_ (.CLK(clknet_leaf_85_wb_clk_i),
    .D(_01122_),
    .Q(\tms1x00.O_pla_ors[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11318_ (.CLK(clknet_leaf_74_wb_clk_i),
    .D(_01123_),
    .Q(\tms1x00.O_pla_ors[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11319_ (.CLK(clknet_leaf_79_wb_clk_i),
    .D(_01124_),
    .Q(\tms1x00.O_pla_ors[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11320_ (.CLK(clknet_leaf_85_wb_clk_i),
    .D(_01125_),
    .Q(\tms1x00.O_pla_ors[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11321_ (.CLK(clknet_leaf_76_wb_clk_i),
    .D(_01126_),
    .Q(\tms1x00.O_pla_ors[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11322_ (.CLK(clknet_leaf_78_wb_clk_i),
    .D(_01127_),
    .Q(\tms1x00.O_pla_ors[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11323_ (.CLK(clknet_leaf_78_wb_clk_i),
    .D(_01128_),
    .Q(\tms1x00.O_pla_ors[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _11324_ (.CLK(clknet_leaf_70_wb_clk_i),
    .D(_01129_),
    .Q(\tms1x00.O_pla_ors[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _11325_ (.CLK(clknet_leaf_77_wb_clk_i),
    .D(_01130_),
    .Q(\tms1x00.O_pla_ors[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _11326_ (.CLK(clknet_leaf_85_wb_clk_i),
    .D(_01131_),
    .Q(\tms1x00.O_pla_ors[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _11327_ (.CLK(clknet_leaf_84_wb_clk_i),
    .D(_01132_),
    .Q(\tms1x00.O_pla_ors[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _11328_ (.CLK(clknet_leaf_85_wb_clk_i),
    .D(_01133_),
    .Q(\tms1x00.O_pla_ors[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _11329_ (.CLK(clknet_leaf_84_wb_clk_i),
    .D(_01134_),
    .Q(\tms1x00.O_pla_ors[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _11330_ (.CLK(clknet_leaf_85_wb_clk_i),
    .D(_01135_),
    .Q(\tms1x00.O_pla_ors[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _11331_ (.CLK(clknet_leaf_76_wb_clk_i),
    .D(_01136_),
    .Q(\tms1x00.O_pla_ors[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _11332_ (.CLK(clknet_leaf_78_wb_clk_i),
    .D(_01137_),
    .Q(\tms1x00.O_pla_ors[0][19] ));
 sky130_fd_sc_hd__dfxtp_4 _11333_ (.CLK(clknet_leaf_88_wb_clk_i),
    .D(_01138_),
    .Q(\tms1x00.X[0] ));
 sky130_fd_sc_hd__dfxtp_4 _11334_ (.CLK(clknet_leaf_88_wb_clk_i),
    .D(_01139_),
    .Q(\tms1x00.X[1] ));
 sky130_fd_sc_hd__dfxtp_1 _11335_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_01140_),
    .Q(\K_override[0] ));
 sky130_fd_sc_hd__dfxtp_1 _11336_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_01141_),
    .Q(\K_override[1] ));
 sky130_fd_sc_hd__dfxtp_1 _11337_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_01142_),
    .Q(\K_override[2] ));
 sky130_fd_sc_hd__dfxtp_1 _11338_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_01143_),
    .Q(\K_override[3] ));
 sky130_fd_sc_hd__dfxtp_1 _11339_ (.CLK(clknet_leaf_73_wb_clk_i),
    .D(_01144_),
    .Q(\tms1x00.O_pla_ands[15][0] ));
 sky130_fd_sc_hd__dfxtp_2 _11340_ (.CLK(clknet_leaf_73_wb_clk_i),
    .D(_01145_),
    .Q(\tms1x00.O_pla_ands[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11341_ (.CLK(clknet_leaf_72_wb_clk_i),
    .D(_01146_),
    .Q(\tms1x00.O_pla_ands[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11342_ (.CLK(clknet_leaf_73_wb_clk_i),
    .D(_01147_),
    .Q(\tms1x00.O_pla_ands[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11343_ (.CLK(clknet_leaf_73_wb_clk_i),
    .D(_01148_),
    .Q(\tms1x00.O_pla_ands[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11344_ (.CLK(clknet_leaf_72_wb_clk_i),
    .D(_01149_),
    .Q(\tms1x00.O_pla_ands[15][5] ));
 sky130_fd_sc_hd__dfxtp_2 _11345_ (.CLK(clknet_leaf_73_wb_clk_i),
    .D(_01150_),
    .Q(\tms1x00.O_pla_ands[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11346_ (.CLK(clknet_leaf_73_wb_clk_i),
    .D(_01151_),
    .Q(\tms1x00.O_pla_ands[15][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11347_ (.CLK(clknet_leaf_72_wb_clk_i),
    .D(_01152_),
    .Q(\tms1x00.O_pla_ands[15][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11348_ (.CLK(clknet_leaf_72_wb_clk_i),
    .D(_01153_),
    .Q(\tms1x00.O_pla_ands[15][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11349_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_01154_),
    .Q(\tms1x00.O_pla_ands[17][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11350_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_01155_),
    .Q(\tms1x00.O_pla_ands[17][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11351_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(_01156_),
    .Q(\tms1x00.O_pla_ands[17][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11352_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(_01157_),
    .Q(\tms1x00.O_pla_ands[17][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11353_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(_01158_),
    .Q(\tms1x00.O_pla_ands[17][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11354_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_01159_),
    .Q(\tms1x00.O_pla_ands[17][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11355_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_01160_),
    .Q(\tms1x00.O_pla_ands[17][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11356_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(_01161_),
    .Q(\tms1x00.O_pla_ands[17][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11357_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(_01162_),
    .Q(\tms1x00.O_pla_ands[17][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11358_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_01163_),
    .Q(\tms1x00.O_pla_ands[17][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11359_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_01164_),
    .Q(\tms1x00.O_pla_ands[16][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11360_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_01165_),
    .Q(\tms1x00.O_pla_ands[16][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11361_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(_01166_),
    .Q(\tms1x00.O_pla_ands[16][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11362_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(_01167_),
    .Q(\tms1x00.O_pla_ands[16][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11363_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(_01168_),
    .Q(\tms1x00.O_pla_ands[16][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11364_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_01169_),
    .Q(\tms1x00.O_pla_ands[16][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11365_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_01170_),
    .Q(\tms1x00.O_pla_ands[16][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11366_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(_01171_),
    .Q(\tms1x00.O_pla_ands[16][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11367_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(_01172_),
    .Q(\tms1x00.O_pla_ands[16][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11368_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_01173_),
    .Q(\tms1x00.O_pla_ands[16][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11369_ (.CLK(clknet_leaf_73_wb_clk_i),
    .D(_01174_),
    .Q(\tms1x00.O_pla_ands[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11370_ (.CLK(clknet_leaf_71_wb_clk_i),
    .D(_01175_),
    .Q(\tms1x00.O_pla_ands[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11371_ (.CLK(clknet_leaf_68_wb_clk_i),
    .D(_01176_),
    .Q(\tms1x00.O_pla_ands[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11372_ (.CLK(clknet_leaf_71_wb_clk_i),
    .D(_01177_),
    .Q(\tms1x00.O_pla_ands[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11373_ (.CLK(clknet_leaf_73_wb_clk_i),
    .D(_01178_),
    .Q(\tms1x00.O_pla_ands[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11374_ (.CLK(clknet_leaf_71_wb_clk_i),
    .D(_01179_),
    .Q(\tms1x00.O_pla_ands[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11375_ (.CLK(clknet_leaf_71_wb_clk_i),
    .D(_01180_),
    .Q(\tms1x00.O_pla_ands[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11376_ (.CLK(clknet_leaf_73_wb_clk_i),
    .D(_01181_),
    .Q(\tms1x00.O_pla_ands[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11377_ (.CLK(clknet_leaf_72_wb_clk_i),
    .D(_01182_),
    .Q(\tms1x00.O_pla_ands[12][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11378_ (.CLK(clknet_leaf_68_wb_clk_i),
    .D(_01183_),
    .Q(\tms1x00.O_pla_ands[12][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11379_ (.CLK(clknet_leaf_69_wb_clk_i),
    .D(_01184_),
    .Q(\tms1x00.O_pla_ands[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11380_ (.CLK(clknet_leaf_70_wb_clk_i),
    .D(_01185_),
    .Q(\tms1x00.O_pla_ands[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11381_ (.CLK(clknet_leaf_70_wb_clk_i),
    .D(_01186_),
    .Q(\tms1x00.O_pla_ands[14][2] ));
 sky130_fd_sc_hd__dfxtp_2 _11382_ (.CLK(clknet_leaf_69_wb_clk_i),
    .D(_01187_),
    .Q(\tms1x00.O_pla_ands[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11383_ (.CLK(clknet_leaf_69_wb_clk_i),
    .D(_01188_),
    .Q(\tms1x00.O_pla_ands[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11384_ (.CLK(clknet_leaf_69_wb_clk_i),
    .D(_01189_),
    .Q(\tms1x00.O_pla_ands[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11385_ (.CLK(clknet_leaf_70_wb_clk_i),
    .D(_01190_),
    .Q(\tms1x00.O_pla_ands[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11386_ (.CLK(clknet_leaf_61_wb_clk_i),
    .D(_01191_),
    .Q(\tms1x00.O_pla_ands[14][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11387_ (.CLK(clknet_leaf_69_wb_clk_i),
    .D(_01192_),
    .Q(\tms1x00.O_pla_ands[14][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11388_ (.CLK(clknet_leaf_69_wb_clk_i),
    .D(_01193_),
    .Q(\tms1x00.O_pla_ands[14][9] ));
 sky130_fd_sc_hd__dfxtp_2 _11389_ (.CLK(clknet_leaf_76_wb_clk_i),
    .D(_01194_),
    .Q(\tms1x00.O_pla_ands[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11390_ (.CLK(clknet_leaf_76_wb_clk_i),
    .D(_01195_),
    .Q(\tms1x00.O_pla_ands[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11391_ (.CLK(clknet_leaf_71_wb_clk_i),
    .D(_01196_),
    .Q(\tms1x00.O_pla_ands[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11392_ (.CLK(clknet_leaf_74_wb_clk_i),
    .D(_01197_),
    .Q(\tms1x00.O_pla_ands[13][3] ));
 sky130_fd_sc_hd__dfxtp_2 _11393_ (.CLK(clknet_leaf_76_wb_clk_i),
    .D(_01198_),
    .Q(\tms1x00.O_pla_ands[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11394_ (.CLK(clknet_leaf_71_wb_clk_i),
    .D(_01199_),
    .Q(\tms1x00.O_pla_ands[13][5] ));
 sky130_fd_sc_hd__dfxtp_2 _11395_ (.CLK(clknet_leaf_74_wb_clk_i),
    .D(_01200_),
    .Q(\tms1x00.O_pla_ands[13][6] ));
 sky130_fd_sc_hd__dfxtp_2 _11396_ (.CLK(clknet_leaf_71_wb_clk_i),
    .D(_01201_),
    .Q(\tms1x00.O_pla_ands[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11397_ (.CLK(clknet_leaf_71_wb_clk_i),
    .D(_01202_),
    .Q(\tms1x00.O_pla_ands[13][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11398_ (.CLK(clknet_leaf_71_wb_clk_i),
    .D(_01203_),
    .Q(\tms1x00.O_pla_ands[13][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11399_ (.CLK(clknet_leaf_112_wb_clk_i),
    .D(_01204_),
    .Q(\tms1x00.ins_pla_ors[7][27] ));
 sky130_fd_sc_hd__dfxtp_1 _11400_ (.CLK(clknet_leaf_112_wb_clk_i),
    .D(_01205_),
    .Q(\tms1x00.ins_pla_ors[7][28] ));
 sky130_fd_sc_hd__dfxtp_1 _11401_ (.CLK(clknet_leaf_120_wb_clk_i),
    .D(_01206_),
    .Q(\tms1x00.ins_pla_ors[7][29] ));
 sky130_fd_sc_hd__dfxtp_2 _11402_ (.CLK(clknet_leaf_74_wb_clk_i),
    .D(_01207_),
    .Q(\tms1x00.O_pla_ands[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11403_ (.CLK(clknet_leaf_74_wb_clk_i),
    .D(_01208_),
    .Q(\tms1x00.O_pla_ands[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11404_ (.CLK(clknet_leaf_73_wb_clk_i),
    .D(_01209_),
    .Q(\tms1x00.O_pla_ands[10][2] ));
 sky130_fd_sc_hd__dfxtp_2 _11405_ (.CLK(clknet_leaf_74_wb_clk_i),
    .D(_01210_),
    .Q(\tms1x00.O_pla_ands[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11406_ (.CLK(clknet_leaf_73_wb_clk_i),
    .D(_01211_),
    .Q(\tms1x00.O_pla_ands[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11407_ (.CLK(clknet_leaf_71_wb_clk_i),
    .D(_01212_),
    .Q(\tms1x00.O_pla_ands[10][5] ));
 sky130_fd_sc_hd__dfxtp_2 _11408_ (.CLK(clknet_leaf_74_wb_clk_i),
    .D(_01213_),
    .Q(\tms1x00.O_pla_ands[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11409_ (.CLK(clknet_leaf_74_wb_clk_i),
    .D(_01214_),
    .Q(\tms1x00.O_pla_ands[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11410_ (.CLK(clknet_leaf_71_wb_clk_i),
    .D(_01215_),
    .Q(\tms1x00.O_pla_ands[10][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11411_ (.CLK(clknet_leaf_74_wb_clk_i),
    .D(_01216_),
    .Q(\tms1x00.O_pla_ands[10][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11412_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_01217_),
    .Q(\tms1x00.O_pla_ands[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11413_ (.CLK(clknet_leaf_67_wb_clk_i),
    .D(_01218_),
    .Q(\tms1x00.O_pla_ands[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11414_ (.CLK(clknet_leaf_67_wb_clk_i),
    .D(_01219_),
    .Q(\tms1x00.O_pla_ands[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11415_ (.CLK(clknet_leaf_67_wb_clk_i),
    .D(_01220_),
    .Q(\tms1x00.O_pla_ands[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11416_ (.CLK(clknet_leaf_67_wb_clk_i),
    .D(_01221_),
    .Q(\tms1x00.O_pla_ands[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11417_ (.CLK(clknet_leaf_67_wb_clk_i),
    .D(_01222_),
    .Q(\tms1x00.O_pla_ands[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11418_ (.CLK(clknet_leaf_67_wb_clk_i),
    .D(_01223_),
    .Q(\tms1x00.O_pla_ands[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11419_ (.CLK(clknet_leaf_67_wb_clk_i),
    .D(_01224_),
    .Q(\tms1x00.O_pla_ands[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11420_ (.CLK(clknet_leaf_67_wb_clk_i),
    .D(_01225_),
    .Q(\tms1x00.O_pla_ands[9][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11421_ (.CLK(clknet_leaf_67_wb_clk_i),
    .D(_01226_),
    .Q(\tms1x00.O_pla_ands[9][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11422_ (.CLK(clknet_leaf_69_wb_clk_i),
    .D(_01227_),
    .Q(\tms1x00.O_pla_ands[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11423_ (.CLK(clknet_leaf_68_wb_clk_i),
    .D(_01228_),
    .Q(\tms1x00.O_pla_ands[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11424_ (.CLK(clknet_leaf_68_wb_clk_i),
    .D(_01229_),
    .Q(\tms1x00.O_pla_ands[11][2] ));
 sky130_fd_sc_hd__dfxtp_2 _11425_ (.CLK(clknet_leaf_69_wb_clk_i),
    .D(_01230_),
    .Q(\tms1x00.O_pla_ands[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11426_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_01231_),
    .Q(\tms1x00.O_pla_ands[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11427_ (.CLK(clknet_leaf_68_wb_clk_i),
    .D(_01232_),
    .Q(\tms1x00.O_pla_ands[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11428_ (.CLK(clknet_leaf_69_wb_clk_i),
    .D(_01233_),
    .Q(\tms1x00.O_pla_ands[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11429_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_01234_),
    .Q(\tms1x00.O_pla_ands[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11430_ (.CLK(clknet_leaf_68_wb_clk_i),
    .D(_01235_),
    .Q(\tms1x00.O_pla_ands[11][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11431_ (.CLK(clknet_leaf_68_wb_clk_i),
    .D(_01236_),
    .Q(\tms1x00.O_pla_ands[11][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11432_ (.CLK(clknet_leaf_94_wb_clk_i),
    .D(_01237_),
    .Q(\tms1x00.ins_pla_ors[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11433_ (.CLK(clknet_leaf_94_wb_clk_i),
    .D(_01238_),
    .Q(\tms1x00.ins_pla_ors[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11434_ (.CLK(clknet_leaf_96_wb_clk_i),
    .D(_01239_),
    .Q(\tms1x00.ins_pla_ors[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11435_ (.CLK(clknet_leaf_94_wb_clk_i),
    .D(_01240_),
    .Q(\tms1x00.ins_pla_ors[3][12] ));
 sky130_fd_sc_hd__dfxtp_2 _11436_ (.CLK(clknet_leaf_106_wb_clk_i),
    .D(_01241_),
    .Q(\tms1x00.ins_pla_ors[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _11437_ (.CLK(clknet_leaf_108_wb_clk_i),
    .D(_01242_),
    .Q(\tms1x00.ins_pla_ors[3][21] ));
 sky130_fd_sc_hd__dfxtp_1 _11438_ (.CLK(clknet_leaf_94_wb_clk_i),
    .D(_01243_),
    .Q(\tms1x00.ins_pla_ors[3][24] ));
 sky130_fd_sc_hd__dfxtp_1 _11439_ (.CLK(clknet_leaf_111_wb_clk_i),
    .D(_01244_),
    .Q(\tms1x00.ins_pla_ors[3][25] ));
 sky130_fd_sc_hd__dfxtp_1 _11440_ (.CLK(clknet_leaf_94_wb_clk_i),
    .D(_01245_),
    .Q(\tms1x00.ins_pla_ors[3][29] ));
 sky130_fd_sc_hd__dfxtp_1 _11441_ (.CLK(clknet_leaf_96_wb_clk_i),
    .D(_01246_),
    .Q(\tms1x00.ins_pla_ors[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11442_ (.CLK(clknet_leaf_96_wb_clk_i),
    .D(_01247_),
    .Q(\tms1x00.ins_pla_ors[6][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11443_ (.CLK(clknet_leaf_105_wb_clk_i),
    .D(_01248_),
    .Q(\tms1x00.ins_pla_ors[6][12] ));
 sky130_fd_sc_hd__dfxtp_2 _11444_ (.CLK(clknet_leaf_94_wb_clk_i),
    .D(_01249_),
    .Q(\tms1x00.ins_pla_ors[6][16] ));
 sky130_fd_sc_hd__dfxtp_1 _11445_ (.CLK(clknet_leaf_94_wb_clk_i),
    .D(_01250_),
    .Q(\tms1x00.ins_pla_ors[6][18] ));
 sky130_fd_sc_hd__dfxtp_1 _11446_ (.CLK(clknet_leaf_105_wb_clk_i),
    .D(_01251_),
    .Q(\tms1x00.ins_pla_ors[6][25] ));
 sky130_fd_sc_hd__dfxtp_1 _11447_ (.CLK(clknet_leaf_108_wb_clk_i),
    .D(_01252_),
    .Q(\tms1x00.ins_pla_ors[6][26] ));
 sky130_fd_sc_hd__dfxtp_1 _11448_ (.CLK(clknet_leaf_105_wb_clk_i),
    .D(_01253_),
    .Q(\tms1x00.ins_pla_ors[6][27] ));
 sky130_fd_sc_hd__dfxtp_1 _11449_ (.CLK(clknet_leaf_112_wb_clk_i),
    .D(_01254_),
    .Q(\tms1x00.ins_pla_ors[6][28] ));
 sky130_fd_sc_hd__dfxtp_1 _11450_ (.CLK(clknet_leaf_105_wb_clk_i),
    .D(_01255_),
    .Q(\tms1x00.ins_pla_ors[6][29] ));
 sky130_fd_sc_hd__dfxtp_2 _11451_ (.CLK(clknet_leaf_91_wb_clk_i),
    .D(_01256_),
    .Q(\tms1x00.ins_pla_ors[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11452_ (.CLK(clknet_leaf_93_wb_clk_i),
    .D(_01257_),
    .Q(\tms1x00.ins_pla_ors[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11453_ (.CLK(clknet_leaf_92_wb_clk_i),
    .D(_01258_),
    .Q(\tms1x00.ins_pla_ors[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11454_ (.CLK(clknet_leaf_90_wb_clk_i),
    .D(_01259_),
    .Q(\tms1x00.ins_pla_ors[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11455_ (.CLK(clknet_leaf_91_wb_clk_i),
    .D(_01260_),
    .Q(\tms1x00.ins_pla_ors[5][7] ));
 sky130_fd_sc_hd__dfxtp_2 _11456_ (.CLK(clknet_leaf_93_wb_clk_i),
    .D(_01261_),
    .Q(\tms1x00.ins_pla_ors[5][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11457_ (.CLK(clknet_leaf_106_wb_clk_i),
    .D(_01262_),
    .Q(\tms1x00.ins_pla_ors[5][16] ));
 sky130_fd_sc_hd__dfxtp_1 _11458_ (.CLK(clknet_leaf_108_wb_clk_i),
    .D(_01263_),
    .Q(\tms1x00.ins_pla_ors[5][21] ));
 sky130_fd_sc_hd__dfxtp_1 _11459_ (.CLK(clknet_leaf_94_wb_clk_i),
    .D(_01264_),
    .Q(\tms1x00.ins_pla_ors[5][24] ));
 sky130_fd_sc_hd__dfxtp_2 _11460_ (.CLK(clknet_leaf_113_wb_clk_i),
    .D(_01265_),
    .Q(\tms1x00.ins_pla_ors[5][26] ));
 sky130_fd_sc_hd__dfxtp_1 _11461_ (.CLK(clknet_leaf_112_wb_clk_i),
    .D(_01266_),
    .Q(\tms1x00.ins_pla_ors[5][27] ));
 sky130_fd_sc_hd__dfxtp_1 _11462_ (.CLK(clknet_leaf_112_wb_clk_i),
    .D(_01267_),
    .Q(\tms1x00.ins_pla_ors[5][28] ));
 sky130_fd_sc_hd__dfxtp_1 _11463_ (.CLK(clknet_leaf_94_wb_clk_i),
    .D(_01268_),
    .Q(\tms1x00.ins_pla_ors[5][29] ));
 sky130_fd_sc_hd__dfxtp_1 _11464_ (.CLK(clknet_leaf_92_wb_clk_i),
    .D(_01269_),
    .Q(\tms1x00.ins_pla_ors[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11465_ (.CLK(clknet_leaf_92_wb_clk_i),
    .D(_01270_),
    .Q(\tms1x00.ins_pla_ors[4][6] ));
 sky130_fd_sc_hd__dfxtp_2 _11466_ (.CLK(clknet_leaf_93_wb_clk_i),
    .D(_01271_),
    .Q(\tms1x00.ins_pla_ors[4][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11467_ (.CLK(clknet_leaf_93_wb_clk_i),
    .D(_01272_),
    .Q(\tms1x00.ins_pla_ors[4][11] ));
 sky130_fd_sc_hd__dfxtp_1 _11468_ (.CLK(clknet_leaf_113_wb_clk_i),
    .D(_01273_),
    .Q(\tms1x00.ins_pla_ors[4][14] ));
 sky130_fd_sc_hd__dfxtp_2 _11469_ (.CLK(clknet_leaf_93_wb_clk_i),
    .D(_01274_),
    .Q(\tms1x00.ins_pla_ors[4][16] ));
 sky130_fd_sc_hd__dfxtp_2 _11470_ (.CLK(clknet_leaf_103_wb_clk_i),
    .D(_01275_),
    .Q(\tms1x00.ins_pla_ors[4][17] ));
 sky130_fd_sc_hd__dfxtp_1 _11471_ (.CLK(clknet_leaf_93_wb_clk_i),
    .D(_01276_),
    .Q(\tms1x00.ins_pla_ors[4][18] ));
 sky130_fd_sc_hd__dfxtp_2 _11472_ (.CLK(clknet_leaf_104_wb_clk_i),
    .D(_01277_),
    .Q(\tms1x00.ins_pla_ors[4][24] ));
 sky130_fd_sc_hd__dfxtp_1 _11473_ (.CLK(clknet_leaf_94_wb_clk_i),
    .D(_01278_),
    .Q(\tms1x00.ins_pla_ors[4][25] ));
 sky130_fd_sc_hd__dfxtp_1 _11474_ (.CLK(clknet_leaf_113_wb_clk_i),
    .D(_01279_),
    .Q(\tms1x00.ins_pla_ors[4][26] ));
 sky130_fd_sc_hd__dfxtp_1 _11475_ (.CLK(clknet_leaf_120_wb_clk_i),
    .D(_01280_),
    .Q(\tms1x00.ins_pla_ors[4][27] ));
 sky130_fd_sc_hd__dfxtp_1 _11476_ (.CLK(clknet_leaf_121_wb_clk_i),
    .D(_01281_),
    .Q(\tms1x00.ins_pla_ors[4][28] ));
 sky130_fd_sc_hd__dfxtp_1 _11477_ (.CLK(clknet_leaf_121_wb_clk_i),
    .D(_01282_),
    .Q(\tms1x00.ins_pla_ors[4][29] ));
 sky130_fd_sc_hd__dfxtp_2 _11478_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_01283_),
    .Q(\tms1x00.O_pla_ands[7][0] ));
 sky130_fd_sc_hd__dfxtp_2 _11479_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_01284_),
    .Q(\tms1x00.O_pla_ands[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11480_ (.CLK(clknet_leaf_63_wb_clk_i),
    .D(_01285_),
    .Q(\tms1x00.O_pla_ands[7][2] ));
 sky130_fd_sc_hd__dfxtp_2 _11481_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_01286_),
    .Q(\tms1x00.O_pla_ands[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11482_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_01287_),
    .Q(\tms1x00.O_pla_ands[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11483_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_01288_),
    .Q(\tms1x00.O_pla_ands[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11484_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_01289_),
    .Q(\tms1x00.O_pla_ands[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11485_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_01290_),
    .Q(\tms1x00.O_pla_ands[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11486_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_01291_),
    .Q(\tms1x00.O_pla_ands[7][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11487_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_01292_),
    .Q(\tms1x00.O_pla_ands[7][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11488_ (.CLK(clknet_leaf_72_wb_clk_i),
    .D(_01293_),
    .Q(\tms1x00.O_pla_ands[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11489_ (.CLK(clknet_leaf_72_wb_clk_i),
    .D(_01294_),
    .Q(\tms1x00.O_pla_ands[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11490_ (.CLK(clknet_leaf_72_wb_clk_i),
    .D(_01295_),
    .Q(\tms1x00.O_pla_ands[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11491_ (.CLK(clknet_leaf_73_wb_clk_i),
    .D(_01296_),
    .Q(\tms1x00.O_pla_ands[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11492_ (.CLK(clknet_leaf_72_wb_clk_i),
    .D(_01297_),
    .Q(\tms1x00.O_pla_ands[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11493_ (.CLK(clknet_leaf_72_wb_clk_i),
    .D(_01298_),
    .Q(\tms1x00.O_pla_ands[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11494_ (.CLK(clknet_leaf_72_wb_clk_i),
    .D(_01299_),
    .Q(\tms1x00.O_pla_ands[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11495_ (.CLK(clknet_leaf_73_wb_clk_i),
    .D(_01300_),
    .Q(\tms1x00.O_pla_ands[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11496_ (.CLK(clknet_leaf_72_wb_clk_i),
    .D(_01301_),
    .Q(\tms1x00.O_pla_ands[8][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11497_ (.CLK(clknet_leaf_72_wb_clk_i),
    .D(_01302_),
    .Q(\tms1x00.O_pla_ands[8][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11498_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_01303_),
    .Q(\tms1x00.O_pla_ands[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11499_ (.CLK(clknet_leaf_64_wb_clk_i),
    .D(_01304_),
    .Q(\tms1x00.O_pla_ands[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11500_ (.CLK(clknet_leaf_65_wb_clk_i),
    .D(_01305_),
    .Q(\tms1x00.O_pla_ands[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11501_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_01306_),
    .Q(\tms1x00.O_pla_ands[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11502_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_01307_),
    .Q(\tms1x00.O_pla_ands[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11503_ (.CLK(clknet_leaf_65_wb_clk_i),
    .D(_01308_),
    .Q(\tms1x00.O_pla_ands[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11504_ (.CLK(clknet_leaf_65_wb_clk_i),
    .D(_01309_),
    .Q(\tms1x00.O_pla_ands[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11505_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_01310_),
    .Q(\tms1x00.O_pla_ands[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11506_ (.CLK(clknet_leaf_65_wb_clk_i),
    .D(_01311_),
    .Q(\tms1x00.O_pla_ands[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11507_ (.CLK(clknet_leaf_65_wb_clk_i),
    .D(_01312_),
    .Q(\tms1x00.O_pla_ands[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11508_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_01313_),
    .Q(\tms1x00.O_pla_ands[25][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11509_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_01314_),
    .Q(\tms1x00.O_pla_ands[25][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11510_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_01315_),
    .Q(\tms1x00.O_pla_ands[25][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11511_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_01316_),
    .Q(\tms1x00.O_pla_ands[25][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11512_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_01317_),
    .Q(\tms1x00.O_pla_ands[25][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11513_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_01318_),
    .Q(\tms1x00.O_pla_ands[25][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11514_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_01319_),
    .Q(\tms1x00.O_pla_ands[25][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11515_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_01320_),
    .Q(\tms1x00.O_pla_ands[25][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11516_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_01321_),
    .Q(\tms1x00.O_pla_ands[25][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11517_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_01322_),
    .Q(\tms1x00.O_pla_ands[25][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11518_ (.CLK(clknet_leaf_61_wb_clk_i),
    .D(_01323_),
    .Q(\tms1x00.O_pla_ands[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11519_ (.CLK(clknet_leaf_63_wb_clk_i),
    .D(_01324_),
    .Q(\tms1x00.O_pla_ands[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11520_ (.CLK(clknet_leaf_62_wb_clk_i),
    .D(_01325_),
    .Q(\tms1x00.O_pla_ands[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11521_ (.CLK(clknet_leaf_61_wb_clk_i),
    .D(_01326_),
    .Q(\tms1x00.O_pla_ands[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11522_ (.CLK(clknet_leaf_61_wb_clk_i),
    .D(_01327_),
    .Q(\tms1x00.O_pla_ands[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11523_ (.CLK(clknet_leaf_63_wb_clk_i),
    .D(_01328_),
    .Q(\tms1x00.O_pla_ands[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11524_ (.CLK(clknet_leaf_62_wb_clk_i),
    .D(_01329_),
    .Q(\tms1x00.O_pla_ands[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11525_ (.CLK(clknet_leaf_61_wb_clk_i),
    .D(_01330_),
    .Q(\tms1x00.O_pla_ands[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11526_ (.CLK(clknet_leaf_63_wb_clk_i),
    .D(_01331_),
    .Q(\tms1x00.O_pla_ands[6][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11527_ (.CLK(clknet_leaf_62_wb_clk_i),
    .D(_01332_),
    .Q(\tms1x00.O_pla_ands[6][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11528_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_01333_),
    .Q(\tms1x00.O_pla_ands[26][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11529_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_01334_),
    .Q(\tms1x00.O_pla_ands[26][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11530_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_01335_),
    .Q(\tms1x00.O_pla_ands[26][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11531_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_01336_),
    .Q(\tms1x00.O_pla_ands[26][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11532_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_01337_),
    .Q(\tms1x00.O_pla_ands[26][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11533_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_01338_),
    .Q(\tms1x00.O_pla_ands[26][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11534_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_01339_),
    .Q(\tms1x00.O_pla_ands[26][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11535_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_01340_),
    .Q(\tms1x00.O_pla_ands[26][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11536_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_01341_),
    .Q(\tms1x00.O_pla_ands[26][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11537_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_01342_),
    .Q(\tms1x00.O_pla_ands[26][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11538_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_01343_),
    .Q(\tms1x00.O_pla_ands[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11539_ (.CLK(clknet_leaf_65_wb_clk_i),
    .D(_01344_),
    .Q(\tms1x00.O_pla_ands[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11540_ (.CLK(clknet_leaf_65_wb_clk_i),
    .D(_01345_),
    .Q(\tms1x00.O_pla_ands[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11541_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_01346_),
    .Q(\tms1x00.O_pla_ands[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11542_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_01347_),
    .Q(\tms1x00.O_pla_ands[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11543_ (.CLK(clknet_leaf_65_wb_clk_i),
    .D(_01348_),
    .Q(\tms1x00.O_pla_ands[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11544_ (.CLK(clknet_leaf_64_wb_clk_i),
    .D(_01349_),
    .Q(\tms1x00.O_pla_ands[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11545_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_01350_),
    .Q(\tms1x00.O_pla_ands[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11546_ (.CLK(clknet_leaf_65_wb_clk_i),
    .D(_01351_),
    .Q(\tms1x00.O_pla_ands[5][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11547_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_01352_),
    .Q(\tms1x00.O_pla_ands[5][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11548_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_01353_),
    .Q(\tms1x00.O_pla_ands[23][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11549_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_01354_),
    .Q(\tms1x00.O_pla_ands[23][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11550_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_01355_),
    .Q(\tms1x00.O_pla_ands[23][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11551_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_01356_),
    .Q(\tms1x00.O_pla_ands[23][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11552_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_01357_),
    .Q(\tms1x00.O_pla_ands[23][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11553_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_01358_),
    .Q(\tms1x00.O_pla_ands[23][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11554_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_01359_),
    .Q(\tms1x00.O_pla_ands[23][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11555_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_01360_),
    .Q(\tms1x00.O_pla_ands[23][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11556_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_01361_),
    .Q(\tms1x00.O_pla_ands[23][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11557_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_01362_),
    .Q(\tms1x00.O_pla_ands[23][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11558_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_01363_),
    .Q(\tms1x00.O_pla_ands[22][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11559_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_01364_),
    .Q(\tms1x00.O_pla_ands[22][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11560_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(_01365_),
    .Q(\tms1x00.O_pla_ands[22][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11561_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_01366_),
    .Q(\tms1x00.O_pla_ands[22][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11562_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_01367_),
    .Q(\tms1x00.O_pla_ands[22][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11563_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(_01368_),
    .Q(\tms1x00.O_pla_ands[22][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11564_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_01369_),
    .Q(\tms1x00.O_pla_ands[22][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11565_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_01370_),
    .Q(\tms1x00.O_pla_ands[22][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11566_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_01371_),
    .Q(\tms1x00.O_pla_ands[22][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11567_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_01372_),
    .Q(\tms1x00.O_pla_ands[22][9] ));
 sky130_fd_sc_hd__dfxtp_2 _11568_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_01373_),
    .Q(\tms1x00.wb_step_state ));
 sky130_fd_sc_hd__dfxtp_2 _11569_ (.CLK(clknet_leaf_81_wb_clk_i),
    .D(_01374_),
    .Q(net146));
 sky130_fd_sc_hd__dfxtp_1 _11570_ (.CLK(clknet_leaf_81_wb_clk_i),
    .D(_01375_),
    .Q(net147));
 sky130_fd_sc_hd__dfxtp_1 _11571_ (.CLK(clknet_leaf_81_wb_clk_i),
    .D(_01376_),
    .Q(net148));
 sky130_fd_sc_hd__dfxtp_1 _11572_ (.CLK(clknet_leaf_80_wb_clk_i),
    .D(_01377_),
    .Q(net149));
 sky130_fd_sc_hd__dfxtp_2 _11573_ (.CLK(clknet_leaf_81_wb_clk_i),
    .D(_01378_),
    .Q(net150));
 sky130_fd_sc_hd__dfxtp_4 _11574_ (.CLK(clknet_leaf_82_wb_clk_i),
    .D(_01379_),
    .Q(net151));
 sky130_fd_sc_hd__dfxtp_4 _11575_ (.CLK(clknet_leaf_82_wb_clk_i),
    .D(_01380_),
    .Q(net152));
 sky130_fd_sc_hd__dfxtp_4 _11576_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_01381_),
    .Q(\tms1x00.rom_addr[0] ));
 sky130_fd_sc_hd__dfxtp_2 _11577_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_01382_),
    .Q(\tms1x00.rom_addr[1] ));
 sky130_fd_sc_hd__dfxtp_2 _11578_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_01383_),
    .Q(net158));
 sky130_fd_sc_hd__dfxtp_2 _11579_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_01384_),
    .Q(net159));
 sky130_fd_sc_hd__dfxtp_1 _11580_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_01385_),
    .Q(net160));
 sky130_fd_sc_hd__dfxtp_1 _11581_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_01386_),
    .Q(net161));
 sky130_fd_sc_hd__dfxtp_1 _11582_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_01387_),
    .Q(net162));
 sky130_fd_sc_hd__dfxtp_1 _11583_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_01388_),
    .Q(net163));
 sky130_fd_sc_hd__dfxtp_1 _11584_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_01389_),
    .Q(net164));
 sky130_fd_sc_hd__dfxtp_1 _11585_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_01390_),
    .Q(net165));
 sky130_fd_sc_hd__dfxtp_1 _11586_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_01391_),
    .Q(net166));
 sky130_fd_sc_hd__dfxtp_4 _11587_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_01392_),
    .Q(net144));
 sky130_fd_sc_hd__dfxtp_1 _11588_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_01393_),
    .Q(\tms1x00.SR[0] ));
 sky130_fd_sc_hd__dfxtp_1 _11589_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_01394_),
    .Q(\tms1x00.SR[1] ));
 sky130_fd_sc_hd__dfxtp_1 _11590_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_01395_),
    .Q(\tms1x00.SR[2] ));
 sky130_fd_sc_hd__dfxtp_1 _11591_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_01396_),
    .Q(\tms1x00.SR[3] ));
 sky130_fd_sc_hd__dfxtp_1 _11592_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_01397_),
    .Q(\tms1x00.SR[4] ));
 sky130_fd_sc_hd__dfxtp_1 _11593_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_01398_),
    .Q(\tms1x00.SR[5] ));
 sky130_fd_sc_hd__dfxtp_4 _11594_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_01399_),
    .Q(\tms1x00.B[1] ));
 sky130_fd_sc_hd__dfxtp_4 _11595_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_01400_),
    .Q(\tms1x00.B[0] ));
 sky130_fd_sc_hd__dfxtp_4 _11596_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_01401_),
    .Q(\tms1x00.ins_arg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _11597_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_01402_),
    .Q(\tms1x00.ins_arg[4] ));
 sky130_fd_sc_hd__dfxtp_4 _11598_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_01403_),
    .Q(\tms1x00.ins_arg[3] ));
 sky130_fd_sc_hd__dfxtp_4 _11599_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_01404_),
    .Q(\tms1x00.ins_arg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _11600_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_01405_),
    .Q(\tms1x00.ins_arg[1] ));
 sky130_fd_sc_hd__dfxtp_4 _11601_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_01406_),
    .Q(\tms1x00.ins_arg[0] ));
 sky130_fd_sc_hd__dfxtp_4 _11602_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_01407_),
    .Q(\tms1x00.cycle[0] ));
 sky130_fd_sc_hd__dfxtp_2 _11603_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_01408_),
    .Q(\tms1x00.cycle[1] ));
 sky130_fd_sc_hd__dfxtp_2 _11604_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_01409_),
    .Q(\tms1x00.cycle[2] ));
 sky130_fd_sc_hd__dfxtp_4 _11605_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(\tms1x00.K_in[0] ),
    .Q(\tms1x00.K_latch[0] ));
 sky130_fd_sc_hd__dfxtp_4 _11606_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(\tms1x00.K_in[1] ),
    .Q(\tms1x00.K_latch[1] ));
 sky130_fd_sc_hd__dfxtp_2 _11607_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(\tms1x00.K_in[2] ),
    .Q(\tms1x00.K_latch[2] ));
 sky130_fd_sc_hd__dfxtp_4 _11608_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(\tms1x00.K_in[3] ),
    .Q(\tms1x00.K_latch[3] ));
 sky130_fd_sc_hd__dfxtp_4 _11609_ (.CLK(clknet_leaf_87_wb_clk_i),
    .D(_01410_),
    .Q(net129));
 sky130_fd_sc_hd__dfxtp_4 _11610_ (.CLK(clknet_leaf_87_wb_clk_i),
    .D(_01411_),
    .Q(net130));
 sky130_fd_sc_hd__dfxtp_4 _11611_ (.CLK(clknet_leaf_83_wb_clk_i),
    .D(_01412_),
    .Q(net131));
 sky130_fd_sc_hd__dfxtp_4 _11612_ (.CLK(clknet_leaf_86_wb_clk_i),
    .D(_01413_),
    .Q(net132));
 sky130_fd_sc_hd__dfxtp_4 _11613_ (.CLK(clknet_leaf_86_wb_clk_i),
    .D(_01414_),
    .Q(net133));
 sky130_fd_sc_hd__dfxtp_4 _11614_ (.CLK(clknet_leaf_87_wb_clk_i),
    .D(_01415_),
    .Q(net134));
 sky130_fd_sc_hd__dfxtp_4 _11615_ (.CLK(clknet_leaf_87_wb_clk_i),
    .D(_01416_),
    .Q(net135));
 sky130_fd_sc_hd__dfxtp_4 _11616_ (.CLK(clknet_leaf_86_wb_clk_i),
    .D(_01417_),
    .Q(net136));
 sky130_fd_sc_hd__dfxtp_4 _11617_ (.CLK(clknet_leaf_87_wb_clk_i),
    .D(_01418_),
    .Q(net137));
 sky130_fd_sc_hd__dfxtp_4 _11618_ (.CLK(clknet_leaf_83_wb_clk_i),
    .D(_01419_),
    .Q(net138));
 sky130_fd_sc_hd__dfxtp_4 _11619_ (.CLK(clknet_leaf_83_wb_clk_i),
    .D(_01420_),
    .Q(net139));
 sky130_fd_sc_hd__dfxtp_4 _11620_ (.CLK(clknet_leaf_86_wb_clk_i),
    .D(_01421_),
    .Q(net140));
 sky130_fd_sc_hd__dfxtp_4 _11621_ (.CLK(clknet_leaf_86_wb_clk_i),
    .D(_01422_),
    .Q(net141));
 sky130_fd_sc_hd__dfxtp_4 _11622_ (.CLK(clknet_leaf_83_wb_clk_i),
    .D(_01423_),
    .Q(net142));
 sky130_fd_sc_hd__dfxtp_4 _11623_ (.CLK(clknet_leaf_87_wb_clk_i),
    .D(_01424_),
    .Q(net143));
 sky130_fd_sc_hd__dfxtp_4 _11624_ (.CLK(clknet_leaf_86_wb_clk_i),
    .D(_01425_),
    .Q(\tms1x00.O_latch[0] ));
 sky130_fd_sc_hd__dfxtp_4 _11625_ (.CLK(clknet_leaf_88_wb_clk_i),
    .D(_01426_),
    .Q(\tms1x00.O_latch[1] ));
 sky130_fd_sc_hd__dfxtp_4 _11626_ (.CLK(clknet_leaf_88_wb_clk_i),
    .D(_01427_),
    .Q(\tms1x00.O_latch[2] ));
 sky130_fd_sc_hd__dfxtp_4 _11627_ (.CLK(clknet_leaf_88_wb_clk_i),
    .D(_01428_),
    .Q(\tms1x00.O_latch[3] ));
 sky130_fd_sc_hd__dfxtp_4 _11628_ (.CLK(clknet_leaf_56_wb_clk_i),
    .D(_01429_),
    .Q(\tms1x00.O_latch[4] ));
 sky130_fd_sc_hd__dfxtp_4 _11629_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_01430_),
    .Q(\tms1x00.CL ));
 sky130_fd_sc_hd__dfxtp_1 _11630_ (.CLK(clknet_leaf_126_wb_clk_i),
    .D(_01431_),
    .Q(\tms1x00.SL ));
 sky130_fd_sc_hd__dfxtp_4 _11631_ (.CLK(clknet_leaf_126_wb_clk_i),
    .D(_01432_),
    .Q(\tms1x00.status ));
 sky130_fd_sc_hd__dfxtp_1 _11632_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_01433_),
    .Q(\tms1x00.CS ));
 sky130_fd_sc_hd__dfxtp_1 _11633_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_01434_),
    .Q(\tms1x00.CB ));
 sky130_fd_sc_hd__dfxtp_2 _11634_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_01435_),
    .Q(\tms1x00.CA ));
 sky130_fd_sc_hd__dfxtp_1 _11635_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_01436_),
    .Q(\tms1x00.PB[0] ));
 sky130_fd_sc_hd__dfxtp_1 _11636_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_01437_),
    .Q(\tms1x00.PB[1] ));
 sky130_fd_sc_hd__dfxtp_1 _11637_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_01438_),
    .Q(\tms1x00.PB[2] ));
 sky130_fd_sc_hd__dfxtp_1 _11638_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_01439_),
    .Q(\tms1x00.PB[3] ));
 sky130_fd_sc_hd__dfxtp_1 _11639_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_01440_),
    .Q(\tms1x00.PA[0] ));
 sky130_fd_sc_hd__dfxtp_1 _11640_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_01441_),
    .Q(\tms1x00.PA[1] ));
 sky130_fd_sc_hd__dfxtp_1 _11641_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_01442_),
    .Q(\tms1x00.PA[2] ));
 sky130_fd_sc_hd__dfxtp_1 _11642_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_01443_),
    .Q(\tms1x00.PA[3] ));
 sky130_fd_sc_hd__dfxtp_2 _11643_ (.CLK(clknet_leaf_90_wb_clk_i),
    .D(_01444_),
    .Q(\tms1x00.P[0] ));
 sky130_fd_sc_hd__dfxtp_1 _11644_ (.CLK(clknet_leaf_91_wb_clk_i),
    .D(_01445_),
    .Q(\tms1x00.P[1] ));
 sky130_fd_sc_hd__dfxtp_1 _11645_ (.CLK(clknet_leaf_89_wb_clk_i),
    .D(_01446_),
    .Q(\tms1x00.P[2] ));
 sky130_fd_sc_hd__dfxtp_1 _11646_ (.CLK(clknet_leaf_89_wb_clk_i),
    .D(_01447_),
    .Q(\tms1x00.P[3] ));
 sky130_fd_sc_hd__dfxtp_2 _11647_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_01448_),
    .Q(\tms1x00.PC[0] ));
 sky130_fd_sc_hd__dfxtp_2 _11648_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_01449_),
    .Q(\tms1x00.PC[1] ));
 sky130_fd_sc_hd__dfxtp_2 _11649_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_01450_),
    .Q(\tms1x00.PC[2] ));
 sky130_fd_sc_hd__dfxtp_2 _11650_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_01451_),
    .Q(\tms1x00.PC[3] ));
 sky130_fd_sc_hd__dfxtp_4 _11651_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_01452_),
    .Q(\tms1x00.PC[4] ));
 sky130_fd_sc_hd__dfxtp_2 _11652_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_01453_),
    .Q(\tms1x00.PC[5] ));
 sky130_fd_sc_hd__dfxtp_2 _11653_ (.CLK(clknet_leaf_87_wb_clk_i),
    .D(_01454_),
    .Q(\tms1x00.Y[0] ));
 sky130_fd_sc_hd__dfxtp_2 _11654_ (.CLK(clknet_leaf_87_wb_clk_i),
    .D(_01455_),
    .Q(\tms1x00.Y[1] ));
 sky130_fd_sc_hd__dfxtp_1 _11655_ (.CLK(clknet_leaf_87_wb_clk_i),
    .D(_01456_),
    .Q(\tms1x00.Y[2] ));
 sky130_fd_sc_hd__dfxtp_1 _11656_ (.CLK(clknet_leaf_87_wb_clk_i),
    .D(_01457_),
    .Q(\tms1x00.Y[3] ));
 sky130_fd_sc_hd__dfxtp_4 _11657_ (.CLK(clknet_leaf_88_wb_clk_i),
    .D(_01458_),
    .Q(\tms1x00.X[2] ));
 sky130_fd_sc_hd__dfxtp_1 _11658_ (.CLK(clknet_leaf_90_wb_clk_i),
    .D(_01459_),
    .Q(\tms1x00.N[0] ));
 sky130_fd_sc_hd__dfxtp_1 _11659_ (.CLK(clknet_leaf_90_wb_clk_i),
    .D(_01460_),
    .Q(\tms1x00.N[1] ));
 sky130_fd_sc_hd__dfxtp_1 _11660_ (.CLK(clknet_leaf_89_wb_clk_i),
    .D(_01461_),
    .Q(\tms1x00.N[2] ));
 sky130_fd_sc_hd__dfxtp_1 _11661_ (.CLK(clknet_leaf_90_wb_clk_i),
    .D(_01462_),
    .Q(\tms1x00.N[3] ));
 sky130_fd_sc_hd__dfxtp_2 _11662_ (.CLK(clknet_leaf_87_wb_clk_i),
    .D(_01463_),
    .Q(\tms1x00.A[0] ));
 sky130_fd_sc_hd__dfxtp_2 _11663_ (.CLK(clknet_leaf_87_wb_clk_i),
    .D(_01464_),
    .Q(\tms1x00.A[1] ));
 sky130_fd_sc_hd__dfxtp_2 _11664_ (.CLK(clknet_leaf_89_wb_clk_i),
    .D(_01465_),
    .Q(\tms1x00.A[2] ));
 sky130_fd_sc_hd__dfxtp_2 _11665_ (.CLK(clknet_leaf_89_wb_clk_i),
    .D(_01466_),
    .Q(\tms1x00.A[3] ));
 sky130_fd_sc_hd__dfxtp_1 _11666_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_01467_),
    .Q(\tms1x00.O_pla_ands[30][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11667_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_01468_),
    .Q(\tms1x00.O_pla_ands[30][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11668_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_01469_),
    .Q(\tms1x00.O_pla_ands[30][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11669_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_01470_),
    .Q(\tms1x00.O_pla_ands[30][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11670_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_01471_),
    .Q(\tms1x00.O_pla_ands[30][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11671_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_01472_),
    .Q(\tms1x00.O_pla_ands[30][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11672_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_01473_),
    .Q(\tms1x00.O_pla_ands[30][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11673_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_01474_),
    .Q(\tms1x00.O_pla_ands[30][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11674_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_01475_),
    .Q(\tms1x00.O_pla_ands[30][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11675_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_01476_),
    .Q(\tms1x00.O_pla_ands[30][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11676_ (.CLK(clknet_leaf_63_wb_clk_i),
    .D(_01477_),
    .Q(\tms1x00.O_pla_ands[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11677_ (.CLK(clknet_leaf_64_wb_clk_i),
    .D(_01478_),
    .Q(\tms1x00.O_pla_ands[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11678_ (.CLK(clknet_leaf_64_wb_clk_i),
    .D(_01479_),
    .Q(\tms1x00.O_pla_ands[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11679_ (.CLK(clknet_leaf_64_wb_clk_i),
    .D(_01480_),
    .Q(\tms1x00.O_pla_ands[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11680_ (.CLK(clknet_leaf_61_wb_clk_i),
    .D(_01481_),
    .Q(\tms1x00.O_pla_ands[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11681_ (.CLK(clknet_leaf_64_wb_clk_i),
    .D(_01482_),
    .Q(\tms1x00.O_pla_ands[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11682_ (.CLK(clknet_leaf_64_wb_clk_i),
    .D(_01483_),
    .Q(\tms1x00.O_pla_ands[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11683_ (.CLK(clknet_leaf_61_wb_clk_i),
    .D(_01484_),
    .Q(\tms1x00.O_pla_ands[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11684_ (.CLK(clknet_leaf_64_wb_clk_i),
    .D(_01485_),
    .Q(\tms1x00.O_pla_ands[4][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11685_ (.CLK(clknet_leaf_63_wb_clk_i),
    .D(_01486_),
    .Q(\tms1x00.O_pla_ands[4][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11686_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_01487_),
    .Q(\tms1x00.O_pla_ands[29][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11687_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_01488_),
    .Q(\tms1x00.O_pla_ands[29][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11688_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_01489_),
    .Q(\tms1x00.O_pla_ands[29][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11689_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_01490_),
    .Q(\tms1x00.O_pla_ands[29][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11690_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_01491_),
    .Q(\tms1x00.O_pla_ands[29][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11691_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_01492_),
    .Q(\tms1x00.O_pla_ands[29][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11692_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_01493_),
    .Q(\tms1x00.O_pla_ands[29][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11693_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_01494_),
    .Q(\tms1x00.O_pla_ands[29][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11694_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_01495_),
    .Q(\tms1x00.O_pla_ands[29][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11695_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_01496_),
    .Q(\tms1x00.O_pla_ands[29][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11696_ (.CLK(clknet_leaf_123_wb_clk_i),
    .D(_01497_),
    .Q(\tms1x00.ins_pla_ors[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11697_ (.CLK(clknet_leaf_124_wb_clk_i),
    .D(_01498_),
    .Q(\tms1x00.ins_pla_ors[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11698_ (.CLK(clknet_leaf_124_wb_clk_i),
    .D(_01499_),
    .Q(\tms1x00.ins_pla_ors[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11699_ (.CLK(clknet_leaf_126_wb_clk_i),
    .D(_01500_),
    .Q(\tms1x00.ins_pla_ors[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11700_ (.CLK(clknet_leaf_125_wb_clk_i),
    .D(_01501_),
    .Q(\tms1x00.ins_pla_ors[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11701_ (.CLK(clknet_leaf_119_wb_clk_i),
    .D(_01502_),
    .Q(\tms1x00.ins_pla_ors[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11702_ (.CLK(clknet_leaf_126_wb_clk_i),
    .D(_01503_),
    .Q(\tms1x00.ins_pla_ors[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11703_ (.CLK(clknet_leaf_125_wb_clk_i),
    .D(_01504_),
    .Q(\tms1x00.ins_pla_ors[9][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11704_ (.CLK(clknet_leaf_134_wb_clk_i),
    .D(_01505_),
    .Q(\tms1x00.ins_pla_ors[9][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11705_ (.CLK(clknet_leaf_116_wb_clk_i),
    .D(_01506_),
    .Q(\tms1x00.ins_pla_ors[9][10] ));
 sky130_fd_sc_hd__dfxtp_2 _11706_ (.CLK(clknet_leaf_134_wb_clk_i),
    .D(_01507_),
    .Q(\tms1x00.ins_pla_ors[9][11] ));
 sky130_fd_sc_hd__dfxtp_1 _11707_ (.CLK(clknet_leaf_135_wb_clk_i),
    .D(_01508_),
    .Q(\tms1x00.ins_pla_ors[9][12] ));
 sky130_fd_sc_hd__dfxtp_2 _11708_ (.CLK(clknet_leaf_135_wb_clk_i),
    .D(_01509_),
    .Q(\tms1x00.ins_pla_ors[9][13] ));
 sky130_fd_sc_hd__dfxtp_1 _11709_ (.CLK(clknet_leaf_135_wb_clk_i),
    .D(_01510_),
    .Q(\tms1x00.ins_pla_ors[9][14] ));
 sky130_fd_sc_hd__dfxtp_1 _11710_ (.CLK(clknet_leaf_133_wb_clk_i),
    .D(_01511_),
    .Q(\tms1x00.ins_pla_ors[9][15] ));
 sky130_fd_sc_hd__dfxtp_1 _11711_ (.CLK(clknet_leaf_122_wb_clk_i),
    .D(_01512_),
    .Q(\tms1x00.ins_pla_ors[9][16] ));
 sky130_fd_sc_hd__dfxtp_2 _11712_ (.CLK(clknet_leaf_114_wb_clk_i),
    .D(_01513_),
    .Q(\tms1x00.ins_pla_ors[9][17] ));
 sky130_fd_sc_hd__dfxtp_1 _11713_ (.CLK(clknet_leaf_123_wb_clk_i),
    .D(_01514_),
    .Q(\tms1x00.ins_pla_ors[9][18] ));
 sky130_fd_sc_hd__dfxtp_2 _11714_ (.CLK(clknet_leaf_116_wb_clk_i),
    .D(_01515_),
    .Q(\tms1x00.ins_pla_ors[9][19] ));
 sky130_fd_sc_hd__dfxtp_2 _11715_ (.CLK(clknet_leaf_115_wb_clk_i),
    .D(_01516_),
    .Q(\tms1x00.ins_pla_ors[9][20] ));
 sky130_fd_sc_hd__dfxtp_1 _11716_ (.CLK(clknet_leaf_135_wb_clk_i),
    .D(_01517_),
    .Q(\tms1x00.ins_pla_ors[9][21] ));
 sky130_fd_sc_hd__dfxtp_2 _11717_ (.CLK(clknet_leaf_116_wb_clk_i),
    .D(_01518_),
    .Q(\tms1x00.ins_pla_ors[9][22] ));
 sky130_fd_sc_hd__dfxtp_2 _11718_ (.CLK(clknet_leaf_115_wb_clk_i),
    .D(_01519_),
    .Q(\tms1x00.ins_pla_ors[9][23] ));
 sky130_fd_sc_hd__dfxtp_2 _11719_ (.CLK(clknet_leaf_115_wb_clk_i),
    .D(_01520_),
    .Q(\tms1x00.ins_pla_ors[9][24] ));
 sky130_fd_sc_hd__dfxtp_1 _11720_ (.CLK(clknet_leaf_116_wb_clk_i),
    .D(_01521_),
    .Q(\tms1x00.ins_pla_ors[9][25] ));
 sky130_fd_sc_hd__dfxtp_1 _11721_ (.CLK(clknet_leaf_117_wb_clk_i),
    .D(_01522_),
    .Q(\tms1x00.ins_pla_ors[9][26] ));
 sky130_fd_sc_hd__dfxtp_2 _11722_ (.CLK(clknet_leaf_117_wb_clk_i),
    .D(_01523_),
    .Q(\tms1x00.ins_pla_ors[9][28] ));
 sky130_fd_sc_hd__dfxtp_1 _11723_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_01524_),
    .Q(\tms1x00.O_pla_ands[27][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11724_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_01525_),
    .Q(\tms1x00.O_pla_ands[27][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11725_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_01526_),
    .Q(\tms1x00.O_pla_ands[27][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11726_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_01527_),
    .Q(\tms1x00.O_pla_ands[27][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11727_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_01528_),
    .Q(\tms1x00.O_pla_ands[27][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11728_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_01529_),
    .Q(\tms1x00.O_pla_ands[27][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11729_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_01530_),
    .Q(\tms1x00.O_pla_ands[27][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11730_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_01531_),
    .Q(\tms1x00.O_pla_ands[27][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11731_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_01532_),
    .Q(\tms1x00.O_pla_ands[27][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11732_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_01533_),
    .Q(\tms1x00.O_pla_ands[27][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11733_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_01534_),
    .Q(\tms1x00.O_pla_ands[28][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11734_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_01535_),
    .Q(\tms1x00.O_pla_ands[28][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11735_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_01536_),
    .Q(\tms1x00.O_pla_ands[28][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11736_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_01537_),
    .Q(\tms1x00.O_pla_ands[28][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11737_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_01538_),
    .Q(\tms1x00.O_pla_ands[28][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11738_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_01539_),
    .Q(\tms1x00.O_pla_ands[28][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11739_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_01540_),
    .Q(\tms1x00.O_pla_ands[28][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11740_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_01541_),
    .Q(\tms1x00.O_pla_ands[28][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11741_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_01542_),
    .Q(\tms1x00.O_pla_ands[28][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11742_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_01543_),
    .Q(\tms1x00.O_pla_ands[28][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11743_ (.CLK(clknet_leaf_132_wb_clk_i),
    .D(_01544_),
    .Q(\tms1x00.ins_pla_ors[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11744_ (.CLK(clknet_leaf_119_wb_clk_i),
    .D(_01545_),
    .Q(\tms1x00.ins_pla_ors[9][27] ));
 sky130_fd_sc_hd__dfxtp_1 _11745_ (.CLK(clknet_leaf_120_wb_clk_i),
    .D(_01546_),
    .Q(\tms1x00.ins_pla_ors[9][29] ));
 sky130_fd_sc_hd__dfxtp_1 _11746_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(_01547_),
    .Q(\tms1x00.O_pla_ands[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11747_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_01548_),
    .Q(\tms1x00.O_pla_ands[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11748_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(_01549_),
    .Q(\tms1x00.O_pla_ands[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11749_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_01550_),
    .Q(\tms1x00.O_pla_ands[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11750_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_01551_),
    .Q(\tms1x00.O_pla_ands[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11751_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_01552_),
    .Q(\tms1x00.O_pla_ands[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11752_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(_01553_),
    .Q(\tms1x00.O_pla_ands[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11753_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_01554_),
    .Q(\tms1x00.O_pla_ands[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11754_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_01555_),
    .Q(\tms1x00.O_pla_ands[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11755_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(_01556_),
    .Q(\tms1x00.O_pla_ands[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11756_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_01557_),
    .Q(\tms1x00.O_pla_ands[24][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11757_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_01558_),
    .Q(\tms1x00.O_pla_ands[24][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11758_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_01559_),
    .Q(\tms1x00.O_pla_ands[24][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11759_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_01560_),
    .Q(\tms1x00.O_pla_ands[24][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11760_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_01561_),
    .Q(\tms1x00.O_pla_ands[24][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11761_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_01562_),
    .Q(\tms1x00.O_pla_ands[24][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11762_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_01563_),
    .Q(\tms1x00.O_pla_ands[24][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11763_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_01564_),
    .Q(\tms1x00.O_pla_ands[24][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11764_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_01565_),
    .Q(\tms1x00.O_pla_ands[24][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11765_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_01566_),
    .Q(\tms1x00.O_pla_ands[24][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11766_ (.CLK(clknet_leaf_130_wb_clk_i),
    .D(_01567_),
    .Q(\tms1x00.ins_pla_ands[31][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11767_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_01568_),
    .Q(\tms1x00.ins_pla_ands[31][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11768_ (.CLK(clknet_leaf_139_wb_clk_i),
    .D(_01569_),
    .Q(\tms1x00.ins_pla_ands[31][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11769_ (.CLK(clknet_leaf_143_wb_clk_i),
    .D(_01570_),
    .Q(\tms1x00.ins_pla_ands[31][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11770_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_01571_),
    .Q(\tms1x00.ins_pla_ands[31][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11771_ (.CLK(clknet_leaf_138_wb_clk_i),
    .D(_01572_),
    .Q(\tms1x00.ins_pla_ands[31][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11772_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_01573_),
    .Q(\tms1x00.ins_pla_ands[31][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11773_ (.CLK(clknet_leaf_142_wb_clk_i),
    .D(_01574_),
    .Q(\tms1x00.ins_pla_ands[31][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11774_ (.CLK(clknet_leaf_143_wb_clk_i),
    .D(_01575_),
    .Q(\tms1x00.ins_pla_ands[31][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11775_ (.CLK(clknet_leaf_143_wb_clk_i),
    .D(_01576_),
    .Q(\tms1x00.ins_pla_ands[31][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11776_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_01577_),
    .Q(\tms1x00.ins_pla_ands[31][10] ));
 sky130_fd_sc_hd__dfxtp_1 _11777_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_01578_),
    .Q(\tms1x00.ins_pla_ands[31][11] ));
 sky130_fd_sc_hd__dfxtp_1 _11778_ (.CLK(clknet_leaf_143_wb_clk_i),
    .D(_01579_),
    .Q(\tms1x00.ins_pla_ands[31][12] ));
 sky130_fd_sc_hd__dfxtp_1 _11779_ (.CLK(clknet_leaf_143_wb_clk_i),
    .D(_01580_),
    .Q(\tms1x00.ins_pla_ands[31][13] ));
 sky130_fd_sc_hd__dfxtp_1 _11780_ (.CLK(clknet_leaf_138_wb_clk_i),
    .D(_01581_),
    .Q(\tms1x00.ins_pla_ands[31][14] ));
 sky130_fd_sc_hd__dfxtp_1 _11781_ (.CLK(clknet_leaf_142_wb_clk_i),
    .D(_01582_),
    .Q(\tms1x00.ins_pla_ands[31][15] ));
 sky130_fd_sc_hd__dfxtp_1 _11782_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_01583_),
    .Q(\tms1x00.O_pla_ands[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11783_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_01584_),
    .Q(\tms1x00.O_pla_ands[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11784_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_01585_),
    .Q(\tms1x00.O_pla_ands[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11785_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_01586_),
    .Q(\tms1x00.O_pla_ands[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11786_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_01587_),
    .Q(\tms1x00.O_pla_ands[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11787_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_01588_),
    .Q(\tms1x00.O_pla_ands[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11788_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_01589_),
    .Q(\tms1x00.O_pla_ands[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11789_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_01590_),
    .Q(\tms1x00.O_pla_ands[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11790_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_01591_),
    .Q(\tms1x00.O_pla_ands[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11791_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_01592_),
    .Q(\tms1x00.O_pla_ands[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11792_ (.CLK(clknet_leaf_67_wb_clk_i),
    .D(_01593_),
    .Q(\tms1x00.O_pla_ands[3][0] ));
 sky130_fd_sc_hd__dfxtp_2 _11793_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_01594_),
    .Q(\tms1x00.O_pla_ands[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11794_ (.CLK(clknet_leaf_65_wb_clk_i),
    .D(_01595_),
    .Q(\tms1x00.O_pla_ands[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11795_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_01596_),
    .Q(\tms1x00.O_pla_ands[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11796_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_01597_),
    .Q(\tms1x00.O_pla_ands[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11797_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_01598_),
    .Q(\tms1x00.O_pla_ands[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11798_ (.CLK(clknet_leaf_65_wb_clk_i),
    .D(_01599_),
    .Q(\tms1x00.O_pla_ands[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11799_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_01600_),
    .Q(\tms1x00.O_pla_ands[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11800_ (.CLK(clknet_leaf_65_wb_clk_i),
    .D(_01601_),
    .Q(\tms1x00.O_pla_ands[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11801_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_01602_),
    .Q(\tms1x00.O_pla_ands[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11802_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_01603_),
    .Q(\tms1x00.O_pla_ands[21][0] ));
 sky130_fd_sc_hd__dfxtp_1 _11803_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_01604_),
    .Q(\tms1x00.O_pla_ands[21][1] ));
 sky130_fd_sc_hd__dfxtp_1 _11804_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(_01605_),
    .Q(\tms1x00.O_pla_ands[21][2] ));
 sky130_fd_sc_hd__dfxtp_1 _11805_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_01606_),
    .Q(\tms1x00.O_pla_ands[21][3] ));
 sky130_fd_sc_hd__dfxtp_1 _11806_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_01607_),
    .Q(\tms1x00.O_pla_ands[21][4] ));
 sky130_fd_sc_hd__dfxtp_1 _11807_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_01608_),
    .Q(\tms1x00.O_pla_ands[21][5] ));
 sky130_fd_sc_hd__dfxtp_1 _11808_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_01609_),
    .Q(\tms1x00.O_pla_ands[21][6] ));
 sky130_fd_sc_hd__dfxtp_1 _11809_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_01610_),
    .Q(\tms1x00.O_pla_ands[21][7] ));
 sky130_fd_sc_hd__dfxtp_1 _11810_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(_01611_),
    .Q(\tms1x00.O_pla_ands[21][8] ));
 sky130_fd_sc_hd__dfxtp_1 _11811_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(_01612_),
    .Q(\tms1x00.O_pla_ands[21][9] ));
 sky130_fd_sc_hd__dfxtp_4 _11812_ (.CLK(clknet_leaf_86_wb_clk_i),
    .D(_01613_),
    .Q(net128));
 sky130_fd_sc_hd__buf_2 _11866_ (.A(net79),
    .X(net168));
 sky130_fd_sc_hd__buf_2 _11867_ (.A(net1004),
    .X(net169));
 sky130_fd_sc_hd__buf_2 _11868_ (.A(net1002),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_2 _11869_ (.A(net991),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_2 _11870_ (.A(net989),
    .X(net172));
 sky130_fd_sc_hd__buf_2 _11871_ (.A(net985),
    .X(net173));
 sky130_fd_sc_hd__buf_2 _11872_ (.A(net984),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_2 _11873_ (.A(net86),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_2 _11874_ (.A(net75),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_0_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_0_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_1_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_1_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_2_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_2_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_3_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_3_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_4_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_4_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_5_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_5_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_6_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_6_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_7_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_7_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_0__f_wb_clk_i (.A(clknet_3_0_0_wb_clk_i),
    .X(clknet_4_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_10__f_wb_clk_i (.A(clknet_3_5_0_wb_clk_i),
    .X(clknet_4_10__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_11__f_wb_clk_i (.A(clknet_3_5_0_wb_clk_i),
    .X(clknet_4_11__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_12__f_wb_clk_i (.A(clknet_3_6_0_wb_clk_i),
    .X(clknet_4_12__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_13__f_wb_clk_i (.A(clknet_3_6_0_wb_clk_i),
    .X(clknet_4_13__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_14__f_wb_clk_i (.A(clknet_3_7_0_wb_clk_i),
    .X(clknet_4_14__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_15__f_wb_clk_i (.A(clknet_3_7_0_wb_clk_i),
    .X(clknet_4_15__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_1__f_wb_clk_i (.A(clknet_3_0_0_wb_clk_i),
    .X(clknet_4_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_2__f_wb_clk_i (.A(clknet_3_1_0_wb_clk_i),
    .X(clknet_4_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_3__f_wb_clk_i (.A(clknet_3_1_0_wb_clk_i),
    .X(clknet_4_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_4__f_wb_clk_i (.A(clknet_3_2_0_wb_clk_i),
    .X(clknet_4_4__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_5__f_wb_clk_i (.A(clknet_3_2_0_wb_clk_i),
    .X(clknet_4_5__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_6__f_wb_clk_i (.A(clknet_3_3_0_wb_clk_i),
    .X(clknet_4_6__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_7__f_wb_clk_i (.A(clknet_3_3_0_wb_clk_i),
    .X(clknet_4_7__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_8__f_wb_clk_i (.A(clknet_3_4_0_wb_clk_i),
    .X(clknet_4_8__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_9__f_wb_clk_i (.A(clknet_3_4_0_wb_clk_i),
    .X(clknet_4_9__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_wb_clk_i (.A(clknet_4_0__leaf_wb_clk_i),
    .X(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_100_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .X(clknet_leaf_100_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_101_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .X(clknet_leaf_101_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_102_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .X(clknet_leaf_102_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_103_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .X(clknet_leaf_103_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_104_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .X(clknet_leaf_104_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_105_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .X(clknet_leaf_105_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_106_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .X(clknet_leaf_106_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_107_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .X(clknet_leaf_107_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_108_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .X(clknet_leaf_108_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_109_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .X(clknet_leaf_109_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .X(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_110_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .X(clknet_leaf_110_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_111_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .X(clknet_leaf_111_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_112_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_112_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_113_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_113_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_114_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_114_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_115_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_115_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_116_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_116_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_117_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_117_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_118_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_118_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_119_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_119_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .X(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_120_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_120_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_121_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_121_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_122_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .X(clknet_leaf_122_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_123_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .X(clknet_leaf_123_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_124_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .X(clknet_leaf_124_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_125_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .X(clknet_leaf_125_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_126_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .X(clknet_leaf_126_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_127_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .X(clknet_leaf_127_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_128_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .X(clknet_leaf_128_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_129_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .X(clknet_leaf_129_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .X(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_130_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .X(clknet_leaf_130_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_131_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .X(clknet_leaf_131_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_132_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .X(clknet_leaf_132_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_133_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .X(clknet_leaf_133_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_134_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .X(clknet_leaf_134_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_135_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .X(clknet_leaf_135_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_136_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .X(clknet_leaf_136_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_137_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .X(clknet_leaf_137_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_138_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .X(clknet_leaf_138_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_139_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .X(clknet_leaf_139_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .X(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_140_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .X(clknet_leaf_140_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_141_wb_clk_i (.A(clknet_4_0__leaf_wb_clk_i),
    .X(clknet_leaf_141_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_142_wb_clk_i (.A(clknet_4_0__leaf_wb_clk_i),
    .X(clknet_leaf_142_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_143_wb_clk_i (.A(clknet_4_0__leaf_wb_clk_i),
    .X(clknet_leaf_143_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_wb_clk_i (.A(clknet_4_0__leaf_wb_clk_i),
    .X(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .X(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .X(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .X(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .X(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .X(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_wb_clk_i (.A(clknet_4_0__leaf_wb_clk_i),
    .X(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .X(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .X(clknet_leaf_21_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .X(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_wb_clk_i (.A(clknet_4_4__leaf_wb_clk_i),
    .X(clknet_leaf_23_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_wb_clk_i (.A(clknet_4_4__leaf_wb_clk_i),
    .X(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_wb_clk_i (.A(clknet_4_4__leaf_wb_clk_i),
    .X(clknet_leaf_25_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_wb_clk_i (.A(clknet_4_4__leaf_wb_clk_i),
    .X(clknet_leaf_26_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_wb_clk_i (.A(clknet_4_4__leaf_wb_clk_i),
    .X(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_wb_clk_i (.A(clknet_4_4__leaf_wb_clk_i),
    .X(clknet_leaf_28_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_wb_clk_i (.A(clknet_4_4__leaf_wb_clk_i),
    .X(clknet_leaf_29_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_wb_clk_i (.A(clknet_4_0__leaf_wb_clk_i),
    .X(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_wb_clk_i (.A(clknet_4_4__leaf_wb_clk_i),
    .X(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_wb_clk_i (.A(clknet_4_4__leaf_wb_clk_i),
    .X(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .X(clknet_leaf_32_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .X(clknet_leaf_33_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .X(clknet_leaf_34_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .X(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .X(clknet_leaf_36_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .X(clknet_leaf_37_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .X(clknet_leaf_38_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .X(clknet_leaf_39_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_wb_clk_i (.A(clknet_4_0__leaf_wb_clk_i),
    .X(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .X(clknet_leaf_40_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .X(clknet_leaf_41_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .X(clknet_leaf_42_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .X(clknet_leaf_43_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .X(clknet_leaf_44_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .X(clknet_leaf_45_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .X(clknet_leaf_46_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .X(clknet_leaf_47_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .X(clknet_leaf_48_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .X(clknet_leaf_49_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .X(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .X(clknet_leaf_50_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .X(clknet_leaf_51_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .X(clknet_leaf_52_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .X(clknet_leaf_53_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .X(clknet_leaf_54_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .X(clknet_leaf_55_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .X(clknet_leaf_56_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .X(clknet_leaf_57_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .X(clknet_leaf_58_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .X(clknet_leaf_59_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .X(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .X(clknet_leaf_60_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_61_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_62_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_63_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_64_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_65_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_66_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_67_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_68_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_69_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .X(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .X(clknet_leaf_70_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .X(clknet_leaf_71_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .X(clknet_leaf_72_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .X(clknet_leaf_73_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .X(clknet_leaf_74_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .X(clknet_leaf_75_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .X(clknet_leaf_76_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .X(clknet_leaf_77_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .X(clknet_leaf_78_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .X(clknet_leaf_79_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .X(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .X(clknet_leaf_80_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .X(clknet_leaf_81_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .X(clknet_leaf_82_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .X(clknet_leaf_83_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .X(clknet_leaf_84_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .X(clknet_leaf_85_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .X(clknet_leaf_86_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .X(clknet_leaf_87_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .X(clknet_leaf_88_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .X(clknet_leaf_89_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .X(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .X(clknet_leaf_90_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .X(clknet_leaf_91_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .X(clknet_leaf_92_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .X(clknet_leaf_93_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .X(clknet_leaf_94_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .X(clknet_leaf_95_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .X(clknet_leaf_96_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_97_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .X(clknet_leaf_97_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_98_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .X(clknet_leaf_98_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_99_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .X(clknet_leaf_99_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .X(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 fanout1000 (.A(net82),
    .X(net1000));
 sky130_fd_sc_hd__clkbuf_8 fanout1001 (.A(net1002),
    .X(net1001));
 sky130_fd_sc_hd__buf_6 fanout1002 (.A(net81),
    .X(net1002));
 sky130_fd_sc_hd__buf_6 fanout1003 (.A(net1004),
    .X(net1003));
 sky130_fd_sc_hd__buf_4 fanout1004 (.A(net80),
    .X(net1004));
 sky130_fd_sc_hd__buf_8 fanout1005 (.A(net79),
    .X(net1005));
 sky130_fd_sc_hd__clkbuf_4 fanout1006 (.A(net79),
    .X(net1006));
 sky130_fd_sc_hd__buf_4 fanout1007 (.A(net1008),
    .X(net1007));
 sky130_fd_sc_hd__buf_6 fanout1008 (.A(net1009),
    .X(net1008));
 sky130_fd_sc_hd__clkbuf_16 fanout1009 (.A(net1010),
    .X(net1009));
 sky130_fd_sc_hd__buf_12 fanout1010 (.A(net117),
    .X(net1010));
 sky130_fd_sc_hd__buf_6 fanout1011 (.A(net1012),
    .X(net1011));
 sky130_fd_sc_hd__clkbuf_16 fanout1012 (.A(net1013),
    .X(net1012));
 sky130_fd_sc_hd__buf_12 fanout1013 (.A(net117),
    .X(net1013));
 sky130_fd_sc_hd__buf_6 fanout1014 (.A(net1018),
    .X(net1014));
 sky130_fd_sc_hd__buf_4 fanout1015 (.A(net1017),
    .X(net1015));
 sky130_fd_sc_hd__buf_2 fanout1016 (.A(net1017),
    .X(net1016));
 sky130_fd_sc_hd__buf_6 fanout1017 (.A(net1018),
    .X(net1017));
 sky130_fd_sc_hd__buf_12 fanout1018 (.A(net1023),
    .X(net1018));
 sky130_fd_sc_hd__buf_6 fanout1019 (.A(net1023),
    .X(net1019));
 sky130_fd_sc_hd__buf_6 fanout1020 (.A(net1021),
    .X(net1020));
 sky130_fd_sc_hd__clkbuf_8 fanout1021 (.A(net1023),
    .X(net1021));
 sky130_fd_sc_hd__buf_6 fanout1022 (.A(net1023),
    .X(net1022));
 sky130_fd_sc_hd__buf_12 fanout1023 (.A(net116),
    .X(net1023));
 sky130_fd_sc_hd__buf_4 fanout1024 (.A(net1026),
    .X(net1024));
 sky130_fd_sc_hd__buf_6 fanout1025 (.A(net1026),
    .X(net1025));
 sky130_fd_sc_hd__buf_12 fanout1026 (.A(net115),
    .X(net1026));
 sky130_fd_sc_hd__buf_6 fanout1027 (.A(net1028),
    .X(net1027));
 sky130_fd_sc_hd__buf_8 fanout1028 (.A(net1029),
    .X(net1028));
 sky130_fd_sc_hd__buf_12 fanout1029 (.A(net115),
    .X(net1029));
 sky130_fd_sc_hd__buf_4 fanout1030 (.A(net1032),
    .X(net1030));
 sky130_fd_sc_hd__buf_6 fanout1031 (.A(net1032),
    .X(net1031));
 sky130_fd_sc_hd__buf_6 fanout1032 (.A(net114),
    .X(net1032));
 sky130_fd_sc_hd__buf_6 fanout1033 (.A(net114),
    .X(net1033));
 sky130_fd_sc_hd__buf_6 fanout1034 (.A(net1035),
    .X(net1034));
 sky130_fd_sc_hd__buf_4 fanout1035 (.A(net1036),
    .X(net1035));
 sky130_fd_sc_hd__buf_6 fanout1036 (.A(net1037),
    .X(net1036));
 sky130_fd_sc_hd__buf_12 fanout1037 (.A(net114),
    .X(net1037));
 sky130_fd_sc_hd__buf_4 fanout1038 (.A(net1039),
    .X(net1038));
 sky130_fd_sc_hd__clkbuf_8 fanout1039 (.A(net1045),
    .X(net1039));
 sky130_fd_sc_hd__buf_8 fanout1040 (.A(net1045),
    .X(net1040));
 sky130_fd_sc_hd__buf_12 fanout1041 (.A(net1045),
    .X(net1041));
 sky130_fd_sc_hd__buf_6 fanout1042 (.A(net1044),
    .X(net1042));
 sky130_fd_sc_hd__buf_6 fanout1043 (.A(net1044),
    .X(net1043));
 sky130_fd_sc_hd__buf_12 fanout1044 (.A(net1045),
    .X(net1044));
 sky130_fd_sc_hd__buf_12 fanout1045 (.A(net113),
    .X(net1045));
 sky130_fd_sc_hd__buf_4 fanout1046 (.A(net1047),
    .X(net1046));
 sky130_fd_sc_hd__buf_4 fanout1047 (.A(net1048),
    .X(net1047));
 sky130_fd_sc_hd__buf_6 fanout1048 (.A(net1049),
    .X(net1048));
 sky130_fd_sc_hd__clkbuf_16 fanout1049 (.A(net112),
    .X(net1049));
 sky130_fd_sc_hd__buf_6 fanout1050 (.A(net1052),
    .X(net1050));
 sky130_fd_sc_hd__buf_4 fanout1051 (.A(net1052),
    .X(net1051));
 sky130_fd_sc_hd__buf_8 fanout1052 (.A(net112),
    .X(net1052));
 sky130_fd_sc_hd__buf_6 fanout1053 (.A(net112),
    .X(net1053));
 sky130_fd_sc_hd__clkbuf_4 fanout1054 (.A(net1055),
    .X(net1054));
 sky130_fd_sc_hd__clkbuf_8 fanout1055 (.A(net1057),
    .X(net1055));
 sky130_fd_sc_hd__buf_6 fanout1056 (.A(net1057),
    .X(net1056));
 sky130_fd_sc_hd__buf_6 fanout1057 (.A(net1058),
    .X(net1057));
 sky130_fd_sc_hd__buf_12 fanout1058 (.A(net111),
    .X(net1058));
 sky130_fd_sc_hd__buf_6 fanout1059 (.A(net1061),
    .X(net1059));
 sky130_fd_sc_hd__buf_6 fanout1060 (.A(net1061),
    .X(net1060));
 sky130_fd_sc_hd__buf_8 fanout1061 (.A(net1062),
    .X(net1061));
 sky130_fd_sc_hd__buf_6 fanout1062 (.A(net111),
    .X(net1062));
 sky130_fd_sc_hd__buf_4 fanout1063 (.A(net1065),
    .X(net1063));
 sky130_fd_sc_hd__buf_2 fanout1064 (.A(net1065),
    .X(net1064));
 sky130_fd_sc_hd__buf_4 fanout1065 (.A(net1071),
    .X(net1065));
 sky130_fd_sc_hd__buf_12 fanout1066 (.A(net1071),
    .X(net1066));
 sky130_fd_sc_hd__buf_6 fanout1067 (.A(net1069),
    .X(net1067));
 sky130_fd_sc_hd__buf_6 fanout1068 (.A(net1069),
    .X(net1068));
 sky130_fd_sc_hd__buf_6 fanout1069 (.A(net1071),
    .X(net1069));
 sky130_fd_sc_hd__buf_6 fanout1070 (.A(net1071),
    .X(net1070));
 sky130_fd_sc_hd__buf_12 fanout1071 (.A(net110),
    .X(net1071));
 sky130_fd_sc_hd__buf_6 fanout1072 (.A(net106),
    .X(net1072));
 sky130_fd_sc_hd__buf_8 fanout1073 (.A(net104),
    .X(net1073));
 sky130_fd_sc_hd__buf_8 fanout1074 (.A(net103),
    .X(net1074));
 sky130_fd_sc_hd__buf_6 fanout1075 (.A(net102),
    .X(net1075));
 sky130_fd_sc_hd__clkbuf_2 fanout1076 (.A(net102),
    .X(net1076));
 sky130_fd_sc_hd__buf_6 fanout1077 (.A(net101),
    .X(net1077));
 sky130_fd_sc_hd__buf_6 fanout1078 (.A(net100),
    .X(net1078));
 sky130_fd_sc_hd__clkbuf_4 fanout1079 (.A(net100),
    .X(net1079));
 sky130_fd_sc_hd__buf_6 fanout212 (.A(net215),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_4 fanout213 (.A(net215),
    .X(net213));
 sky130_fd_sc_hd__buf_6 fanout214 (.A(net215),
    .X(net214));
 sky130_fd_sc_hd__buf_6 fanout215 (.A(_03791_),
    .X(net215));
 sky130_fd_sc_hd__buf_4 fanout216 (.A(_03715_),
    .X(net216));
 sky130_fd_sc_hd__buf_2 fanout217 (.A(_03715_),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_8 fanout218 (.A(_03594_),
    .X(net218));
 sky130_fd_sc_hd__buf_2 fanout219 (.A(_03594_),
    .X(net219));
 sky130_fd_sc_hd__buf_6 fanout220 (.A(net221),
    .X(net220));
 sky130_fd_sc_hd__clkbuf_4 fanout221 (.A(_03591_),
    .X(net221));
 sky130_fd_sc_hd__buf_6 fanout222 (.A(net224),
    .X(net222));
 sky130_fd_sc_hd__buf_8 fanout223 (.A(net224),
    .X(net223));
 sky130_fd_sc_hd__buf_12 fanout224 (.A(_03532_),
    .X(net224));
 sky130_fd_sc_hd__buf_6 fanout225 (.A(_03529_),
    .X(net225));
 sky130_fd_sc_hd__buf_4 fanout226 (.A(_03529_),
    .X(net226));
 sky130_fd_sc_hd__buf_8 fanout227 (.A(_03528_),
    .X(net227));
 sky130_fd_sc_hd__buf_6 fanout228 (.A(net230),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_2 fanout229 (.A(net230),
    .X(net229));
 sky130_fd_sc_hd__buf_8 fanout230 (.A(_03490_),
    .X(net230));
 sky130_fd_sc_hd__buf_6 fanout231 (.A(net233),
    .X(net231));
 sky130_fd_sc_hd__buf_6 fanout232 (.A(net233),
    .X(net232));
 sky130_fd_sc_hd__buf_6 fanout233 (.A(_03455_),
    .X(net233));
 sky130_fd_sc_hd__buf_8 fanout234 (.A(_03423_),
    .X(net234));
 sky130_fd_sc_hd__buf_6 fanout235 (.A(_05045_),
    .X(net235));
 sky130_fd_sc_hd__buf_4 fanout236 (.A(_05045_),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_16 fanout237 (.A(_05006_),
    .X(net237));
 sky130_fd_sc_hd__buf_6 fanout238 (.A(_05005_),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_4 fanout239 (.A(_05005_),
    .X(net239));
 sky130_fd_sc_hd__buf_4 fanout240 (.A(_04574_),
    .X(net240));
 sky130_fd_sc_hd__buf_2 fanout241 (.A(_04574_),
    .X(net241));
 sky130_fd_sc_hd__buf_4 fanout242 (.A(_04571_),
    .X(net242));
 sky130_fd_sc_hd__buf_2 fanout243 (.A(_04571_),
    .X(net243));
 sky130_fd_sc_hd__buf_4 fanout244 (.A(net245),
    .X(net244));
 sky130_fd_sc_hd__buf_6 fanout245 (.A(_04282_),
    .X(net245));
 sky130_fd_sc_hd__clkbuf_4 fanout246 (.A(net247),
    .X(net246));
 sky130_fd_sc_hd__buf_4 fanout247 (.A(_04281_),
    .X(net247));
 sky130_fd_sc_hd__buf_6 fanout248 (.A(net250),
    .X(net248));
 sky130_fd_sc_hd__buf_2 fanout249 (.A(net250),
    .X(net249));
 sky130_fd_sc_hd__buf_6 fanout250 (.A(_04258_),
    .X(net250));
 sky130_fd_sc_hd__buf_6 fanout251 (.A(_04214_),
    .X(net251));
 sky130_fd_sc_hd__buf_6 fanout252 (.A(_04214_),
    .X(net252));
 sky130_fd_sc_hd__buf_6 fanout253 (.A(net254),
    .X(net253));
 sky130_fd_sc_hd__buf_8 fanout254 (.A(_04167_),
    .X(net254));
 sky130_fd_sc_hd__buf_6 fanout255 (.A(_04157_),
    .X(net255));
 sky130_fd_sc_hd__clkbuf_4 fanout256 (.A(_04157_),
    .X(net256));
 sky130_fd_sc_hd__buf_6 fanout257 (.A(_04130_),
    .X(net257));
 sky130_fd_sc_hd__buf_6 fanout258 (.A(_04130_),
    .X(net258));
 sky130_fd_sc_hd__buf_6 fanout259 (.A(_04113_),
    .X(net259));
 sky130_fd_sc_hd__buf_6 fanout260 (.A(net261),
    .X(net260));
 sky130_fd_sc_hd__buf_8 fanout261 (.A(_04091_),
    .X(net261));
 sky130_fd_sc_hd__buf_4 fanout262 (.A(_04073_),
    .X(net262));
 sky130_fd_sc_hd__buf_2 fanout263 (.A(_04073_),
    .X(net263));
 sky130_fd_sc_hd__buf_6 fanout264 (.A(net265),
    .X(net264));
 sky130_fd_sc_hd__clkbuf_16 fanout265 (.A(_04038_),
    .X(net265));
 sky130_fd_sc_hd__buf_6 fanout266 (.A(_04028_),
    .X(net266));
 sky130_fd_sc_hd__buf_6 fanout267 (.A(_04003_),
    .X(net267));
 sky130_fd_sc_hd__buf_6 fanout268 (.A(net269),
    .X(net268));
 sky130_fd_sc_hd__buf_8 fanout269 (.A(_03978_),
    .X(net269));
 sky130_fd_sc_hd__clkbuf_8 fanout270 (.A(_03953_),
    .X(net270));
 sky130_fd_sc_hd__clkbuf_4 fanout271 (.A(_03953_),
    .X(net271));
 sky130_fd_sc_hd__buf_6 fanout272 (.A(_03945_),
    .X(net272));
 sky130_fd_sc_hd__buf_4 fanout273 (.A(_03945_),
    .X(net273));
 sky130_fd_sc_hd__buf_4 fanout274 (.A(net275),
    .X(net274));
 sky130_fd_sc_hd__buf_4 fanout275 (.A(_03923_),
    .X(net275));
 sky130_fd_sc_hd__clkbuf_8 fanout276 (.A(_03912_),
    .X(net276));
 sky130_fd_sc_hd__clkbuf_4 fanout277 (.A(_03912_),
    .X(net277));
 sky130_fd_sc_hd__buf_6 fanout278 (.A(_03860_),
    .X(net278));
 sky130_fd_sc_hd__clkbuf_4 fanout279 (.A(_03860_),
    .X(net279));
 sky130_fd_sc_hd__buf_8 fanout280 (.A(net282),
    .X(net280));
 sky130_fd_sc_hd__buf_8 fanout281 (.A(net282),
    .X(net281));
 sky130_fd_sc_hd__buf_6 fanout282 (.A(_03822_),
    .X(net282));
 sky130_fd_sc_hd__buf_6 fanout283 (.A(net286),
    .X(net283));
 sky130_fd_sc_hd__buf_6 fanout284 (.A(net286),
    .X(net284));
 sky130_fd_sc_hd__clkbuf_4 fanout285 (.A(net286),
    .X(net285));
 sky130_fd_sc_hd__clkbuf_8 fanout286 (.A(_03796_),
    .X(net286));
 sky130_fd_sc_hd__buf_4 fanout287 (.A(net289),
    .X(net287));
 sky130_fd_sc_hd__buf_4 fanout288 (.A(net289),
    .X(net288));
 sky130_fd_sc_hd__buf_4 fanout289 (.A(_03795_),
    .X(net289));
 sky130_fd_sc_hd__buf_6 fanout290 (.A(_03793_),
    .X(net290));
 sky130_fd_sc_hd__buf_6 fanout291 (.A(net292),
    .X(net291));
 sky130_fd_sc_hd__buf_8 fanout292 (.A(_03790_),
    .X(net292));
 sky130_fd_sc_hd__buf_8 fanout293 (.A(net295),
    .X(net293));
 sky130_fd_sc_hd__buf_8 fanout294 (.A(net295),
    .X(net294));
 sky130_fd_sc_hd__buf_8 fanout295 (.A(_03769_),
    .X(net295));
 sky130_fd_sc_hd__buf_6 fanout296 (.A(_03721_),
    .X(net296));
 sky130_fd_sc_hd__buf_6 fanout297 (.A(net298),
    .X(net297));
 sky130_fd_sc_hd__buf_6 fanout298 (.A(_03719_),
    .X(net298));
 sky130_fd_sc_hd__clkbuf_8 fanout299 (.A(_03716_),
    .X(net299));
 sky130_fd_sc_hd__buf_4 fanout300 (.A(_03714_),
    .X(net300));
 sky130_fd_sc_hd__buf_6 fanout301 (.A(_03709_),
    .X(net301));
 sky130_fd_sc_hd__buf_8 fanout302 (.A(net305),
    .X(net302));
 sky130_fd_sc_hd__buf_6 fanout303 (.A(net305),
    .X(net303));
 sky130_fd_sc_hd__buf_6 fanout304 (.A(net305),
    .X(net304));
 sky130_fd_sc_hd__buf_6 fanout305 (.A(_03674_),
    .X(net305));
 sky130_fd_sc_hd__clkbuf_8 fanout306 (.A(net307),
    .X(net306));
 sky130_fd_sc_hd__buf_6 fanout307 (.A(_03638_),
    .X(net307));
 sky130_fd_sc_hd__buf_6 fanout308 (.A(_03638_),
    .X(net308));
 sky130_fd_sc_hd__buf_4 fanout309 (.A(net310),
    .X(net309));
 sky130_fd_sc_hd__clkbuf_8 fanout310 (.A(_03637_),
    .X(net310));
 sky130_fd_sc_hd__buf_6 fanout311 (.A(_03637_),
    .X(net311));
 sky130_fd_sc_hd__buf_6 fanout312 (.A(net313),
    .X(net312));
 sky130_fd_sc_hd__buf_6 fanout313 (.A(net314),
    .X(net313));
 sky130_fd_sc_hd__buf_8 fanout314 (.A(_03632_),
    .X(net314));
 sky130_fd_sc_hd__buf_12 fanout315 (.A(_03600_),
    .X(net315));
 sky130_fd_sc_hd__buf_6 fanout316 (.A(_03597_),
    .X(net316));
 sky130_fd_sc_hd__buf_8 fanout317 (.A(_03595_),
    .X(net317));
 sky130_fd_sc_hd__buf_6 fanout318 (.A(_03593_),
    .X(net318));
 sky130_fd_sc_hd__buf_6 fanout319 (.A(_03590_),
    .X(net319));
 sky130_fd_sc_hd__buf_6 fanout320 (.A(_03546_),
    .X(net320));
 sky130_fd_sc_hd__buf_8 fanout321 (.A(_03546_),
    .X(net321));
 sky130_fd_sc_hd__clkbuf_4 fanout322 (.A(_03546_),
    .X(net322));
 sky130_fd_sc_hd__buf_8 fanout323 (.A(_03531_),
    .X(net323));
 sky130_fd_sc_hd__buf_6 fanout324 (.A(_03531_),
    .X(net324));
 sky130_fd_sc_hd__buf_12 fanout325 (.A(_03526_),
    .X(net325));
 sky130_fd_sc_hd__clkbuf_4 fanout326 (.A(_03526_),
    .X(net326));
 sky130_fd_sc_hd__buf_8 fanout327 (.A(net329),
    .X(net327));
 sky130_fd_sc_hd__buf_8 fanout328 (.A(net329),
    .X(net328));
 sky130_fd_sc_hd__buf_8 fanout329 (.A(_03522_),
    .X(net329));
 sky130_fd_sc_hd__buf_6 fanout330 (.A(net331),
    .X(net330));
 sky130_fd_sc_hd__buf_8 fanout331 (.A(_03503_),
    .X(net331));
 sky130_fd_sc_hd__buf_6 fanout332 (.A(net335),
    .X(net332));
 sky130_fd_sc_hd__clkbuf_4 fanout333 (.A(net335),
    .X(net333));
 sky130_fd_sc_hd__buf_4 fanout334 (.A(net335),
    .X(net334));
 sky130_fd_sc_hd__clkbuf_8 fanout335 (.A(_03488_),
    .X(net335));
 sky130_fd_sc_hd__buf_6 fanout336 (.A(_03453_),
    .X(net336));
 sky130_fd_sc_hd__buf_6 fanout337 (.A(_03453_),
    .X(net337));
 sky130_fd_sc_hd__buf_8 fanout338 (.A(_03421_),
    .X(net338));
 sky130_fd_sc_hd__buf_8 fanout339 (.A(_04528_),
    .X(net339));
 sky130_fd_sc_hd__clkbuf_16 fanout340 (.A(_04306_),
    .X(net340));
 sky130_fd_sc_hd__buf_12 fanout341 (.A(net342),
    .X(net341));
 sky130_fd_sc_hd__buf_6 fanout342 (.A(_03976_),
    .X(net342));
 sky130_fd_sc_hd__buf_12 fanout343 (.A(_03585_),
    .X(net343));
 sky130_fd_sc_hd__buf_12 fanout344 (.A(_03533_),
    .X(net344));
 sky130_fd_sc_hd__buf_8 fanout345 (.A(_03501_),
    .X(net345));
 sky130_fd_sc_hd__buf_6 fanout346 (.A(_03501_),
    .X(net346));
 sky130_fd_sc_hd__clkbuf_8 fanout347 (.A(_03483_),
    .X(net347));
 sky130_fd_sc_hd__buf_6 fanout348 (.A(net349),
    .X(net348));
 sky130_fd_sc_hd__buf_8 fanout349 (.A(_03470_),
    .X(net349));
 sky130_fd_sc_hd__buf_4 fanout350 (.A(_03469_),
    .X(net350));
 sky130_fd_sc_hd__buf_6 fanout351 (.A(net352),
    .X(net351));
 sky130_fd_sc_hd__buf_6 fanout352 (.A(_03469_),
    .X(net352));
 sky130_fd_sc_hd__buf_12 fanout353 (.A(_03439_),
    .X(net353));
 sky130_fd_sc_hd__clkbuf_16 fanout354 (.A(_03427_),
    .X(net354));
 sky130_fd_sc_hd__buf_12 fanout355 (.A(net356),
    .X(net355));
 sky130_fd_sc_hd__buf_6 fanout356 (.A(_03419_),
    .X(net356));
 sky130_fd_sc_hd__buf_6 fanout357 (.A(net358),
    .X(net357));
 sky130_fd_sc_hd__buf_8 fanout358 (.A(_03357_),
    .X(net358));
 sky130_fd_sc_hd__buf_6 fanout359 (.A(net360),
    .X(net359));
 sky130_fd_sc_hd__buf_8 fanout360 (.A(_03356_),
    .X(net360));
 sky130_fd_sc_hd__buf_4 fanout361 (.A(_03351_),
    .X(net361));
 sky130_fd_sc_hd__clkbuf_4 fanout362 (.A(_04525_),
    .X(net362));
 sky130_fd_sc_hd__buf_8 fanout363 (.A(_03486_),
    .X(net363));
 sky130_fd_sc_hd__buf_6 fanout364 (.A(_03458_),
    .X(net364));
 sky130_fd_sc_hd__clkbuf_8 fanout365 (.A(_03458_),
    .X(net365));
 sky130_fd_sc_hd__buf_8 fanout366 (.A(_03457_),
    .X(net366));
 sky130_fd_sc_hd__buf_6 fanout367 (.A(net368),
    .X(net367));
 sky130_fd_sc_hd__buf_8 fanout368 (.A(_03436_),
    .X(net368));
 sky130_fd_sc_hd__buf_6 fanout369 (.A(net370),
    .X(net369));
 sky130_fd_sc_hd__buf_6 fanout370 (.A(_03432_),
    .X(net370));
 sky130_fd_sc_hd__buf_4 fanout371 (.A(net372),
    .X(net371));
 sky130_fd_sc_hd__buf_6 fanout372 (.A(net373),
    .X(net372));
 sky130_fd_sc_hd__buf_12 fanout373 (.A(_03432_),
    .X(net373));
 sky130_fd_sc_hd__buf_6 fanout374 (.A(net378),
    .X(net374));
 sky130_fd_sc_hd__buf_6 fanout375 (.A(net378),
    .X(net375));
 sky130_fd_sc_hd__buf_6 fanout376 (.A(net377),
    .X(net376));
 sky130_fd_sc_hd__buf_12 fanout377 (.A(net378),
    .X(net377));
 sky130_fd_sc_hd__buf_12 fanout378 (.A(_03431_),
    .X(net378));
 sky130_fd_sc_hd__buf_6 fanout379 (.A(net381),
    .X(net379));
 sky130_fd_sc_hd__buf_6 fanout380 (.A(net381),
    .X(net380));
 sky130_fd_sc_hd__buf_8 fanout381 (.A(net382),
    .X(net381));
 sky130_fd_sc_hd__buf_6 fanout382 (.A(_03431_),
    .X(net382));
 sky130_fd_sc_hd__buf_6 fanout383 (.A(net384),
    .X(net383));
 sky130_fd_sc_hd__buf_12 fanout384 (.A(_03426_),
    .X(net384));
 sky130_fd_sc_hd__buf_12 fanout385 (.A(net388),
    .X(net385));
 sky130_fd_sc_hd__buf_6 fanout386 (.A(net388),
    .X(net386));
 sky130_fd_sc_hd__buf_4 fanout387 (.A(net388),
    .X(net387));
 sky130_fd_sc_hd__buf_6 fanout388 (.A(_03426_),
    .X(net388));
 sky130_fd_sc_hd__buf_6 fanout389 (.A(net390),
    .X(net389));
 sky130_fd_sc_hd__buf_6 fanout390 (.A(net396),
    .X(net390));
 sky130_fd_sc_hd__buf_6 fanout391 (.A(net392),
    .X(net391));
 sky130_fd_sc_hd__buf_8 fanout392 (.A(net396),
    .X(net392));
 sky130_fd_sc_hd__buf_6 fanout393 (.A(net395),
    .X(net393));
 sky130_fd_sc_hd__buf_6 fanout394 (.A(net395),
    .X(net394));
 sky130_fd_sc_hd__buf_6 fanout395 (.A(net396),
    .X(net395));
 sky130_fd_sc_hd__buf_12 fanout396 (.A(_03425_),
    .X(net396));
 sky130_fd_sc_hd__clkbuf_16 fanout397 (.A(_03424_),
    .X(net397));
 sky130_fd_sc_hd__buf_6 fanout398 (.A(_01973_),
    .X(net398));
 sky130_fd_sc_hd__buf_4 fanout399 (.A(_01973_),
    .X(net399));
 sky130_fd_sc_hd__buf_8 fanout400 (.A(_01962_),
    .X(net400));
 sky130_fd_sc_hd__clkbuf_8 fanout401 (.A(_01962_),
    .X(net401));
 sky130_fd_sc_hd__buf_6 fanout402 (.A(_01951_),
    .X(net402));
 sky130_fd_sc_hd__buf_4 fanout403 (.A(_01951_),
    .X(net403));
 sky130_fd_sc_hd__buf_6 fanout404 (.A(_01940_),
    .X(net404));
 sky130_fd_sc_hd__buf_4 fanout405 (.A(_01940_),
    .X(net405));
 sky130_fd_sc_hd__buf_6 fanout406 (.A(_01929_),
    .X(net406));
 sky130_fd_sc_hd__clkbuf_8 fanout407 (.A(_01929_),
    .X(net407));
 sky130_fd_sc_hd__buf_8 fanout408 (.A(_01918_),
    .X(net408));
 sky130_fd_sc_hd__buf_4 fanout409 (.A(_01918_),
    .X(net409));
 sky130_fd_sc_hd__buf_8 fanout410 (.A(_01907_),
    .X(net410));
 sky130_fd_sc_hd__buf_4 fanout411 (.A(_01907_),
    .X(net411));
 sky130_fd_sc_hd__buf_8 fanout412 (.A(_01896_),
    .X(net412));
 sky130_fd_sc_hd__buf_4 fanout413 (.A(_01896_),
    .X(net413));
 sky130_fd_sc_hd__buf_8 fanout414 (.A(_01885_),
    .X(net414));
 sky130_fd_sc_hd__clkbuf_8 fanout415 (.A(_01885_),
    .X(net415));
 sky130_fd_sc_hd__buf_8 fanout416 (.A(_01874_),
    .X(net416));
 sky130_fd_sc_hd__buf_4 fanout417 (.A(_01874_),
    .X(net417));
 sky130_fd_sc_hd__buf_8 fanout418 (.A(_01863_),
    .X(net418));
 sky130_fd_sc_hd__clkbuf_8 fanout419 (.A(_01863_),
    .X(net419));
 sky130_fd_sc_hd__clkbuf_16 fanout420 (.A(_01852_),
    .X(net420));
 sky130_fd_sc_hd__buf_6 fanout421 (.A(_01852_),
    .X(net421));
 sky130_fd_sc_hd__buf_6 fanout422 (.A(_01841_),
    .X(net422));
 sky130_fd_sc_hd__clkbuf_4 fanout423 (.A(_01841_),
    .X(net423));
 sky130_fd_sc_hd__buf_8 fanout424 (.A(_01830_),
    .X(net424));
 sky130_fd_sc_hd__clkbuf_4 fanout425 (.A(_01830_),
    .X(net425));
 sky130_fd_sc_hd__buf_8 fanout426 (.A(_01820_),
    .X(net426));
 sky130_fd_sc_hd__buf_6 fanout427 (.A(_01820_),
    .X(net427));
 sky130_fd_sc_hd__buf_6 fanout428 (.A(net429),
    .X(net428));
 sky130_fd_sc_hd__buf_6 fanout429 (.A(_01809_),
    .X(net429));
 sky130_fd_sc_hd__buf_6 fanout430 (.A(_01798_),
    .X(net430));
 sky130_fd_sc_hd__buf_4 fanout431 (.A(_01798_),
    .X(net431));
 sky130_fd_sc_hd__buf_8 fanout432 (.A(_01787_),
    .X(net432));
 sky130_fd_sc_hd__buf_4 fanout433 (.A(_01787_),
    .X(net433));
 sky130_fd_sc_hd__buf_8 fanout434 (.A(_01777_),
    .X(net434));
 sky130_fd_sc_hd__buf_4 fanout435 (.A(_01777_),
    .X(net435));
 sky130_fd_sc_hd__clkbuf_16 fanout436 (.A(_01763_),
    .X(net436));
 sky130_fd_sc_hd__buf_4 fanout437 (.A(_01763_),
    .X(net437));
 sky130_fd_sc_hd__buf_8 fanout438 (.A(_01753_),
    .X(net438));
 sky130_fd_sc_hd__clkbuf_4 fanout439 (.A(_01753_),
    .X(net439));
 sky130_fd_sc_hd__buf_8 fanout440 (.A(_01743_),
    .X(net440));
 sky130_fd_sc_hd__buf_4 fanout441 (.A(_01743_),
    .X(net441));
 sky130_fd_sc_hd__buf_8 fanout442 (.A(_01729_),
    .X(net442));
 sky130_fd_sc_hd__buf_4 fanout443 (.A(_01729_),
    .X(net443));
 sky130_fd_sc_hd__buf_8 fanout444 (.A(_01718_),
    .X(net444));
 sky130_fd_sc_hd__buf_4 fanout445 (.A(_01718_),
    .X(net445));
 sky130_fd_sc_hd__buf_6 fanout446 (.A(net447),
    .X(net446));
 sky130_fd_sc_hd__buf_6 fanout447 (.A(_01707_),
    .X(net447));
 sky130_fd_sc_hd__buf_8 fanout448 (.A(_01696_),
    .X(net448));
 sky130_fd_sc_hd__buf_4 fanout449 (.A(_01696_),
    .X(net449));
 sky130_fd_sc_hd__buf_6 fanout450 (.A(_01685_),
    .X(net450));
 sky130_fd_sc_hd__clkbuf_4 fanout451 (.A(_01685_),
    .X(net451));
 sky130_fd_sc_hd__buf_8 fanout452 (.A(_01674_),
    .X(net452));
 sky130_fd_sc_hd__clkbuf_8 fanout453 (.A(_01674_),
    .X(net453));
 sky130_fd_sc_hd__buf_6 fanout454 (.A(_01663_),
    .X(net454));
 sky130_fd_sc_hd__buf_4 fanout455 (.A(_01663_),
    .X(net455));
 sky130_fd_sc_hd__buf_8 fanout456 (.A(_01652_),
    .X(net456));
 sky130_fd_sc_hd__buf_4 fanout457 (.A(_01652_),
    .X(net457));
 sky130_fd_sc_hd__buf_6 fanout458 (.A(_03372_),
    .X(net458));
 sky130_fd_sc_hd__buf_4 fanout459 (.A(net460),
    .X(net459));
 sky130_fd_sc_hd__buf_6 fanout460 (.A(net478),
    .X(net460));
 sky130_fd_sc_hd__buf_8 fanout461 (.A(net462),
    .X(net461));
 sky130_fd_sc_hd__buf_8 fanout462 (.A(net478),
    .X(net462));
 sky130_fd_sc_hd__buf_4 fanout463 (.A(net465),
    .X(net463));
 sky130_fd_sc_hd__buf_4 fanout464 (.A(net465),
    .X(net464));
 sky130_fd_sc_hd__clkbuf_4 fanout465 (.A(net467),
    .X(net465));
 sky130_fd_sc_hd__buf_6 fanout466 (.A(net467),
    .X(net466));
 sky130_fd_sc_hd__clkbuf_4 fanout467 (.A(net468),
    .X(net467));
 sky130_fd_sc_hd__buf_6 fanout468 (.A(net478),
    .X(net468));
 sky130_fd_sc_hd__buf_6 fanout469 (.A(net470),
    .X(net469));
 sky130_fd_sc_hd__buf_6 fanout470 (.A(net478),
    .X(net470));
 sky130_fd_sc_hd__buf_4 fanout471 (.A(net477),
    .X(net471));
 sky130_fd_sc_hd__buf_2 fanout472 (.A(net477),
    .X(net472));
 sky130_fd_sc_hd__buf_4 fanout473 (.A(net474),
    .X(net473));
 sky130_fd_sc_hd__clkbuf_4 fanout474 (.A(net477),
    .X(net474));
 sky130_fd_sc_hd__buf_4 fanout475 (.A(net476),
    .X(net475));
 sky130_fd_sc_hd__clkbuf_8 fanout476 (.A(net477),
    .X(net476));
 sky130_fd_sc_hd__buf_4 fanout477 (.A(net478),
    .X(net477));
 sky130_fd_sc_hd__buf_6 fanout478 (.A(_03355_),
    .X(net478));
 sky130_fd_sc_hd__buf_4 fanout479 (.A(net481),
    .X(net479));
 sky130_fd_sc_hd__clkbuf_4 fanout480 (.A(net481),
    .X(net480));
 sky130_fd_sc_hd__buf_8 fanout481 (.A(net510),
    .X(net481));
 sky130_fd_sc_hd__buf_4 fanout482 (.A(net489),
    .X(net482));
 sky130_fd_sc_hd__buf_4 fanout483 (.A(net484),
    .X(net483));
 sky130_fd_sc_hd__buf_6 fanout484 (.A(net489),
    .X(net484));
 sky130_fd_sc_hd__buf_6 fanout485 (.A(net488),
    .X(net485));
 sky130_fd_sc_hd__buf_4 fanout486 (.A(net487),
    .X(net486));
 sky130_fd_sc_hd__buf_4 fanout487 (.A(net488),
    .X(net487));
 sky130_fd_sc_hd__buf_4 fanout488 (.A(net489),
    .X(net488));
 sky130_fd_sc_hd__clkbuf_8 fanout489 (.A(net510),
    .X(net489));
 sky130_fd_sc_hd__buf_6 fanout490 (.A(net493),
    .X(net490));
 sky130_fd_sc_hd__buf_4 fanout491 (.A(net493),
    .X(net491));
 sky130_fd_sc_hd__clkbuf_4 fanout492 (.A(net493),
    .X(net492));
 sky130_fd_sc_hd__buf_4 fanout493 (.A(net510),
    .X(net493));
 sky130_fd_sc_hd__buf_4 fanout494 (.A(net496),
    .X(net494));
 sky130_fd_sc_hd__buf_2 fanout495 (.A(net496),
    .X(net495));
 sky130_fd_sc_hd__clkbuf_8 fanout496 (.A(net510),
    .X(net496));
 sky130_fd_sc_hd__buf_4 fanout497 (.A(net498),
    .X(net497));
 sky130_fd_sc_hd__buf_4 fanout498 (.A(net510),
    .X(net498));
 sky130_fd_sc_hd__buf_4 fanout499 (.A(net509),
    .X(net499));
 sky130_fd_sc_hd__clkbuf_4 fanout500 (.A(net509),
    .X(net500));
 sky130_fd_sc_hd__buf_4 fanout501 (.A(net502),
    .X(net501));
 sky130_fd_sc_hd__buf_4 fanout502 (.A(net509),
    .X(net502));
 sky130_fd_sc_hd__buf_4 fanout503 (.A(net505),
    .X(net503));
 sky130_fd_sc_hd__buf_4 fanout504 (.A(net505),
    .X(net504));
 sky130_fd_sc_hd__buf_4 fanout505 (.A(net509),
    .X(net505));
 sky130_fd_sc_hd__buf_4 fanout506 (.A(net508),
    .X(net506));
 sky130_fd_sc_hd__clkbuf_4 fanout507 (.A(net508),
    .X(net507));
 sky130_fd_sc_hd__clkbuf_8 fanout508 (.A(net509),
    .X(net508));
 sky130_fd_sc_hd__buf_4 fanout509 (.A(net510),
    .X(net509));
 sky130_fd_sc_hd__buf_8 fanout510 (.A(_03355_),
    .X(net510));
 sky130_fd_sc_hd__clkbuf_16 fanout511 (.A(net512),
    .X(net511));
 sky130_fd_sc_hd__buf_6 fanout512 (.A(net518),
    .X(net512));
 sky130_fd_sc_hd__clkbuf_4 fanout513 (.A(net514),
    .X(net513));
 sky130_fd_sc_hd__buf_4 fanout514 (.A(net517),
    .X(net514));
 sky130_fd_sc_hd__clkbuf_4 fanout515 (.A(net517),
    .X(net515));
 sky130_fd_sc_hd__buf_4 fanout516 (.A(net517),
    .X(net516));
 sky130_fd_sc_hd__buf_6 fanout517 (.A(net518),
    .X(net517));
 sky130_fd_sc_hd__buf_4 fanout518 (.A(net525),
    .X(net518));
 sky130_fd_sc_hd__buf_8 fanout519 (.A(net521),
    .X(net519));
 sky130_fd_sc_hd__clkbuf_2 fanout520 (.A(net521),
    .X(net520));
 sky130_fd_sc_hd__clkbuf_4 fanout521 (.A(net522),
    .X(net521));
 sky130_fd_sc_hd__buf_4 fanout522 (.A(net525),
    .X(net522));
 sky130_fd_sc_hd__buf_4 fanout523 (.A(net525),
    .X(net523));
 sky130_fd_sc_hd__buf_4 fanout524 (.A(net525),
    .X(net524));
 sky130_fd_sc_hd__buf_4 fanout525 (.A(net536),
    .X(net525));
 sky130_fd_sc_hd__clkbuf_4 fanout526 (.A(net527),
    .X(net526));
 sky130_fd_sc_hd__buf_4 fanout527 (.A(net529),
    .X(net527));
 sky130_fd_sc_hd__buf_4 fanout528 (.A(net529),
    .X(net528));
 sky130_fd_sc_hd__clkbuf_4 fanout529 (.A(net530),
    .X(net529));
 sky130_fd_sc_hd__buf_4 fanout530 (.A(net536),
    .X(net530));
 sky130_fd_sc_hd__buf_4 fanout531 (.A(net533),
    .X(net531));
 sky130_fd_sc_hd__buf_4 fanout532 (.A(net533),
    .X(net532));
 sky130_fd_sc_hd__clkbuf_4 fanout533 (.A(net536),
    .X(net533));
 sky130_fd_sc_hd__clkbuf_8 fanout534 (.A(net536),
    .X(net534));
 sky130_fd_sc_hd__buf_8 fanout535 (.A(net536),
    .X(net535));
 sky130_fd_sc_hd__buf_6 fanout536 (.A(_03354_),
    .X(net536));
 sky130_fd_sc_hd__clkbuf_4 fanout537 (.A(net539),
    .X(net537));
 sky130_fd_sc_hd__clkbuf_4 fanout538 (.A(net539),
    .X(net538));
 sky130_fd_sc_hd__buf_4 fanout539 (.A(net555),
    .X(net539));
 sky130_fd_sc_hd__buf_4 fanout540 (.A(net543),
    .X(net540));
 sky130_fd_sc_hd__buf_4 fanout541 (.A(net543),
    .X(net541));
 sky130_fd_sc_hd__clkbuf_2 fanout542 (.A(net543),
    .X(net542));
 sky130_fd_sc_hd__clkbuf_4 fanout543 (.A(net555),
    .X(net543));
 sky130_fd_sc_hd__clkbuf_4 fanout544 (.A(net545),
    .X(net544));
 sky130_fd_sc_hd__buf_2 fanout545 (.A(net555),
    .X(net545));
 sky130_fd_sc_hd__clkbuf_4 fanout546 (.A(net547),
    .X(net546));
 sky130_fd_sc_hd__buf_4 fanout547 (.A(net548),
    .X(net547));
 sky130_fd_sc_hd__buf_2 fanout548 (.A(net555),
    .X(net548));
 sky130_fd_sc_hd__buf_4 fanout549 (.A(net554),
    .X(net549));
 sky130_fd_sc_hd__clkbuf_4 fanout550 (.A(net554),
    .X(net550));
 sky130_fd_sc_hd__clkbuf_2 fanout551 (.A(net554),
    .X(net551));
 sky130_fd_sc_hd__clkbuf_4 fanout552 (.A(net553),
    .X(net552));
 sky130_fd_sc_hd__buf_2 fanout553 (.A(net554),
    .X(net553));
 sky130_fd_sc_hd__buf_4 fanout554 (.A(net555),
    .X(net554));
 sky130_fd_sc_hd__buf_6 fanout555 (.A(_03354_),
    .X(net555));
 sky130_fd_sc_hd__clkbuf_4 fanout556 (.A(net566),
    .X(net556));
 sky130_fd_sc_hd__buf_6 fanout557 (.A(net566),
    .X(net557));
 sky130_fd_sc_hd__buf_4 fanout558 (.A(net560),
    .X(net558));
 sky130_fd_sc_hd__clkbuf_8 fanout559 (.A(net560),
    .X(net559));
 sky130_fd_sc_hd__buf_4 fanout560 (.A(net565),
    .X(net560));
 sky130_fd_sc_hd__clkbuf_4 fanout561 (.A(net565),
    .X(net561));
 sky130_fd_sc_hd__buf_2 fanout562 (.A(net565),
    .X(net562));
 sky130_fd_sc_hd__buf_4 fanout563 (.A(net565),
    .X(net563));
 sky130_fd_sc_hd__buf_2 fanout564 (.A(net565),
    .X(net564));
 sky130_fd_sc_hd__clkbuf_4 fanout565 (.A(net566),
    .X(net565));
 sky130_fd_sc_hd__buf_4 fanout566 (.A(_03354_),
    .X(net566));
 sky130_fd_sc_hd__clkbuf_4 fanout567 (.A(net573),
    .X(net567));
 sky130_fd_sc_hd__clkbuf_2 fanout568 (.A(net573),
    .X(net568));
 sky130_fd_sc_hd__clkbuf_4 fanout569 (.A(net573),
    .X(net569));
 sky130_fd_sc_hd__clkbuf_4 fanout570 (.A(net571),
    .X(net570));
 sky130_fd_sc_hd__buf_2 fanout571 (.A(net572),
    .X(net571));
 sky130_fd_sc_hd__clkbuf_4 fanout572 (.A(net573),
    .X(net572));
 sky130_fd_sc_hd__clkbuf_4 fanout573 (.A(net578),
    .X(net573));
 sky130_fd_sc_hd__buf_4 fanout574 (.A(net578),
    .X(net574));
 sky130_fd_sc_hd__buf_4 fanout575 (.A(net578),
    .X(net575));
 sky130_fd_sc_hd__buf_4 fanout576 (.A(net578),
    .X(net576));
 sky130_fd_sc_hd__clkbuf_4 fanout577 (.A(net578),
    .X(net577));
 sky130_fd_sc_hd__buf_4 fanout578 (.A(_03354_),
    .X(net578));
 sky130_fd_sc_hd__clkbuf_8 fanout579 (.A(_02313_),
    .X(net579));
 sky130_fd_sc_hd__buf_2 fanout580 (.A(_02313_),
    .X(net580));
 sky130_fd_sc_hd__buf_6 fanout581 (.A(_02313_),
    .X(net581));
 sky130_fd_sc_hd__clkbuf_16 fanout582 (.A(_02312_),
    .X(net582));
 sky130_fd_sc_hd__buf_2 fanout583 (.A(_02312_),
    .X(net583));
 sky130_fd_sc_hd__buf_8 fanout584 (.A(_02312_),
    .X(net584));
 sky130_fd_sc_hd__buf_4 fanout585 (.A(_02312_),
    .X(net585));
 sky130_fd_sc_hd__clkbuf_8 fanout586 (.A(_02228_),
    .X(net586));
 sky130_fd_sc_hd__buf_4 fanout587 (.A(_02228_),
    .X(net587));
 sky130_fd_sc_hd__buf_6 fanout588 (.A(_02228_),
    .X(net588));
 sky130_fd_sc_hd__clkbuf_8 fanout589 (.A(net590),
    .X(net589));
 sky130_fd_sc_hd__buf_12 fanout590 (.A(_02227_),
    .X(net590));
 sky130_fd_sc_hd__buf_6 fanout591 (.A(net592),
    .X(net591));
 sky130_fd_sc_hd__buf_12 fanout592 (.A(net167),
    .X(net592));
 sky130_fd_sc_hd__buf_6 fanout593 (.A(_04522_),
    .X(net593));
 sky130_fd_sc_hd__clkbuf_16 fanout594 (.A(_03733_),
    .X(net594));
 sky130_fd_sc_hd__buf_4 fanout595 (.A(_03733_),
    .X(net595));
 sky130_fd_sc_hd__clkbuf_16 fanout596 (.A(_03732_),
    .X(net596));
 sky130_fd_sc_hd__clkbuf_4 fanout597 (.A(_03732_),
    .X(net597));
 sky130_fd_sc_hd__buf_6 fanout598 (.A(_03352_),
    .X(net598));
 sky130_fd_sc_hd__buf_6 fanout599 (.A(_02283_),
    .X(net599));
 sky130_fd_sc_hd__buf_8 fanout600 (.A(_02268_),
    .X(net600));
 sky130_fd_sc_hd__buf_4 fanout601 (.A(_02268_),
    .X(net601));
 sky130_fd_sc_hd__clkbuf_8 fanout602 (.A(net603),
    .X(net602));
 sky130_fd_sc_hd__buf_4 fanout603 (.A(net607),
    .X(net603));
 sky130_fd_sc_hd__clkbuf_8 fanout604 (.A(net607),
    .X(net604));
 sky130_fd_sc_hd__buf_8 fanout605 (.A(net607),
    .X(net605));
 sky130_fd_sc_hd__buf_4 fanout606 (.A(net607),
    .X(net606));
 sky130_fd_sc_hd__clkbuf_8 fanout607 (.A(_02231_),
    .X(net607));
 sky130_fd_sc_hd__buf_6 fanout608 (.A(net612),
    .X(net608));
 sky130_fd_sc_hd__clkbuf_4 fanout609 (.A(net612),
    .X(net609));
 sky130_fd_sc_hd__buf_4 fanout610 (.A(net612),
    .X(net610));
 sky130_fd_sc_hd__buf_6 fanout611 (.A(net612),
    .X(net611));
 sky130_fd_sc_hd__buf_4 fanout612 (.A(net615),
    .X(net612));
 sky130_fd_sc_hd__buf_4 fanout613 (.A(net614),
    .X(net613));
 sky130_fd_sc_hd__clkbuf_4 fanout614 (.A(net615),
    .X(net614));
 sky130_fd_sc_hd__clkbuf_4 fanout615 (.A(_02231_),
    .X(net615));
 sky130_fd_sc_hd__buf_6 fanout616 (.A(net621),
    .X(net616));
 sky130_fd_sc_hd__buf_2 fanout617 (.A(net621),
    .X(net617));
 sky130_fd_sc_hd__buf_6 fanout618 (.A(net621),
    .X(net618));
 sky130_fd_sc_hd__buf_6 fanout619 (.A(net621),
    .X(net619));
 sky130_fd_sc_hd__clkbuf_4 fanout620 (.A(net621),
    .X(net620));
 sky130_fd_sc_hd__buf_8 fanout621 (.A(_02231_),
    .X(net621));
 sky130_fd_sc_hd__buf_4 fanout622 (.A(net626),
    .X(net622));
 sky130_fd_sc_hd__buf_4 fanout623 (.A(net626),
    .X(net623));
 sky130_fd_sc_hd__buf_8 fanout624 (.A(net625),
    .X(net624));
 sky130_fd_sc_hd__buf_6 fanout625 (.A(net626),
    .X(net625));
 sky130_fd_sc_hd__buf_4 fanout626 (.A(_02231_),
    .X(net626));
 sky130_fd_sc_hd__clkbuf_16 fanout627 (.A(_02230_),
    .X(net627));
 sky130_fd_sc_hd__buf_12 fanout628 (.A(_02230_),
    .X(net628));
 sky130_fd_sc_hd__clkbuf_8 fanout629 (.A(net630),
    .X(net629));
 sky130_fd_sc_hd__buf_12 fanout630 (.A(_02224_),
    .X(net630));
 sky130_fd_sc_hd__buf_6 fanout631 (.A(net632),
    .X(net631));
 sky130_fd_sc_hd__clkbuf_4 fanout632 (.A(net633),
    .X(net632));
 sky130_fd_sc_hd__clkbuf_2 fanout633 (.A(net637),
    .X(net633));
 sky130_fd_sc_hd__clkbuf_4 fanout634 (.A(net635),
    .X(net634));
 sky130_fd_sc_hd__buf_4 fanout635 (.A(net636),
    .X(net635));
 sky130_fd_sc_hd__buf_4 fanout636 (.A(net637),
    .X(net636));
 sky130_fd_sc_hd__buf_8 fanout637 (.A(_01641_),
    .X(net637));
 sky130_fd_sc_hd__clkbuf_16 fanout638 (.A(_01621_),
    .X(net638));
 sky130_fd_sc_hd__clkbuf_16 fanout639 (.A(_01621_),
    .X(net639));
 sky130_fd_sc_hd__clkbuf_16 fanout640 (.A(_01620_),
    .X(net640));
 sky130_fd_sc_hd__buf_8 fanout641 (.A(_01620_),
    .X(net641));
 sky130_fd_sc_hd__buf_6 fanout642 (.A(net643),
    .X(net642));
 sky130_fd_sc_hd__buf_8 fanout643 (.A(_01619_),
    .X(net643));
 sky130_fd_sc_hd__buf_6 fanout644 (.A(_01618_),
    .X(net644));
 sky130_fd_sc_hd__buf_6 fanout645 (.A(_01618_),
    .X(net645));
 sky130_fd_sc_hd__buf_6 fanout646 (.A(net647),
    .X(net646));
 sky130_fd_sc_hd__buf_8 fanout647 (.A(_01617_),
    .X(net647));
 sky130_fd_sc_hd__buf_4 fanout648 (.A(_01614_),
    .X(net648));
 sky130_fd_sc_hd__buf_2 fanout649 (.A(_01614_),
    .X(net649));
 sky130_fd_sc_hd__buf_4 fanout650 (.A(net651),
    .X(net650));
 sky130_fd_sc_hd__clkbuf_4 fanout651 (.A(net652),
    .X(net651));
 sky130_fd_sc_hd__buf_4 fanout652 (.A(\tms1x00.Y[3] ),
    .X(net652));
 sky130_fd_sc_hd__clkbuf_4 fanout653 (.A(net654),
    .X(net653));
 sky130_fd_sc_hd__clkbuf_4 fanout654 (.A(\tms1x00.Y[2] ),
    .X(net654));
 sky130_fd_sc_hd__clkbuf_4 fanout655 (.A(\tms1x00.Y[1] ),
    .X(net655));
 sky130_fd_sc_hd__buf_4 fanout656 (.A(\tms1x00.Y[0] ),
    .X(net656));
 sky130_fd_sc_hd__buf_6 fanout657 (.A(\tms1x00.O_latch[4] ),
    .X(net657));
 sky130_fd_sc_hd__buf_8 fanout658 (.A(\tms1x00.O_latch[4] ),
    .X(net658));
 sky130_fd_sc_hd__clkbuf_16 fanout659 (.A(\tms1x00.O_latch[3] ),
    .X(net659));
 sky130_fd_sc_hd__buf_12 fanout660 (.A(\tms1x00.O_latch[3] ),
    .X(net660));
 sky130_fd_sc_hd__buf_8 fanout661 (.A(\tms1x00.O_latch[2] ),
    .X(net661));
 sky130_fd_sc_hd__buf_6 fanout662 (.A(\tms1x00.O_latch[2] ),
    .X(net662));
 sky130_fd_sc_hd__buf_6 fanout663 (.A(\tms1x00.O_latch[1] ),
    .X(net663));
 sky130_fd_sc_hd__buf_8 fanout664 (.A(\tms1x00.O_latch[1] ),
    .X(net664));
 sky130_fd_sc_hd__buf_12 fanout665 (.A(net666),
    .X(net665));
 sky130_fd_sc_hd__buf_12 fanout666 (.A(\tms1x00.O_latch[0] ),
    .X(net666));
 sky130_fd_sc_hd__buf_8 fanout667 (.A(net669),
    .X(net667));
 sky130_fd_sc_hd__buf_8 fanout668 (.A(net669),
    .X(net668));
 sky130_fd_sc_hd__buf_12 fanout669 (.A(\tms1x00.ins_arg[0] ),
    .X(net669));
 sky130_fd_sc_hd__buf_8 fanout670 (.A(net671),
    .X(net670));
 sky130_fd_sc_hd__clkbuf_16 fanout671 (.A(\tms1x00.ins_arg[0] ),
    .X(net671));
 sky130_fd_sc_hd__clkbuf_16 fanout672 (.A(net676),
    .X(net672));
 sky130_fd_sc_hd__buf_8 fanout673 (.A(net676),
    .X(net673));
 sky130_fd_sc_hd__buf_6 fanout674 (.A(net675),
    .X(net674));
 sky130_fd_sc_hd__buf_6 fanout675 (.A(net676),
    .X(net675));
 sky130_fd_sc_hd__clkbuf_16 fanout676 (.A(\tms1x00.ins_arg[1] ),
    .X(net676));
 sky130_fd_sc_hd__buf_6 fanout677 (.A(net678),
    .X(net677));
 sky130_fd_sc_hd__buf_4 fanout678 (.A(net679),
    .X(net678));
 sky130_fd_sc_hd__buf_12 fanout679 (.A(net680),
    .X(net679));
 sky130_fd_sc_hd__buf_12 fanout680 (.A(\tms1x00.ins_arg[2] ),
    .X(net680));
 sky130_fd_sc_hd__buf_8 fanout681 (.A(net682),
    .X(net681));
 sky130_fd_sc_hd__buf_6 fanout682 (.A(net683),
    .X(net682));
 sky130_fd_sc_hd__buf_8 fanout683 (.A(\tms1x00.ins_arg[3] ),
    .X(net683));
 sky130_fd_sc_hd__buf_8 fanout684 (.A(net685),
    .X(net684));
 sky130_fd_sc_hd__buf_6 fanout685 (.A(\tms1x00.ins_arg[3] ),
    .X(net685));
 sky130_fd_sc_hd__buf_8 fanout686 (.A(net690),
    .X(net686));
 sky130_fd_sc_hd__buf_8 fanout687 (.A(net690),
    .X(net687));
 sky130_fd_sc_hd__buf_6 fanout688 (.A(net689),
    .X(net688));
 sky130_fd_sc_hd__buf_6 fanout689 (.A(net690),
    .X(net689));
 sky130_fd_sc_hd__buf_12 fanout690 (.A(\tms1x00.ins_arg[4] ),
    .X(net690));
 sky130_fd_sc_hd__clkbuf_16 fanout691 (.A(net692),
    .X(net691));
 sky130_fd_sc_hd__buf_12 fanout692 (.A(\tms1x00.ins_arg[5] ),
    .X(net692));
 sky130_fd_sc_hd__buf_8 fanout693 (.A(net694),
    .X(net693));
 sky130_fd_sc_hd__clkbuf_8 fanout694 (.A(net695),
    .X(net694));
 sky130_fd_sc_hd__clkbuf_4 fanout695 (.A(\tms1x00.ins_arg[5] ),
    .X(net695));
 sky130_fd_sc_hd__clkbuf_16 fanout696 (.A(net697),
    .X(net696));
 sky130_fd_sc_hd__buf_12 fanout697 (.A(\tms1x00.B[0] ),
    .X(net697));
 sky130_fd_sc_hd__buf_8 fanout698 (.A(net699),
    .X(net698));
 sky130_fd_sc_hd__buf_6 fanout699 (.A(\tms1x00.B[0] ),
    .X(net699));
 sky130_fd_sc_hd__clkbuf_16 fanout700 (.A(net701),
    .X(net700));
 sky130_fd_sc_hd__buf_12 fanout701 (.A(\tms1x00.B[1] ),
    .X(net701));
 sky130_fd_sc_hd__buf_8 fanout702 (.A(net703),
    .X(net702));
 sky130_fd_sc_hd__buf_6 fanout703 (.A(net704),
    .X(net703));
 sky130_fd_sc_hd__buf_4 fanout704 (.A(\tms1x00.B[1] ),
    .X(net704));
 sky130_fd_sc_hd__buf_12 fanout705 (.A(net144),
    .X(net705));
 sky130_fd_sc_hd__clkbuf_8 fanout706 (.A(net707),
    .X(net706));
 sky130_fd_sc_hd__buf_4 fanout707 (.A(_03569_),
    .X(net707));
 sky130_fd_sc_hd__buf_6 fanout708 (.A(_03568_),
    .X(net708));
 sky130_fd_sc_hd__clkbuf_4 fanout709 (.A(_03568_),
    .X(net709));
 sky130_fd_sc_hd__buf_6 fanout710 (.A(_03472_),
    .X(net710));
 sky130_fd_sc_hd__buf_8 fanout711 (.A(_02281_),
    .X(net711));
 sky130_fd_sc_hd__buf_4 fanout712 (.A(net713),
    .X(net712));
 sky130_fd_sc_hd__buf_6 fanout713 (.A(_02280_),
    .X(net713));
 sky130_fd_sc_hd__clkbuf_8 fanout714 (.A(net716),
    .X(net714));
 sky130_fd_sc_hd__buf_6 fanout715 (.A(net716),
    .X(net715));
 sky130_fd_sc_hd__buf_4 fanout716 (.A(net726),
    .X(net716));
 sky130_fd_sc_hd__clkbuf_16 fanout717 (.A(net719),
    .X(net717));
 sky130_fd_sc_hd__buf_4 fanout718 (.A(net719),
    .X(net718));
 sky130_fd_sc_hd__buf_4 fanout719 (.A(net726),
    .X(net719));
 sky130_fd_sc_hd__buf_4 fanout720 (.A(net721),
    .X(net720));
 sky130_fd_sc_hd__clkbuf_4 fanout721 (.A(net726),
    .X(net721));
 sky130_fd_sc_hd__clkbuf_8 fanout722 (.A(net723),
    .X(net722));
 sky130_fd_sc_hd__buf_4 fanout723 (.A(net726),
    .X(net723));
 sky130_fd_sc_hd__clkbuf_8 fanout724 (.A(net725),
    .X(net724));
 sky130_fd_sc_hd__buf_4 fanout725 (.A(net726),
    .X(net725));
 sky130_fd_sc_hd__buf_8 fanout726 (.A(net738),
    .X(net726));
 sky130_fd_sc_hd__buf_6 fanout727 (.A(net728),
    .X(net727));
 sky130_fd_sc_hd__buf_4 fanout728 (.A(net738),
    .X(net728));
 sky130_fd_sc_hd__buf_8 fanout729 (.A(net731),
    .X(net729));
 sky130_fd_sc_hd__buf_6 fanout730 (.A(net731),
    .X(net730));
 sky130_fd_sc_hd__buf_6 fanout731 (.A(net738),
    .X(net731));
 sky130_fd_sc_hd__buf_6 fanout732 (.A(net734),
    .X(net732));
 sky130_fd_sc_hd__buf_6 fanout733 (.A(net734),
    .X(net733));
 sky130_fd_sc_hd__buf_6 fanout734 (.A(net738),
    .X(net734));
 sky130_fd_sc_hd__clkbuf_8 fanout735 (.A(net737),
    .X(net735));
 sky130_fd_sc_hd__clkbuf_4 fanout736 (.A(net737),
    .X(net736));
 sky130_fd_sc_hd__clkbuf_16 fanout737 (.A(net738),
    .X(net737));
 sky130_fd_sc_hd__buf_12 fanout738 (.A(_02245_),
    .X(net738));
 sky130_fd_sc_hd__buf_12 fanout739 (.A(net741),
    .X(net739));
 sky130_fd_sc_hd__buf_8 fanout740 (.A(net741),
    .X(net740));
 sky130_fd_sc_hd__buf_12 fanout741 (.A(_02244_),
    .X(net741));
 sky130_fd_sc_hd__buf_4 fanout742 (.A(net743),
    .X(net742));
 sky130_fd_sc_hd__clkbuf_4 fanout743 (.A(net744),
    .X(net743));
 sky130_fd_sc_hd__buf_6 fanout744 (.A(net755),
    .X(net744));
 sky130_fd_sc_hd__buf_8 fanout745 (.A(net755),
    .X(net745));
 sky130_fd_sc_hd__buf_4 fanout746 (.A(net755),
    .X(net746));
 sky130_fd_sc_hd__clkbuf_8 fanout747 (.A(net749),
    .X(net747));
 sky130_fd_sc_hd__buf_6 fanout748 (.A(net749),
    .X(net748));
 sky130_fd_sc_hd__buf_4 fanout749 (.A(net755),
    .X(net749));
 sky130_fd_sc_hd__buf_4 fanout750 (.A(net751),
    .X(net750));
 sky130_fd_sc_hd__buf_6 fanout751 (.A(net754),
    .X(net751));
 sky130_fd_sc_hd__buf_4 fanout752 (.A(net753),
    .X(net752));
 sky130_fd_sc_hd__buf_6 fanout753 (.A(net754),
    .X(net753));
 sky130_fd_sc_hd__buf_4 fanout754 (.A(net755),
    .X(net754));
 sky130_fd_sc_hd__buf_8 fanout755 (.A(_02243_),
    .X(net755));
 sky130_fd_sc_hd__buf_6 fanout756 (.A(net757),
    .X(net756));
 sky130_fd_sc_hd__buf_6 fanout757 (.A(net761),
    .X(net757));
 sky130_fd_sc_hd__buf_6 fanout758 (.A(net761),
    .X(net758));
 sky130_fd_sc_hd__buf_6 fanout759 (.A(net761),
    .X(net759));
 sky130_fd_sc_hd__buf_2 fanout760 (.A(net761),
    .X(net760));
 sky130_fd_sc_hd__buf_6 fanout761 (.A(_02243_),
    .X(net761));
 sky130_fd_sc_hd__buf_6 fanout762 (.A(net763),
    .X(net762));
 sky130_fd_sc_hd__buf_4 fanout763 (.A(net764),
    .X(net763));
 sky130_fd_sc_hd__buf_4 fanout764 (.A(net765),
    .X(net764));
 sky130_fd_sc_hd__buf_6 fanout765 (.A(_02243_),
    .X(net765));
 sky130_fd_sc_hd__buf_12 fanout766 (.A(net768),
    .X(net766));
 sky130_fd_sc_hd__clkbuf_16 fanout767 (.A(net768),
    .X(net767));
 sky130_fd_sc_hd__buf_12 fanout768 (.A(_02242_),
    .X(net768));
 sky130_fd_sc_hd__buf_6 fanout769 (.A(net771),
    .X(net769));
 sky130_fd_sc_hd__clkbuf_8 fanout770 (.A(net771),
    .X(net770));
 sky130_fd_sc_hd__buf_6 fanout771 (.A(net782),
    .X(net771));
 sky130_fd_sc_hd__buf_6 fanout772 (.A(net782),
    .X(net772));
 sky130_fd_sc_hd__buf_4 fanout773 (.A(net782),
    .X(net773));
 sky130_fd_sc_hd__buf_6 fanout774 (.A(net778),
    .X(net774));
 sky130_fd_sc_hd__buf_4 fanout775 (.A(net776),
    .X(net775));
 sky130_fd_sc_hd__clkbuf_4 fanout776 (.A(net777),
    .X(net776));
 sky130_fd_sc_hd__buf_4 fanout777 (.A(net778),
    .X(net777));
 sky130_fd_sc_hd__buf_4 fanout778 (.A(net782),
    .X(net778));
 sky130_fd_sc_hd__buf_4 fanout779 (.A(net780),
    .X(net779));
 sky130_fd_sc_hd__buf_4 fanout780 (.A(net781),
    .X(net780));
 sky130_fd_sc_hd__clkbuf_4 fanout781 (.A(net782),
    .X(net781));
 sky130_fd_sc_hd__buf_6 fanout782 (.A(net793),
    .X(net782));
 sky130_fd_sc_hd__buf_6 fanout783 (.A(net784),
    .X(net783));
 sky130_fd_sc_hd__buf_6 fanout784 (.A(net793),
    .X(net784));
 sky130_fd_sc_hd__buf_6 fanout785 (.A(net787),
    .X(net785));
 sky130_fd_sc_hd__buf_6 fanout786 (.A(net787),
    .X(net786));
 sky130_fd_sc_hd__buf_6 fanout787 (.A(net793),
    .X(net787));
 sky130_fd_sc_hd__buf_4 fanout788 (.A(net789),
    .X(net788));
 sky130_fd_sc_hd__buf_4 fanout789 (.A(net793),
    .X(net789));
 sky130_fd_sc_hd__buf_8 fanout790 (.A(net792),
    .X(net790));
 sky130_fd_sc_hd__clkbuf_4 fanout791 (.A(net792),
    .X(net791));
 sky130_fd_sc_hd__clkbuf_8 fanout792 (.A(net793),
    .X(net792));
 sky130_fd_sc_hd__buf_12 fanout793 (.A(_02241_),
    .X(net793));
 sky130_fd_sc_hd__buf_12 fanout794 (.A(_02240_),
    .X(net794));
 sky130_fd_sc_hd__clkbuf_16 fanout795 (.A(_02240_),
    .X(net795));
 sky130_fd_sc_hd__buf_6 fanout796 (.A(net797),
    .X(net796));
 sky130_fd_sc_hd__buf_6 fanout797 (.A(net800),
    .X(net797));
 sky130_fd_sc_hd__buf_6 fanout798 (.A(net799),
    .X(net798));
 sky130_fd_sc_hd__buf_6 fanout799 (.A(net800),
    .X(net799));
 sky130_fd_sc_hd__buf_6 fanout800 (.A(net819),
    .X(net800));
 sky130_fd_sc_hd__buf_4 fanout801 (.A(net802),
    .X(net801));
 sky130_fd_sc_hd__buf_4 fanout802 (.A(net804),
    .X(net802));
 sky130_fd_sc_hd__buf_6 fanout803 (.A(net804),
    .X(net803));
 sky130_fd_sc_hd__buf_4 fanout804 (.A(net805),
    .X(net804));
 sky130_fd_sc_hd__buf_6 fanout805 (.A(net819),
    .X(net805));
 sky130_fd_sc_hd__buf_6 fanout806 (.A(net808),
    .X(net806));
 sky130_fd_sc_hd__buf_6 fanout807 (.A(net808),
    .X(net807));
 sky130_fd_sc_hd__buf_4 fanout808 (.A(net819),
    .X(net808));
 sky130_fd_sc_hd__buf_6 fanout809 (.A(net811),
    .X(net809));
 sky130_fd_sc_hd__buf_8 fanout810 (.A(net811),
    .X(net810));
 sky130_fd_sc_hd__buf_6 fanout811 (.A(net819),
    .X(net811));
 sky130_fd_sc_hd__buf_4 fanout812 (.A(net815),
    .X(net812));
 sky130_fd_sc_hd__buf_4 fanout813 (.A(net814),
    .X(net813));
 sky130_fd_sc_hd__clkbuf_8 fanout814 (.A(net815),
    .X(net814));
 sky130_fd_sc_hd__clkbuf_4 fanout815 (.A(net819),
    .X(net815));
 sky130_fd_sc_hd__buf_8 fanout816 (.A(net818),
    .X(net816));
 sky130_fd_sc_hd__buf_4 fanout817 (.A(net818),
    .X(net817));
 sky130_fd_sc_hd__buf_6 fanout818 (.A(net819),
    .X(net818));
 sky130_fd_sc_hd__buf_12 fanout819 (.A(_02239_),
    .X(net819));
 sky130_fd_sc_hd__buf_12 fanout820 (.A(net822),
    .X(net820));
 sky130_fd_sc_hd__buf_12 fanout821 (.A(net822),
    .X(net821));
 sky130_fd_sc_hd__buf_12 fanout822 (.A(_02238_),
    .X(net822));
 sky130_fd_sc_hd__buf_6 fanout823 (.A(net824),
    .X(net823));
 sky130_fd_sc_hd__clkbuf_4 fanout824 (.A(net826),
    .X(net824));
 sky130_fd_sc_hd__buf_6 fanout825 (.A(net826),
    .X(net825));
 sky130_fd_sc_hd__buf_4 fanout826 (.A(net828),
    .X(net826));
 sky130_fd_sc_hd__buf_8 fanout827 (.A(net828),
    .X(net827));
 sky130_fd_sc_hd__buf_6 fanout828 (.A(net846),
    .X(net828));
 sky130_fd_sc_hd__buf_4 fanout829 (.A(net831),
    .X(net829));
 sky130_fd_sc_hd__buf_6 fanout830 (.A(net831),
    .X(net830));
 sky130_fd_sc_hd__buf_4 fanout831 (.A(net846),
    .X(net831));
 sky130_fd_sc_hd__buf_4 fanout832 (.A(net833),
    .X(net832));
 sky130_fd_sc_hd__buf_4 fanout833 (.A(net836),
    .X(net833));
 sky130_fd_sc_hd__clkbuf_8 fanout834 (.A(net836),
    .X(net834));
 sky130_fd_sc_hd__buf_4 fanout835 (.A(net836),
    .X(net835));
 sky130_fd_sc_hd__buf_4 fanout836 (.A(net846),
    .X(net836));
 sky130_fd_sc_hd__buf_6 fanout837 (.A(net838),
    .X(net837));
 sky130_fd_sc_hd__buf_6 fanout838 (.A(net846),
    .X(net838));
 sky130_fd_sc_hd__buf_6 fanout839 (.A(net841),
    .X(net839));
 sky130_fd_sc_hd__buf_6 fanout840 (.A(net841),
    .X(net840));
 sky130_fd_sc_hd__buf_6 fanout841 (.A(net846),
    .X(net841));
 sky130_fd_sc_hd__buf_4 fanout842 (.A(net843),
    .X(net842));
 sky130_fd_sc_hd__buf_6 fanout843 (.A(net844),
    .X(net843));
 sky130_fd_sc_hd__buf_6 fanout844 (.A(net845),
    .X(net844));
 sky130_fd_sc_hd__buf_6 fanout845 (.A(net846),
    .X(net845));
 sky130_fd_sc_hd__buf_12 fanout846 (.A(_02237_),
    .X(net846));
 sky130_fd_sc_hd__buf_12 fanout847 (.A(net849),
    .X(net847));
 sky130_fd_sc_hd__clkbuf_16 fanout848 (.A(net849),
    .X(net848));
 sky130_fd_sc_hd__buf_12 fanout849 (.A(_02236_),
    .X(net849));
 sky130_fd_sc_hd__buf_6 fanout850 (.A(net861),
    .X(net850));
 sky130_fd_sc_hd__clkbuf_8 fanout851 (.A(net861),
    .X(net851));
 sky130_fd_sc_hd__buf_8 fanout852 (.A(net861),
    .X(net852));
 sky130_fd_sc_hd__buf_4 fanout853 (.A(net861),
    .X(net853));
 sky130_fd_sc_hd__buf_4 fanout854 (.A(net857),
    .X(net854));
 sky130_fd_sc_hd__buf_6 fanout855 (.A(net856),
    .X(net855));
 sky130_fd_sc_hd__buf_4 fanout856 (.A(net857),
    .X(net856));
 sky130_fd_sc_hd__clkbuf_4 fanout857 (.A(net860),
    .X(net857));
 sky130_fd_sc_hd__buf_6 fanout858 (.A(net859),
    .X(net858));
 sky130_fd_sc_hd__buf_6 fanout859 (.A(net860),
    .X(net859));
 sky130_fd_sc_hd__buf_4 fanout860 (.A(net861),
    .X(net860));
 sky130_fd_sc_hd__buf_8 fanout861 (.A(_02235_),
    .X(net861));
 sky130_fd_sc_hd__buf_6 fanout862 (.A(net863),
    .X(net862));
 sky130_fd_sc_hd__buf_6 fanout863 (.A(net867),
    .X(net863));
 sky130_fd_sc_hd__clkbuf_16 fanout864 (.A(net867),
    .X(net864));
 sky130_fd_sc_hd__buf_2 fanout865 (.A(net867),
    .X(net865));
 sky130_fd_sc_hd__buf_6 fanout866 (.A(net867),
    .X(net866));
 sky130_fd_sc_hd__buf_8 fanout867 (.A(net873),
    .X(net867));
 sky130_fd_sc_hd__buf_6 fanout868 (.A(net870),
    .X(net868));
 sky130_fd_sc_hd__buf_4 fanout869 (.A(net870),
    .X(net869));
 sky130_fd_sc_hd__buf_6 fanout870 (.A(net873),
    .X(net870));
 sky130_fd_sc_hd__buf_6 fanout871 (.A(net872),
    .X(net871));
 sky130_fd_sc_hd__buf_6 fanout872 (.A(net873),
    .X(net872));
 sky130_fd_sc_hd__buf_8 fanout873 (.A(_02235_),
    .X(net873));
 sky130_fd_sc_hd__buf_12 fanout874 (.A(net876),
    .X(net874));
 sky130_fd_sc_hd__clkbuf_16 fanout875 (.A(net876),
    .X(net875));
 sky130_fd_sc_hd__buf_12 fanout876 (.A(_02234_),
    .X(net876));
 sky130_fd_sc_hd__buf_6 fanout877 (.A(net878),
    .X(net877));
 sky130_fd_sc_hd__buf_6 fanout878 (.A(net887),
    .X(net878));
 sky130_fd_sc_hd__buf_4 fanout879 (.A(net880),
    .X(net879));
 sky130_fd_sc_hd__buf_6 fanout880 (.A(net881),
    .X(net880));
 sky130_fd_sc_hd__clkbuf_4 fanout881 (.A(net887),
    .X(net881));
 sky130_fd_sc_hd__buf_4 fanout882 (.A(net883),
    .X(net882));
 sky130_fd_sc_hd__buf_4 fanout883 (.A(net886),
    .X(net883));
 sky130_fd_sc_hd__buf_6 fanout884 (.A(net886),
    .X(net884));
 sky130_fd_sc_hd__buf_6 fanout885 (.A(net886),
    .X(net885));
 sky130_fd_sc_hd__buf_8 fanout886 (.A(net887),
    .X(net886));
 sky130_fd_sc_hd__buf_8 fanout887 (.A(net901),
    .X(net887));
 sky130_fd_sc_hd__buf_6 fanout888 (.A(net889),
    .X(net888));
 sky130_fd_sc_hd__clkbuf_16 fanout889 (.A(net893),
    .X(net889));
 sky130_fd_sc_hd__clkbuf_4 fanout890 (.A(net893),
    .X(net890));
 sky130_fd_sc_hd__buf_6 fanout891 (.A(net892),
    .X(net891));
 sky130_fd_sc_hd__buf_8 fanout892 (.A(net893),
    .X(net892));
 sky130_fd_sc_hd__buf_8 fanout893 (.A(net901),
    .X(net893));
 sky130_fd_sc_hd__buf_4 fanout894 (.A(net895),
    .X(net894));
 sky130_fd_sc_hd__clkbuf_4 fanout895 (.A(net901),
    .X(net895));
 sky130_fd_sc_hd__clkbuf_8 fanout896 (.A(net897),
    .X(net896));
 sky130_fd_sc_hd__clkbuf_8 fanout897 (.A(net901),
    .X(net897));
 sky130_fd_sc_hd__buf_8 fanout898 (.A(net900),
    .X(net898));
 sky130_fd_sc_hd__buf_4 fanout899 (.A(net900),
    .X(net899));
 sky130_fd_sc_hd__buf_6 fanout900 (.A(net901),
    .X(net900));
 sky130_fd_sc_hd__buf_8 fanout901 (.A(_02233_),
    .X(net901));
 sky130_fd_sc_hd__buf_12 fanout902 (.A(net904),
    .X(net902));
 sky130_fd_sc_hd__clkbuf_16 fanout903 (.A(net904),
    .X(net903));
 sky130_fd_sc_hd__buf_12 fanout904 (.A(_02232_),
    .X(net904));
 sky130_fd_sc_hd__buf_12 fanout905 (.A(_01636_),
    .X(net905));
 sky130_fd_sc_hd__buf_4 fanout906 (.A(_01635_),
    .X(net906));
 sky130_fd_sc_hd__clkbuf_4 fanout907 (.A(_01635_),
    .X(net907));
 sky130_fd_sc_hd__buf_4 fanout908 (.A(net909),
    .X(net908));
 sky130_fd_sc_hd__clkbuf_2 fanout909 (.A(net910),
    .X(net909));
 sky130_fd_sc_hd__buf_6 fanout910 (.A(_01635_),
    .X(net910));
 sky130_fd_sc_hd__buf_6 fanout911 (.A(net913),
    .X(net911));
 sky130_fd_sc_hd__buf_4 fanout912 (.A(net913),
    .X(net912));
 sky130_fd_sc_hd__buf_6 fanout913 (.A(net922),
    .X(net913));
 sky130_fd_sc_hd__buf_4 fanout914 (.A(net916),
    .X(net914));
 sky130_fd_sc_hd__clkbuf_4 fanout915 (.A(net916),
    .X(net915));
 sky130_fd_sc_hd__buf_6 fanout916 (.A(net917),
    .X(net916));
 sky130_fd_sc_hd__buf_8 fanout917 (.A(net922),
    .X(net917));
 sky130_fd_sc_hd__buf_6 fanout918 (.A(net919),
    .X(net918));
 sky130_fd_sc_hd__buf_6 fanout919 (.A(net920),
    .X(net919));
 sky130_fd_sc_hd__buf_6 fanout920 (.A(net922),
    .X(net920));
 sky130_fd_sc_hd__clkbuf_8 fanout921 (.A(net922),
    .X(net921));
 sky130_fd_sc_hd__buf_8 fanout922 (.A(_01634_),
    .X(net922));
 sky130_fd_sc_hd__buf_8 fanout923 (.A(net926),
    .X(net923));
 sky130_fd_sc_hd__clkbuf_4 fanout924 (.A(net926),
    .X(net924));
 sky130_fd_sc_hd__buf_12 fanout925 (.A(net926),
    .X(net925));
 sky130_fd_sc_hd__buf_12 fanout926 (.A(_01633_),
    .X(net926));
 sky130_fd_sc_hd__clkbuf_4 fanout927 (.A(net928),
    .X(net927));
 sky130_fd_sc_hd__clkbuf_4 fanout928 (.A(net929),
    .X(net928));
 sky130_fd_sc_hd__buf_6 fanout929 (.A(net930),
    .X(net929));
 sky130_fd_sc_hd__buf_6 fanout930 (.A(net99),
    .X(net930));
 sky130_fd_sc_hd__buf_6 fanout931 (.A(net932),
    .X(net931));
 sky130_fd_sc_hd__buf_4 fanout932 (.A(net933),
    .X(net932));
 sky130_fd_sc_hd__buf_6 fanout933 (.A(net934),
    .X(net933));
 sky130_fd_sc_hd__buf_6 fanout934 (.A(net99),
    .X(net934));
 sky130_fd_sc_hd__buf_6 fanout935 (.A(net937),
    .X(net935));
 sky130_fd_sc_hd__buf_2 fanout936 (.A(net937),
    .X(net936));
 sky130_fd_sc_hd__buf_12 fanout937 (.A(net98),
    .X(net937));
 sky130_fd_sc_hd__buf_6 fanout938 (.A(net939),
    .X(net938));
 sky130_fd_sc_hd__buf_12 fanout939 (.A(net97),
    .X(net939));
 sky130_fd_sc_hd__buf_6 fanout940 (.A(net941),
    .X(net940));
 sky130_fd_sc_hd__clkbuf_16 fanout941 (.A(net96),
    .X(net941));
 sky130_fd_sc_hd__buf_6 fanout942 (.A(net943),
    .X(net942));
 sky130_fd_sc_hd__clkbuf_16 fanout943 (.A(net95),
    .X(net943));
 sky130_fd_sc_hd__buf_6 fanout944 (.A(net945),
    .X(net944));
 sky130_fd_sc_hd__buf_4 fanout945 (.A(net94),
    .X(net945));
 sky130_fd_sc_hd__buf_8 fanout946 (.A(net94),
    .X(net946));
 sky130_fd_sc_hd__buf_2 fanout947 (.A(net94),
    .X(net947));
 sky130_fd_sc_hd__buf_6 fanout948 (.A(net950),
    .X(net948));
 sky130_fd_sc_hd__buf_6 fanout949 (.A(net950),
    .X(net949));
 sky130_fd_sc_hd__buf_8 fanout950 (.A(net94),
    .X(net950));
 sky130_fd_sc_hd__buf_8 fanout951 (.A(net958),
    .X(net951));
 sky130_fd_sc_hd__clkbuf_8 fanout952 (.A(net958),
    .X(net952));
 sky130_fd_sc_hd__buf_8 fanout953 (.A(net958),
    .X(net953));
 sky130_fd_sc_hd__buf_2 fanout954 (.A(net958),
    .X(net954));
 sky130_fd_sc_hd__buf_6 fanout955 (.A(net957),
    .X(net955));
 sky130_fd_sc_hd__clkbuf_2 fanout956 (.A(net957),
    .X(net956));
 sky130_fd_sc_hd__buf_6 fanout957 (.A(net958),
    .X(net957));
 sky130_fd_sc_hd__buf_12 fanout958 (.A(net93),
    .X(net958));
 sky130_fd_sc_hd__buf_8 fanout959 (.A(net960),
    .X(net959));
 sky130_fd_sc_hd__clkbuf_16 fanout960 (.A(net92),
    .X(net960));
 sky130_fd_sc_hd__buf_6 fanout961 (.A(net962),
    .X(net961));
 sky130_fd_sc_hd__buf_6 fanout962 (.A(net92),
    .X(net962));
 sky130_fd_sc_hd__buf_6 fanout963 (.A(net965),
    .X(net963));
 sky130_fd_sc_hd__buf_4 fanout964 (.A(net965),
    .X(net964));
 sky130_fd_sc_hd__buf_12 fanout965 (.A(net967),
    .X(net965));
 sky130_fd_sc_hd__buf_8 fanout966 (.A(net967),
    .X(net966));
 sky130_fd_sc_hd__clkbuf_16 fanout967 (.A(net91),
    .X(net967));
 sky130_fd_sc_hd__buf_12 fanout968 (.A(net90),
    .X(net968));
 sky130_fd_sc_hd__buf_4 fanout969 (.A(net90),
    .X(net969));
 sky130_fd_sc_hd__buf_6 fanout970 (.A(net971),
    .X(net970));
 sky130_fd_sc_hd__clkbuf_16 fanout971 (.A(net90),
    .X(net971));
 sky130_fd_sc_hd__buf_12 fanout972 (.A(net89),
    .X(net972));
 sky130_fd_sc_hd__clkbuf_8 fanout973 (.A(net89),
    .X(net973));
 sky130_fd_sc_hd__buf_6 fanout974 (.A(net975),
    .X(net974));
 sky130_fd_sc_hd__clkbuf_16 fanout975 (.A(net89),
    .X(net975));
 sky130_fd_sc_hd__buf_6 fanout976 (.A(net978),
    .X(net976));
 sky130_fd_sc_hd__buf_6 fanout977 (.A(net978),
    .X(net977));
 sky130_fd_sc_hd__buf_8 fanout978 (.A(net983),
    .X(net978));
 sky130_fd_sc_hd__buf_6 fanout979 (.A(net983),
    .X(net979));
 sky130_fd_sc_hd__buf_6 fanout980 (.A(net981),
    .X(net980));
 sky130_fd_sc_hd__buf_8 fanout981 (.A(net982),
    .X(net981));
 sky130_fd_sc_hd__clkbuf_16 fanout982 (.A(net983),
    .X(net982));
 sky130_fd_sc_hd__clkbuf_16 fanout983 (.A(net88),
    .X(net983));
 sky130_fd_sc_hd__buf_12 fanout984 (.A(net85),
    .X(net984));
 sky130_fd_sc_hd__buf_8 fanout985 (.A(net84),
    .X(net985));
 sky130_fd_sc_hd__buf_4 fanout986 (.A(net987),
    .X(net986));
 sky130_fd_sc_hd__buf_12 fanout987 (.A(net989),
    .X(net987));
 sky130_fd_sc_hd__buf_6 fanout988 (.A(net989),
    .X(net988));
 sky130_fd_sc_hd__buf_12 fanout989 (.A(net83),
    .X(net989));
 sky130_fd_sc_hd__buf_6 fanout990 (.A(net991),
    .X(net990));
 sky130_fd_sc_hd__clkbuf_16 fanout991 (.A(net995),
    .X(net991));
 sky130_fd_sc_hd__clkbuf_8 fanout992 (.A(net994),
    .X(net992));
 sky130_fd_sc_hd__buf_4 fanout993 (.A(net994),
    .X(net993));
 sky130_fd_sc_hd__buf_12 fanout994 (.A(net995),
    .X(net994));
 sky130_fd_sc_hd__clkbuf_16 fanout995 (.A(net1000),
    .X(net995));
 sky130_fd_sc_hd__buf_6 fanout996 (.A(net997),
    .X(net996));
 sky130_fd_sc_hd__buf_6 fanout997 (.A(net999),
    .X(net997));
 sky130_fd_sc_hd__buf_8 fanout998 (.A(net999),
    .X(net998));
 sky130_fd_sc_hd__buf_12 fanout999 (.A(net1000),
    .X(net999));
 sky130_fd_sc_hd__buf_2 hold1 (.A(feedback_delay),
    .X(net1133));
 sky130_fd_sc_hd__clkbuf_4 input1 (.A(io_in[5]),
    .X(net1));
 sky130_fd_sc_hd__buf_2 input10 (.A(rom_value[0]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_4 input100 (.A(wbs_dat_i[20]),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_4 input101 (.A(wbs_dat_i[21]),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_2 input102 (.A(wbs_dat_i[22]),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_8 input103 (.A(wbs_dat_i[23]),
    .X(net103));
 sky130_fd_sc_hd__buf_4 input104 (.A(wbs_dat_i[24]),
    .X(net104));
 sky130_fd_sc_hd__buf_6 input105 (.A(wbs_dat_i[25]),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_2 input106 (.A(wbs_dat_i[26]),
    .X(net106));
 sky130_fd_sc_hd__buf_4 input107 (.A(wbs_dat_i[27]),
    .X(net107));
 sky130_fd_sc_hd__buf_4 input108 (.A(wbs_dat_i[28]),
    .X(net108));
 sky130_fd_sc_hd__buf_6 input109 (.A(wbs_dat_i[29]),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(rom_value[10]),
    .X(net11));
 sky130_fd_sc_hd__buf_2 input110 (.A(wbs_dat_i[2]),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_8 input111 (.A(wbs_dat_i[3]),
    .X(net111));
 sky130_fd_sc_hd__buf_6 input112 (.A(wbs_dat_i[4]),
    .X(net112));
 sky130_fd_sc_hd__buf_2 input113 (.A(wbs_dat_i[5]),
    .X(net113));
 sky130_fd_sc_hd__buf_6 input114 (.A(wbs_dat_i[6]),
    .X(net114));
 sky130_fd_sc_hd__buf_6 input115 (.A(wbs_dat_i[7]),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_4 input116 (.A(wbs_dat_i[8]),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_16 input117 (.A(wbs_dat_i[9]),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_2 input118 (.A(wbs_stb_i),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_16 input119 (.A(wbs_we_i),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(rom_value[11]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 input13 (.A(rom_value[12]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(rom_value[13]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 input15 (.A(rom_value[14]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(rom_value[15]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(rom_value[16]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(rom_value[17]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(rom_value[18]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(io_in[6]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(rom_value[19]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(rom_value[1]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(rom_value[20]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(rom_value[21]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(rom_value[22]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(rom_value[23]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(rom_value[24]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(rom_value[25]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_2 input28 (.A(rom_value[26]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_2 input29 (.A(rom_value[27]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(io_in[7]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input30 (.A(rom_value[28]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_2 input31 (.A(rom_value[29]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 input32 (.A(rom_value[2]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(rom_value[30]),
    .X(net33));
 sky130_fd_sc_hd__buf_2 input34 (.A(rom_value[31]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 input35 (.A(rom_value[3]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 input36 (.A(rom_value[4]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_2 input37 (.A(rom_value[5]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_2 input38 (.A(rom_value[6]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_2 input39 (.A(rom_value[7]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(io_in[8]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input40 (.A(rom_value[8]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_2 input41 (.A(rom_value[9]),
    .X(net41));
 sky130_fd_sc_hd__buf_2 input42 (.A(wb_rom_val[0]),
    .X(net42));
 sky130_fd_sc_hd__buf_2 input43 (.A(wb_rom_val[10]),
    .X(net43));
 sky130_fd_sc_hd__buf_2 input44 (.A(wb_rom_val[11]),
    .X(net44));
 sky130_fd_sc_hd__buf_2 input45 (.A(wb_rom_val[12]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_4 input46 (.A(wb_rom_val[13]),
    .X(net46));
 sky130_fd_sc_hd__buf_2 input47 (.A(wb_rom_val[14]),
    .X(net47));
 sky130_fd_sc_hd__buf_2 input48 (.A(wb_rom_val[15]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_4 input49 (.A(wb_rom_val[16]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(io_in[9]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_4 input50 (.A(wb_rom_val[17]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_4 input51 (.A(wb_rom_val[18]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_4 input52 (.A(wb_rom_val[19]),
    .X(net52));
 sky130_fd_sc_hd__buf_2 input53 (.A(wb_rom_val[1]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_4 input54 (.A(wb_rom_val[20]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_4 input55 (.A(wb_rom_val[21]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_4 input56 (.A(wb_rom_val[22]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_4 input57 (.A(wb_rom_val[23]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_4 input58 (.A(wb_rom_val[24]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_4 input59 (.A(wb_rom_val[25]),
    .X(net59));
 sky130_fd_sc_hd__buf_4 input6 (.A(ram_val_in[0]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_4 input60 (.A(wb_rom_val[26]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_4 input61 (.A(wb_rom_val[27]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_4 input62 (.A(wb_rom_val[28]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_4 input63 (.A(wb_rom_val[29]),
    .X(net63));
 sky130_fd_sc_hd__buf_2 input64 (.A(wb_rom_val[2]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_4 input65 (.A(wb_rom_val[30]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_4 input66 (.A(wb_rom_val[31]),
    .X(net66));
 sky130_fd_sc_hd__buf_2 input67 (.A(wb_rom_val[3]),
    .X(net67));
 sky130_fd_sc_hd__buf_2 input68 (.A(wb_rom_val[4]),
    .X(net68));
 sky130_fd_sc_hd__buf_2 input69 (.A(wb_rom_val[5]),
    .X(net69));
 sky130_fd_sc_hd__buf_4 input7 (.A(ram_val_in[1]),
    .X(net7));
 sky130_fd_sc_hd__buf_2 input70 (.A(wb_rom_val[6]),
    .X(net70));
 sky130_fd_sc_hd__buf_2 input71 (.A(wb_rom_val[7]),
    .X(net71));
 sky130_fd_sc_hd__buf_2 input72 (.A(wb_rom_val[8]),
    .X(net72));
 sky130_fd_sc_hd__buf_2 input73 (.A(wb_rom_val[9]),
    .X(net73));
 sky130_fd_sc_hd__buf_12 input74 (.A(wb_rst_i),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_4 input75 (.A(wbs_adr_i[10]),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_4 input76 (.A(wbs_adr_i[16]),
    .X(net76));
 sky130_fd_sc_hd__buf_6 input77 (.A(wbs_adr_i[17]),
    .X(net77));
 sky130_fd_sc_hd__buf_8 input78 (.A(wbs_adr_i[23]),
    .X(net78));
 sky130_fd_sc_hd__buf_2 input79 (.A(wbs_adr_i[2]),
    .X(net79));
 sky130_fd_sc_hd__buf_4 input8 (.A(ram_val_in[2]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input80 (.A(wbs_adr_i[3]),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_2 input81 (.A(wbs_adr_i[4]),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_2 input82 (.A(wbs_adr_i[5]),
    .X(net82));
 sky130_fd_sc_hd__buf_2 input83 (.A(wbs_adr_i[6]),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_4 input84 (.A(wbs_adr_i[7]),
    .X(net84));
 sky130_fd_sc_hd__buf_4 input85 (.A(wbs_adr_i[8]),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_4 input86 (.A(wbs_adr_i[9]),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_2 input87 (.A(wbs_cyc_i),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_2 input88 (.A(wbs_dat_i[0]),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_16 input89 (.A(wbs_dat_i[10]),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_8 input9 (.A(ram_val_in[3]),
    .X(net9));
 sky130_fd_sc_hd__buf_8 input90 (.A(wbs_dat_i[11]),
    .X(net90));
 sky130_fd_sc_hd__buf_2 input91 (.A(wbs_dat_i[12]),
    .X(net91));
 sky130_fd_sc_hd__buf_8 input92 (.A(wbs_dat_i[13]),
    .X(net92));
 sky130_fd_sc_hd__buf_2 input93 (.A(wbs_dat_i[14]),
    .X(net93));
 sky130_fd_sc_hd__buf_8 input94 (.A(wbs_dat_i[15]),
    .X(net94));
 sky130_fd_sc_hd__buf_4 input95 (.A(wbs_dat_i[16]),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_2 input96 (.A(wbs_dat_i[17]),
    .X(net96));
 sky130_fd_sc_hd__buf_6 input97 (.A(wbs_dat_i[18]),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_4 input98 (.A(wbs_dat_i[19]),
    .X(net98));
 sky130_fd_sc_hd__buf_4 input99 (.A(wbs_dat_i[1]),
    .X(net99));
 sky130_fd_sc_hd__buf_4 output120 (.A(net120),
    .X(io_out[10]));
 sky130_fd_sc_hd__buf_4 output121 (.A(net121),
    .X(io_out[11]));
 sky130_fd_sc_hd__buf_4 output122 (.A(net122),
    .X(io_out[12]));
 sky130_fd_sc_hd__buf_4 output123 (.A(net123),
    .X(io_out[13]));
 sky130_fd_sc_hd__buf_4 output124 (.A(net124),
    .X(io_out[14]));
 sky130_fd_sc_hd__buf_4 output125 (.A(net125),
    .X(io_out[15]));
 sky130_fd_sc_hd__buf_4 output126 (.A(net126),
    .X(io_out[16]));
 sky130_fd_sc_hd__buf_4 output127 (.A(net127),
    .X(io_out[17]));
 sky130_fd_sc_hd__buf_4 output128 (.A(net128),
    .X(io_out[18]));
 sky130_fd_sc_hd__buf_4 output129 (.A(net129),
    .X(io_out[19]));
 sky130_fd_sc_hd__buf_4 output130 (.A(net130),
    .X(io_out[20]));
 sky130_fd_sc_hd__buf_4 output131 (.A(net131),
    .X(io_out[21]));
 sky130_fd_sc_hd__buf_4 output132 (.A(net132),
    .X(io_out[22]));
 sky130_fd_sc_hd__buf_4 output133 (.A(net133),
    .X(io_out[23]));
 sky130_fd_sc_hd__buf_4 output134 (.A(net134),
    .X(io_out[24]));
 sky130_fd_sc_hd__buf_4 output135 (.A(net135),
    .X(io_out[25]));
 sky130_fd_sc_hd__buf_4 output136 (.A(net136),
    .X(io_out[26]));
 sky130_fd_sc_hd__buf_4 output137 (.A(net137),
    .X(io_out[27]));
 sky130_fd_sc_hd__buf_4 output138 (.A(net138),
    .X(io_out[28]));
 sky130_fd_sc_hd__buf_4 output139 (.A(net139),
    .X(io_out[29]));
 sky130_fd_sc_hd__buf_4 output140 (.A(net140),
    .X(io_out[30]));
 sky130_fd_sc_hd__buf_4 output141 (.A(net141),
    .X(io_out[31]));
 sky130_fd_sc_hd__buf_4 output142 (.A(net142),
    .X(io_out[32]));
 sky130_fd_sc_hd__buf_4 output143 (.A(net143),
    .X(io_out[33]));
 sky130_fd_sc_hd__buf_4 output144 (.A(net144),
    .X(io_out[36]));
 sky130_fd_sc_hd__buf_4 output145 (.A(net145),
    .X(io_out[37]));
 sky130_fd_sc_hd__buf_4 output146 (.A(net146),
    .X(ram_addr[0]));
 sky130_fd_sc_hd__buf_4 output147 (.A(net147),
    .X(ram_addr[1]));
 sky130_fd_sc_hd__buf_4 output148 (.A(net148),
    .X(ram_addr[2]));
 sky130_fd_sc_hd__buf_4 output149 (.A(net149),
    .X(ram_addr[3]));
 sky130_fd_sc_hd__buf_4 output150 (.A(net150),
    .X(ram_addr[4]));
 sky130_fd_sc_hd__buf_4 output151 (.A(net151),
    .X(ram_addr[5]));
 sky130_fd_sc_hd__buf_4 output152 (.A(net152),
    .X(ram_addr[6]));
 sky130_fd_sc_hd__buf_4 output153 (.A(net153),
    .X(ram_val_out[0]));
 sky130_fd_sc_hd__buf_4 output154 (.A(net154),
    .X(ram_val_out[1]));
 sky130_fd_sc_hd__buf_4 output155 (.A(net155),
    .X(ram_val_out[2]));
 sky130_fd_sc_hd__buf_4 output156 (.A(net156),
    .X(ram_val_out[3]));
 sky130_fd_sc_hd__buf_4 output157 (.A(net157),
    .X(ram_we));
 sky130_fd_sc_hd__buf_4 output158 (.A(net158),
    .X(rom_addr[0]));
 sky130_fd_sc_hd__buf_4 output159 (.A(net159),
    .X(rom_addr[1]));
 sky130_fd_sc_hd__buf_4 output160 (.A(net160),
    .X(rom_addr[2]));
 sky130_fd_sc_hd__buf_4 output161 (.A(net161),
    .X(rom_addr[3]));
 sky130_fd_sc_hd__buf_4 output162 (.A(net162),
    .X(rom_addr[4]));
 sky130_fd_sc_hd__buf_4 output163 (.A(net163),
    .X(rom_addr[5]));
 sky130_fd_sc_hd__buf_4 output164 (.A(net164),
    .X(rom_addr[6]));
 sky130_fd_sc_hd__buf_4 output165 (.A(net165),
    .X(rom_addr[7]));
 sky130_fd_sc_hd__buf_4 output166 (.A(net166),
    .X(rom_addr[8]));
 sky130_fd_sc_hd__buf_4 output167 (.A(net592),
    .X(rom_csb));
 sky130_fd_sc_hd__buf_4 output168 (.A(net168),
    .X(wb_rom_adrb[0]));
 sky130_fd_sc_hd__buf_4 output169 (.A(net169),
    .X(wb_rom_adrb[1]));
 sky130_fd_sc_hd__buf_4 output170 (.A(net170),
    .X(wb_rom_adrb[2]));
 sky130_fd_sc_hd__buf_4 output171 (.A(net171),
    .X(wb_rom_adrb[3]));
 sky130_fd_sc_hd__buf_4 output172 (.A(net172),
    .X(wb_rom_adrb[4]));
 sky130_fd_sc_hd__buf_4 output173 (.A(net173),
    .X(wb_rom_adrb[5]));
 sky130_fd_sc_hd__buf_4 output174 (.A(net174),
    .X(wb_rom_adrb[6]));
 sky130_fd_sc_hd__buf_4 output175 (.A(net175),
    .X(wb_rom_adrb[7]));
 sky130_fd_sc_hd__buf_4 output176 (.A(net176),
    .X(wb_rom_adrb[8]));
 sky130_fd_sc_hd__buf_4 output177 (.A(net177),
    .X(wb_rom_csb));
 sky130_fd_sc_hd__buf_4 output178 (.A(net178),
    .X(wb_rom_web));
 sky130_fd_sc_hd__buf_4 output179 (.A(net179),
    .X(wbs_ack_o));
 sky130_fd_sc_hd__buf_4 output180 (.A(net180),
    .X(wbs_dat_o[0]));
 sky130_fd_sc_hd__buf_4 output181 (.A(net181),
    .X(wbs_dat_o[10]));
 sky130_fd_sc_hd__buf_4 output182 (.A(net182),
    .X(wbs_dat_o[11]));
 sky130_fd_sc_hd__buf_4 output183 (.A(net183),
    .X(wbs_dat_o[12]));
 sky130_fd_sc_hd__buf_4 output184 (.A(net184),
    .X(wbs_dat_o[13]));
 sky130_fd_sc_hd__buf_4 output185 (.A(net185),
    .X(wbs_dat_o[14]));
 sky130_fd_sc_hd__buf_4 output186 (.A(net186),
    .X(wbs_dat_o[15]));
 sky130_fd_sc_hd__buf_4 output187 (.A(net187),
    .X(wbs_dat_o[16]));
 sky130_fd_sc_hd__buf_4 output188 (.A(net188),
    .X(wbs_dat_o[17]));
 sky130_fd_sc_hd__buf_4 output189 (.A(net189),
    .X(wbs_dat_o[18]));
 sky130_fd_sc_hd__buf_4 output190 (.A(net190),
    .X(wbs_dat_o[19]));
 sky130_fd_sc_hd__buf_4 output191 (.A(net191),
    .X(wbs_dat_o[1]));
 sky130_fd_sc_hd__buf_4 output192 (.A(net192),
    .X(wbs_dat_o[20]));
 sky130_fd_sc_hd__buf_4 output193 (.A(net193),
    .X(wbs_dat_o[21]));
 sky130_fd_sc_hd__buf_4 output194 (.A(net194),
    .X(wbs_dat_o[22]));
 sky130_fd_sc_hd__buf_4 output195 (.A(net195),
    .X(wbs_dat_o[23]));
 sky130_fd_sc_hd__buf_4 output196 (.A(net196),
    .X(wbs_dat_o[24]));
 sky130_fd_sc_hd__buf_4 output197 (.A(net197),
    .X(wbs_dat_o[25]));
 sky130_fd_sc_hd__buf_4 output198 (.A(net198),
    .X(wbs_dat_o[26]));
 sky130_fd_sc_hd__buf_4 output199 (.A(net199),
    .X(wbs_dat_o[27]));
 sky130_fd_sc_hd__buf_4 output200 (.A(net200),
    .X(wbs_dat_o[28]));
 sky130_fd_sc_hd__buf_4 output201 (.A(net201),
    .X(wbs_dat_o[29]));
 sky130_fd_sc_hd__buf_4 output202 (.A(net202),
    .X(wbs_dat_o[2]));
 sky130_fd_sc_hd__buf_4 output203 (.A(net203),
    .X(wbs_dat_o[30]));
 sky130_fd_sc_hd__buf_4 output204 (.A(net204),
    .X(wbs_dat_o[31]));
 sky130_fd_sc_hd__buf_4 output205 (.A(net205),
    .X(wbs_dat_o[3]));
 sky130_fd_sc_hd__buf_4 output206 (.A(net206),
    .X(wbs_dat_o[4]));
 sky130_fd_sc_hd__buf_4 output207 (.A(net207),
    .X(wbs_dat_o[5]));
 sky130_fd_sc_hd__buf_4 output208 (.A(net208),
    .X(wbs_dat_o[6]));
 sky130_fd_sc_hd__buf_4 output209 (.A(net209),
    .X(wbs_dat_o[7]));
 sky130_fd_sc_hd__buf_4 output210 (.A(net210),
    .X(wbs_dat_o[8]));
 sky130_fd_sc_hd__buf_4 output211 (.A(net211),
    .X(wbs_dat_o[9]));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1080 (.LO(net1080));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1081 (.LO(net1081));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1082 (.LO(net1082));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1083 (.LO(net1083));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1084 (.LO(net1084));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1085 (.LO(net1085));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1086 (.LO(net1086));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1087 (.LO(net1087));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1088 (.LO(net1088));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1089 (.LO(net1089));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1090 (.LO(net1090));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1091 (.LO(net1091));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1092 (.LO(net1092));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1093 (.LO(net1093));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1094 (.LO(net1094));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1095 (.LO(net1095));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1096 (.LO(net1096));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1097 (.LO(net1097));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1098 (.LO(net1098));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1099 (.LO(net1099));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1100 (.LO(net1100));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1101 (.LO(net1101));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1102 (.LO(net1102));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1103 (.LO(net1103));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1104 (.LO(net1104));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1105 (.LO(net1105));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1106 (.LO(net1106));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1107 (.LO(net1107));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1108 (.LO(net1108));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1109 (.LO(net1109));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1110 (.LO(net1110));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1111 (.LO(net1111));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1112 (.LO(net1112));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1113 (.LO(net1113));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1114 (.LO(net1114));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1115 (.LO(net1115));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1116 (.LO(net1116));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1117 (.LO(net1117));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1118 (.LO(net1118));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1119 (.LO(net1119));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1120 (.LO(net1120));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1121 (.LO(net1121));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1122 (.LO(net1122));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1123 (.HI(net1123));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1124 (.HI(net1124));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1125 (.HI(net1125));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1126 (.HI(net1126));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1127 (.HI(net1127));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1128 (.HI(net1128));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1129 (.HI(net1129));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1130 (.HI(net1130));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1131 (.HI(net1131));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_1132 (.HI(net1132));
 assign io_oeb[0] = net1123;
 assign io_oeb[10] = net1080;
 assign io_oeb[11] = net1081;
 assign io_oeb[12] = net1082;
 assign io_oeb[13] = net1083;
 assign io_oeb[14] = net1084;
 assign io_oeb[15] = net1085;
 assign io_oeb[16] = net1086;
 assign io_oeb[17] = net1087;
 assign io_oeb[18] = net1088;
 assign io_oeb[19] = net1089;
 assign io_oeb[1] = net1124;
 assign io_oeb[20] = net1090;
 assign io_oeb[21] = net1091;
 assign io_oeb[22] = net1092;
 assign io_oeb[23] = net1093;
 assign io_oeb[24] = net1094;
 assign io_oeb[25] = net1095;
 assign io_oeb[26] = net1096;
 assign io_oeb[27] = net1097;
 assign io_oeb[28] = net1098;
 assign io_oeb[29] = net1099;
 assign io_oeb[2] = net1125;
 assign io_oeb[30] = net1100;
 assign io_oeb[31] = net1101;
 assign io_oeb[32] = net1102;
 assign io_oeb[33] = net1103;
 assign io_oeb[34] = net1104;
 assign io_oeb[35] = net1105;
 assign io_oeb[36] = net1106;
 assign io_oeb[37] = net1107;
 assign io_oeb[3] = net1126;
 assign io_oeb[4] = net1127;
 assign io_oeb[5] = net1128;
 assign io_oeb[6] = net1129;
 assign io_oeb[7] = net1130;
 assign io_oeb[8] = net1131;
 assign io_oeb[9] = net1132;
 assign io_out[0] = net1108;
 assign io_out[1] = net1109;
 assign io_out[2] = net1110;
 assign io_out[34] = net1118;
 assign io_out[35] = net1119;
 assign io_out[3] = net1111;
 assign io_out[4] = net1112;
 assign io_out[5] = net1113;
 assign io_out[6] = net1114;
 assign io_out[7] = net1115;
 assign io_out[8] = net1116;
 assign io_out[9] = net1117;
 assign irq[0] = net1120;
 assign irq[1] = net1121;
 assign irq[2] = net1122;
endmodule

