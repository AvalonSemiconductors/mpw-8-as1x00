VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_tms1x00
  CLASS BLOCK ;
  FOREIGN wrapped_tms1x00 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1000.000 BY 1000.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 996.000 6.350 1000.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.270 996.000 268.550 1000.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.490 996.000 294.770 1000.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.710 996.000 320.990 1000.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.930 996.000 347.210 1000.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.150 996.000 373.430 1000.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 996.000 399.650 1000.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.590 996.000 425.870 1000.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.810 996.000 452.090 1000.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.030 996.000 478.310 1000.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.250 996.000 504.530 1000.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 996.000 32.570 1000.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.470 996.000 530.750 1000.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.690 996.000 556.970 1000.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.910 996.000 583.190 1000.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.130 996.000 609.410 1000.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 635.350 996.000 635.630 1000.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.570 996.000 661.850 1000.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 687.790 996.000 688.070 1000.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.010 996.000 714.290 1000.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.230 996.000 740.510 1000.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.450 996.000 766.730 1000.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 996.000 58.790 1000.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.670 996.000 792.950 1000.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.890 996.000 819.170 1000.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 845.110 996.000 845.390 1000.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.330 996.000 871.610 1000.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 897.550 996.000 897.830 1000.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 923.770 996.000 924.050 1000.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.990 996.000 950.270 1000.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 976.210 996.000 976.490 1000.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 996.000 85.010 1000.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.950 996.000 111.230 1000.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.170 996.000 137.450 1000.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 996.000 163.670 1000.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.610 996.000 189.890 1000.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 996.000 216.110 1000.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.050 996.000 242.330 1000.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 996.000 15.090 1000.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 996.000 277.290 1000.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.230 996.000 303.510 1000.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.450 996.000 329.730 1000.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.670 996.000 355.950 1000.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.890 996.000 382.170 1000.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.110 996.000 408.390 1000.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.330 996.000 434.610 1000.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 996.000 460.830 1000.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.770 996.000 487.050 1000.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.990 996.000 513.270 1000.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 996.000 41.310 1000.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.210 996.000 539.490 1000.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.430 996.000 565.710 1000.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.650 996.000 591.930 1000.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.870 996.000 618.150 1000.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.090 996.000 644.370 1000.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.310 996.000 670.590 1000.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.530 996.000 696.810 1000.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.750 996.000 723.030 1000.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.970 996.000 749.250 1000.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.190 996.000 775.470 1000.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 996.000 67.530 1000.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.410 996.000 801.690 1000.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 827.630 996.000 827.910 1000.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.850 996.000 854.130 1000.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 880.070 996.000 880.350 1000.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 906.290 996.000 906.570 1000.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.510 996.000 932.790 1000.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 958.730 996.000 959.010 1000.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 984.950 996.000 985.230 1000.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 996.000 93.750 1000.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 996.000 119.970 1000.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.910 996.000 146.190 1000.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.130 996.000 172.410 1000.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.350 996.000 198.630 1000.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.570 996.000 224.850 1000.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.790 996.000 251.070 1000.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 996.000 23.830 1000.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.750 996.000 286.030 1000.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.970 996.000 312.250 1000.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 996.000 338.470 1000.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.410 996.000 364.690 1000.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.630 996.000 390.910 1000.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.850 996.000 417.130 1000.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.070 996.000 443.350 1000.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.290 996.000 469.570 1000.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.510 996.000 495.790 1000.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.730 996.000 522.010 1000.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 996.000 50.050 1000.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.950 996.000 548.230 1000.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.170 996.000 574.450 1000.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 600.390 996.000 600.670 1000.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.610 996.000 626.890 1000.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.830 996.000 653.110 1000.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.050 996.000 679.330 1000.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.270 996.000 705.550 1000.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.490 996.000 731.770 1000.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 757.710 996.000 757.990 1000.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.930 996.000 784.210 1000.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 996.000 76.270 1000.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 810.150 996.000 810.430 1000.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 836.370 996.000 836.650 1000.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 862.590 996.000 862.870 1000.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.810 996.000 889.090 1000.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.030 996.000 915.310 1000.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 941.250 996.000 941.530 1000.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 967.470 996.000 967.750 1000.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 993.690 996.000 993.970 1000.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 996.000 102.490 1000.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.430 996.000 128.710 1000.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 996.000 154.930 1000.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.870 996.000 181.150 1000.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.090 996.000 207.370 1000.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.310 996.000 233.590 1000.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.530 996.000 259.810 1000.000 ;
    END
  END io_out[9]
  PIN oram_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END oram_addr[0]
  PIN oram_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END oram_addr[1]
  PIN oram_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 4.000 131.200 ;
    END
  END oram_addr[2]
  PIN oram_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 4.000 178.800 ;
    END
  END oram_addr[3]
  PIN oram_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.800 4.000 226.400 ;
    END
  END oram_addr[4]
  PIN oram_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 273.400 4.000 274.000 ;
    END
  END oram_addr[5]
  PIN oram_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.000 4.000 321.600 ;
    END
  END oram_addr[6]
  PIN oram_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 368.600 4.000 369.200 ;
    END
  END oram_addr[7]
  PIN oram_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 416.200 4.000 416.800 ;
    END
  END oram_addr[8]
  PIN oram_csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 11.600 4.000 12.200 ;
    END
  END oram_csb
  PIN oram_value[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 4.000 59.800 ;
    END
  END oram_value[0]
  PIN oram_value[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 487.600 4.000 488.200 ;
    END
  END oram_value[10]
  PIN oram_value[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 511.400 4.000 512.000 ;
    END
  END oram_value[11]
  PIN oram_value[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 535.200 4.000 535.800 ;
    END
  END oram_value[12]
  PIN oram_value[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 559.000 4.000 559.600 ;
    END
  END oram_value[13]
  PIN oram_value[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 582.800 4.000 583.400 ;
    END
  END oram_value[14]
  PIN oram_value[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 606.600 4.000 607.200 ;
    END
  END oram_value[15]
  PIN oram_value[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 630.400 4.000 631.000 ;
    END
  END oram_value[16]
  PIN oram_value[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 654.200 4.000 654.800 ;
    END
  END oram_value[17]
  PIN oram_value[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 678.000 4.000 678.600 ;
    END
  END oram_value[18]
  PIN oram_value[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 701.800 4.000 702.400 ;
    END
  END oram_value[19]
  PIN oram_value[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.800 4.000 107.400 ;
    END
  END oram_value[1]
  PIN oram_value[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 725.600 4.000 726.200 ;
    END
  END oram_value[20]
  PIN oram_value[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 749.400 4.000 750.000 ;
    END
  END oram_value[21]
  PIN oram_value[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 773.200 4.000 773.800 ;
    END
  END oram_value[22]
  PIN oram_value[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 797.000 4.000 797.600 ;
    END
  END oram_value[23]
  PIN oram_value[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 820.800 4.000 821.400 ;
    END
  END oram_value[24]
  PIN oram_value[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 844.600 4.000 845.200 ;
    END
  END oram_value[25]
  PIN oram_value[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 868.400 4.000 869.000 ;
    END
  END oram_value[26]
  PIN oram_value[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 892.200 4.000 892.800 ;
    END
  END oram_value[27]
  PIN oram_value[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 916.000 4.000 916.600 ;
    END
  END oram_value[28]
  PIN oram_value[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 939.800 4.000 940.400 ;
    END
  END oram_value[29]
  PIN oram_value[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 154.400 4.000 155.000 ;
    END
  END oram_value[2]
  PIN oram_value[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 963.600 4.000 964.200 ;
    END
  END oram_value[30]
  PIN oram_value[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 987.400 4.000 988.000 ;
    END
  END oram_value[31]
  PIN oram_value[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.000 4.000 202.600 ;
    END
  END oram_value[3]
  PIN oram_value[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 249.600 4.000 250.200 ;
    END
  END oram_value[4]
  PIN oram_value[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.200 4.000 297.800 ;
    END
  END oram_value[5]
  PIN oram_value[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.800 4.000 345.400 ;
    END
  END oram_value[6]
  PIN oram_value[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 392.400 4.000 393.000 ;
    END
  END oram_value[7]
  PIN oram_value[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 440.000 4.000 440.600 ;
    END
  END oram_value[8]
  PIN oram_value[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.800 4.000 464.400 ;
    END
  END oram_value[9]
  PIN ram_adrb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 59.880 1000.000 60.480 ;
    END
  END ram_adrb[0]
  PIN ram_adrb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 106.120 1000.000 106.720 ;
    END
  END ram_adrb[1]
  PIN ram_adrb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 152.360 1000.000 152.960 ;
    END
  END ram_adrb[2]
  PIN ram_adrb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 198.600 1000.000 199.200 ;
    END
  END ram_adrb[3]
  PIN ram_adrb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 244.840 1000.000 245.440 ;
    END
  END ram_adrb[4]
  PIN ram_adrb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 291.080 1000.000 291.680 ;
    END
  END ram_adrb[5]
  PIN ram_adrb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 337.320 1000.000 337.920 ;
    END
  END ram_adrb[6]
  PIN ram_adrb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 383.560 1000.000 384.160 ;
    END
  END ram_adrb[7]
  PIN ram_adrb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 429.800 1000.000 430.400 ;
    END
  END ram_adrb[8]
  PIN ram_csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 13.640 1000.000 14.240 ;
    END
  END ram_csb
  PIN ram_val[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 83.000 1000.000 83.600 ;
    END
  END ram_val[0]
  PIN ram_val[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 499.160 1000.000 499.760 ;
    END
  END ram_val[10]
  PIN ram_val[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 522.280 1000.000 522.880 ;
    END
  END ram_val[11]
  PIN ram_val[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 545.400 1000.000 546.000 ;
    END
  END ram_val[12]
  PIN ram_val[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 568.520 1000.000 569.120 ;
    END
  END ram_val[13]
  PIN ram_val[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 591.640 1000.000 592.240 ;
    END
  END ram_val[14]
  PIN ram_val[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 614.760 1000.000 615.360 ;
    END
  END ram_val[15]
  PIN ram_val[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 637.880 1000.000 638.480 ;
    END
  END ram_val[16]
  PIN ram_val[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 661.000 1000.000 661.600 ;
    END
  END ram_val[17]
  PIN ram_val[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 684.120 1000.000 684.720 ;
    END
  END ram_val[18]
  PIN ram_val[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 707.240 1000.000 707.840 ;
    END
  END ram_val[19]
  PIN ram_val[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 129.240 1000.000 129.840 ;
    END
  END ram_val[1]
  PIN ram_val[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 730.360 1000.000 730.960 ;
    END
  END ram_val[20]
  PIN ram_val[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 753.480 1000.000 754.080 ;
    END
  END ram_val[21]
  PIN ram_val[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 776.600 1000.000 777.200 ;
    END
  END ram_val[22]
  PIN ram_val[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 799.720 1000.000 800.320 ;
    END
  END ram_val[23]
  PIN ram_val[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 822.840 1000.000 823.440 ;
    END
  END ram_val[24]
  PIN ram_val[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 845.960 1000.000 846.560 ;
    END
  END ram_val[25]
  PIN ram_val[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 869.080 1000.000 869.680 ;
    END
  END ram_val[26]
  PIN ram_val[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 892.200 1000.000 892.800 ;
    END
  END ram_val[27]
  PIN ram_val[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 915.320 1000.000 915.920 ;
    END
  END ram_val[28]
  PIN ram_val[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 938.440 1000.000 939.040 ;
    END
  END ram_val[29]
  PIN ram_val[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 175.480 1000.000 176.080 ;
    END
  END ram_val[2]
  PIN ram_val[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 961.560 1000.000 962.160 ;
    END
  END ram_val[30]
  PIN ram_val[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 984.680 1000.000 985.280 ;
    END
  END ram_val[31]
  PIN ram_val[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 221.720 1000.000 222.320 ;
    END
  END ram_val[3]
  PIN ram_val[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 267.960 1000.000 268.560 ;
    END
  END ram_val[4]
  PIN ram_val[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 314.200 1000.000 314.800 ;
    END
  END ram_val[5]
  PIN ram_val[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 360.440 1000.000 361.040 ;
    END
  END ram_val[6]
  PIN ram_val[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 406.680 1000.000 407.280 ;
    END
  END ram_val[7]
  PIN ram_val[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 452.920 1000.000 453.520 ;
    END
  END ram_val[8]
  PIN ram_val[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 476.040 1000.000 476.640 ;
    END
  END ram_val[9]
  PIN ram_web
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 36.760 1000.000 37.360 ;
    END
  END ram_web
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 987.600 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 987.600 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 0.000 12.330 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.710 0.000 21.990 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 0.000 31.650 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 0.000 70.290 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.810 0.000 360.090 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.790 0.000 389.070 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.770 0.000 418.050 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.750 0.000 447.030 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.730 0.000 476.010 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.710 0.000 504.990 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.690 0.000 533.970 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.670 0.000 562.950 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.650 0.000 591.930 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.630 0.000 620.910 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.990 0.000 99.270 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.610 0.000 649.890 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 678.590 0.000 678.870 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.570 0.000 707.850 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 736.550 0.000 736.830 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.530 0.000 765.810 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.510 0.000 794.790 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 823.490 0.000 823.770 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.470 0.000 852.750 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 881.450 0.000 881.730 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 910.430 0.000 910.710 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.970 0.000 128.250 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 939.410 0.000 939.690 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 968.390 0.000 968.670 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.950 0.000 157.230 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 0.000 186.210 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.910 0.000 215.190 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.890 0.000 244.170 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.870 0.000 273.150 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.850 0.000 302.130 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.830 0.000 331.110 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 0.000 41.310 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.670 0.000 79.950 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.470 0.000 369.750 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.450 0.000 398.730 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.430 0.000 427.710 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.410 0.000 456.690 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.390 0.000 485.670 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.370 0.000 514.650 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.350 0.000 543.630 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.330 0.000 572.610 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 601.310 0.000 601.590 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.290 0.000 630.570 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 0.000 108.930 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 659.270 0.000 659.550 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.250 0.000 688.530 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.230 0.000 717.510 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.210 0.000 746.490 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.190 0.000 775.470 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 804.170 0.000 804.450 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 833.150 0.000 833.430 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 862.130 0.000 862.410 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 891.110 0.000 891.390 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 920.090 0.000 920.370 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.630 0.000 137.910 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.070 0.000 949.350 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 978.050 0.000 978.330 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.610 0.000 166.890 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.590 0.000 195.870 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.570 0.000 224.850 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.550 0.000 253.830 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.530 0.000 282.810 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.510 0.000 311.790 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.490 0.000 340.770 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 0.000 89.610 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.130 0.000 379.410 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.110 0.000 408.390 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.090 0.000 437.370 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.070 0.000 466.350 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.050 0.000 495.330 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.030 0.000 524.310 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.010 0.000 553.290 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.990 0.000 582.270 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.970 0.000 611.250 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.950 0.000 640.230 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.310 0.000 118.590 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.930 0.000 669.210 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.910 0.000 698.190 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 726.890 0.000 727.170 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 755.870 0.000 756.150 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.850 0.000 785.130 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 813.830 0.000 814.110 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 842.810 0.000 843.090 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.790 0.000 872.070 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 900.770 0.000 901.050 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 929.750 0.000 930.030 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 958.730 0.000 959.010 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 987.710 0.000 987.990 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.270 0.000 176.550 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.250 0.000 205.530 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.230 0.000 234.510 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.210 0.000 263.490 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.190 0.000 292.470 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.170 0.000 321.450 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.150 0.000 350.430 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 0.000 60.630 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 994.060 987.445 ;
      LAYER met1 ;
        RECT 5.520 1.060 995.370 987.600 ;
      LAYER met2 ;
        RECT 6.990 995.720 14.530 996.610 ;
        RECT 15.370 995.720 23.270 996.610 ;
        RECT 24.110 995.720 32.010 996.610 ;
        RECT 32.850 995.720 40.750 996.610 ;
        RECT 41.590 995.720 49.490 996.610 ;
        RECT 50.330 995.720 58.230 996.610 ;
        RECT 59.070 995.720 66.970 996.610 ;
        RECT 67.810 995.720 75.710 996.610 ;
        RECT 76.550 995.720 84.450 996.610 ;
        RECT 85.290 995.720 93.190 996.610 ;
        RECT 94.030 995.720 101.930 996.610 ;
        RECT 102.770 995.720 110.670 996.610 ;
        RECT 111.510 995.720 119.410 996.610 ;
        RECT 120.250 995.720 128.150 996.610 ;
        RECT 128.990 995.720 136.890 996.610 ;
        RECT 137.730 995.720 145.630 996.610 ;
        RECT 146.470 995.720 154.370 996.610 ;
        RECT 155.210 995.720 163.110 996.610 ;
        RECT 163.950 995.720 171.850 996.610 ;
        RECT 172.690 995.720 180.590 996.610 ;
        RECT 181.430 995.720 189.330 996.610 ;
        RECT 190.170 995.720 198.070 996.610 ;
        RECT 198.910 995.720 206.810 996.610 ;
        RECT 207.650 995.720 215.550 996.610 ;
        RECT 216.390 995.720 224.290 996.610 ;
        RECT 225.130 995.720 233.030 996.610 ;
        RECT 233.870 995.720 241.770 996.610 ;
        RECT 242.610 995.720 250.510 996.610 ;
        RECT 251.350 995.720 259.250 996.610 ;
        RECT 260.090 995.720 267.990 996.610 ;
        RECT 268.830 995.720 276.730 996.610 ;
        RECT 277.570 995.720 285.470 996.610 ;
        RECT 286.310 995.720 294.210 996.610 ;
        RECT 295.050 995.720 302.950 996.610 ;
        RECT 303.790 995.720 311.690 996.610 ;
        RECT 312.530 995.720 320.430 996.610 ;
        RECT 321.270 995.720 329.170 996.610 ;
        RECT 330.010 995.720 337.910 996.610 ;
        RECT 338.750 995.720 346.650 996.610 ;
        RECT 347.490 995.720 355.390 996.610 ;
        RECT 356.230 995.720 364.130 996.610 ;
        RECT 364.970 995.720 372.870 996.610 ;
        RECT 373.710 995.720 381.610 996.610 ;
        RECT 382.450 995.720 390.350 996.610 ;
        RECT 391.190 995.720 399.090 996.610 ;
        RECT 399.930 995.720 407.830 996.610 ;
        RECT 408.670 995.720 416.570 996.610 ;
        RECT 417.410 995.720 425.310 996.610 ;
        RECT 426.150 995.720 434.050 996.610 ;
        RECT 434.890 995.720 442.790 996.610 ;
        RECT 443.630 995.720 451.530 996.610 ;
        RECT 452.370 995.720 460.270 996.610 ;
        RECT 461.110 995.720 469.010 996.610 ;
        RECT 469.850 995.720 477.750 996.610 ;
        RECT 478.590 995.720 486.490 996.610 ;
        RECT 487.330 995.720 495.230 996.610 ;
        RECT 496.070 995.720 503.970 996.610 ;
        RECT 504.810 995.720 512.710 996.610 ;
        RECT 513.550 995.720 521.450 996.610 ;
        RECT 522.290 995.720 530.190 996.610 ;
        RECT 531.030 995.720 538.930 996.610 ;
        RECT 539.770 995.720 547.670 996.610 ;
        RECT 548.510 995.720 556.410 996.610 ;
        RECT 557.250 995.720 565.150 996.610 ;
        RECT 565.990 995.720 573.890 996.610 ;
        RECT 574.730 995.720 582.630 996.610 ;
        RECT 583.470 995.720 591.370 996.610 ;
        RECT 592.210 995.720 600.110 996.610 ;
        RECT 600.950 995.720 608.850 996.610 ;
        RECT 609.690 995.720 617.590 996.610 ;
        RECT 618.430 995.720 626.330 996.610 ;
        RECT 627.170 995.720 635.070 996.610 ;
        RECT 635.910 995.720 643.810 996.610 ;
        RECT 644.650 995.720 652.550 996.610 ;
        RECT 653.390 995.720 661.290 996.610 ;
        RECT 662.130 995.720 670.030 996.610 ;
        RECT 670.870 995.720 678.770 996.610 ;
        RECT 679.610 995.720 687.510 996.610 ;
        RECT 688.350 995.720 696.250 996.610 ;
        RECT 697.090 995.720 704.990 996.610 ;
        RECT 705.830 995.720 713.730 996.610 ;
        RECT 714.570 995.720 722.470 996.610 ;
        RECT 723.310 995.720 731.210 996.610 ;
        RECT 732.050 995.720 739.950 996.610 ;
        RECT 740.790 995.720 748.690 996.610 ;
        RECT 749.530 995.720 757.430 996.610 ;
        RECT 758.270 995.720 766.170 996.610 ;
        RECT 767.010 995.720 774.910 996.610 ;
        RECT 775.750 995.720 783.650 996.610 ;
        RECT 784.490 995.720 792.390 996.610 ;
        RECT 793.230 995.720 801.130 996.610 ;
        RECT 801.970 995.720 809.870 996.610 ;
        RECT 810.710 995.720 818.610 996.610 ;
        RECT 819.450 995.720 827.350 996.610 ;
        RECT 828.190 995.720 836.090 996.610 ;
        RECT 836.930 995.720 844.830 996.610 ;
        RECT 845.670 995.720 853.570 996.610 ;
        RECT 854.410 995.720 862.310 996.610 ;
        RECT 863.150 995.720 871.050 996.610 ;
        RECT 871.890 995.720 879.790 996.610 ;
        RECT 880.630 995.720 888.530 996.610 ;
        RECT 889.370 995.720 897.270 996.610 ;
        RECT 898.110 995.720 906.010 996.610 ;
        RECT 906.850 995.720 914.750 996.610 ;
        RECT 915.590 995.720 923.490 996.610 ;
        RECT 924.330 995.720 932.230 996.610 ;
        RECT 933.070 995.720 940.970 996.610 ;
        RECT 941.810 995.720 949.710 996.610 ;
        RECT 950.550 995.720 958.450 996.610 ;
        RECT 959.290 995.720 967.190 996.610 ;
        RECT 968.030 995.720 975.930 996.610 ;
        RECT 976.770 995.720 984.670 996.610 ;
        RECT 985.510 995.720 993.410 996.610 ;
        RECT 994.250 995.720 995.340 996.610 ;
        RECT 6.990 4.280 995.340 995.720 ;
        RECT 6.990 0.155 11.770 4.280 ;
        RECT 12.610 0.155 21.430 4.280 ;
        RECT 22.270 0.155 31.090 4.280 ;
        RECT 31.930 0.155 40.750 4.280 ;
        RECT 41.590 0.155 50.410 4.280 ;
        RECT 51.250 0.155 60.070 4.280 ;
        RECT 60.910 0.155 69.730 4.280 ;
        RECT 70.570 0.155 79.390 4.280 ;
        RECT 80.230 0.155 89.050 4.280 ;
        RECT 89.890 0.155 98.710 4.280 ;
        RECT 99.550 0.155 108.370 4.280 ;
        RECT 109.210 0.155 118.030 4.280 ;
        RECT 118.870 0.155 127.690 4.280 ;
        RECT 128.530 0.155 137.350 4.280 ;
        RECT 138.190 0.155 147.010 4.280 ;
        RECT 147.850 0.155 156.670 4.280 ;
        RECT 157.510 0.155 166.330 4.280 ;
        RECT 167.170 0.155 175.990 4.280 ;
        RECT 176.830 0.155 185.650 4.280 ;
        RECT 186.490 0.155 195.310 4.280 ;
        RECT 196.150 0.155 204.970 4.280 ;
        RECT 205.810 0.155 214.630 4.280 ;
        RECT 215.470 0.155 224.290 4.280 ;
        RECT 225.130 0.155 233.950 4.280 ;
        RECT 234.790 0.155 243.610 4.280 ;
        RECT 244.450 0.155 253.270 4.280 ;
        RECT 254.110 0.155 262.930 4.280 ;
        RECT 263.770 0.155 272.590 4.280 ;
        RECT 273.430 0.155 282.250 4.280 ;
        RECT 283.090 0.155 291.910 4.280 ;
        RECT 292.750 0.155 301.570 4.280 ;
        RECT 302.410 0.155 311.230 4.280 ;
        RECT 312.070 0.155 320.890 4.280 ;
        RECT 321.730 0.155 330.550 4.280 ;
        RECT 331.390 0.155 340.210 4.280 ;
        RECT 341.050 0.155 349.870 4.280 ;
        RECT 350.710 0.155 359.530 4.280 ;
        RECT 360.370 0.155 369.190 4.280 ;
        RECT 370.030 0.155 378.850 4.280 ;
        RECT 379.690 0.155 388.510 4.280 ;
        RECT 389.350 0.155 398.170 4.280 ;
        RECT 399.010 0.155 407.830 4.280 ;
        RECT 408.670 0.155 417.490 4.280 ;
        RECT 418.330 0.155 427.150 4.280 ;
        RECT 427.990 0.155 436.810 4.280 ;
        RECT 437.650 0.155 446.470 4.280 ;
        RECT 447.310 0.155 456.130 4.280 ;
        RECT 456.970 0.155 465.790 4.280 ;
        RECT 466.630 0.155 475.450 4.280 ;
        RECT 476.290 0.155 485.110 4.280 ;
        RECT 485.950 0.155 494.770 4.280 ;
        RECT 495.610 0.155 504.430 4.280 ;
        RECT 505.270 0.155 514.090 4.280 ;
        RECT 514.930 0.155 523.750 4.280 ;
        RECT 524.590 0.155 533.410 4.280 ;
        RECT 534.250 0.155 543.070 4.280 ;
        RECT 543.910 0.155 552.730 4.280 ;
        RECT 553.570 0.155 562.390 4.280 ;
        RECT 563.230 0.155 572.050 4.280 ;
        RECT 572.890 0.155 581.710 4.280 ;
        RECT 582.550 0.155 591.370 4.280 ;
        RECT 592.210 0.155 601.030 4.280 ;
        RECT 601.870 0.155 610.690 4.280 ;
        RECT 611.530 0.155 620.350 4.280 ;
        RECT 621.190 0.155 630.010 4.280 ;
        RECT 630.850 0.155 639.670 4.280 ;
        RECT 640.510 0.155 649.330 4.280 ;
        RECT 650.170 0.155 658.990 4.280 ;
        RECT 659.830 0.155 668.650 4.280 ;
        RECT 669.490 0.155 678.310 4.280 ;
        RECT 679.150 0.155 687.970 4.280 ;
        RECT 688.810 0.155 697.630 4.280 ;
        RECT 698.470 0.155 707.290 4.280 ;
        RECT 708.130 0.155 716.950 4.280 ;
        RECT 717.790 0.155 726.610 4.280 ;
        RECT 727.450 0.155 736.270 4.280 ;
        RECT 737.110 0.155 745.930 4.280 ;
        RECT 746.770 0.155 755.590 4.280 ;
        RECT 756.430 0.155 765.250 4.280 ;
        RECT 766.090 0.155 774.910 4.280 ;
        RECT 775.750 0.155 784.570 4.280 ;
        RECT 785.410 0.155 794.230 4.280 ;
        RECT 795.070 0.155 803.890 4.280 ;
        RECT 804.730 0.155 813.550 4.280 ;
        RECT 814.390 0.155 823.210 4.280 ;
        RECT 824.050 0.155 832.870 4.280 ;
        RECT 833.710 0.155 842.530 4.280 ;
        RECT 843.370 0.155 852.190 4.280 ;
        RECT 853.030 0.155 861.850 4.280 ;
        RECT 862.690 0.155 871.510 4.280 ;
        RECT 872.350 0.155 881.170 4.280 ;
        RECT 882.010 0.155 890.830 4.280 ;
        RECT 891.670 0.155 900.490 4.280 ;
        RECT 901.330 0.155 910.150 4.280 ;
        RECT 910.990 0.155 919.810 4.280 ;
        RECT 920.650 0.155 929.470 4.280 ;
        RECT 930.310 0.155 939.130 4.280 ;
        RECT 939.970 0.155 948.790 4.280 ;
        RECT 949.630 0.155 958.450 4.280 ;
        RECT 959.290 0.155 968.110 4.280 ;
        RECT 968.950 0.155 977.770 4.280 ;
        RECT 978.610 0.155 987.430 4.280 ;
        RECT 988.270 0.155 995.340 4.280 ;
      LAYER met3 ;
        RECT 4.400 987.000 996.000 987.865 ;
        RECT 4.000 985.680 996.000 987.000 ;
        RECT 4.000 984.280 995.600 985.680 ;
        RECT 4.000 964.600 996.000 984.280 ;
        RECT 4.400 963.200 996.000 964.600 ;
        RECT 4.000 962.560 996.000 963.200 ;
        RECT 4.000 961.160 995.600 962.560 ;
        RECT 4.000 940.800 996.000 961.160 ;
        RECT 4.400 939.440 996.000 940.800 ;
        RECT 4.400 939.400 995.600 939.440 ;
        RECT 4.000 938.040 995.600 939.400 ;
        RECT 4.000 917.000 996.000 938.040 ;
        RECT 4.400 916.320 996.000 917.000 ;
        RECT 4.400 915.600 995.600 916.320 ;
        RECT 4.000 914.920 995.600 915.600 ;
        RECT 4.000 893.200 996.000 914.920 ;
        RECT 4.400 891.800 995.600 893.200 ;
        RECT 4.000 870.080 996.000 891.800 ;
        RECT 4.000 869.400 995.600 870.080 ;
        RECT 4.400 868.680 995.600 869.400 ;
        RECT 4.400 868.000 996.000 868.680 ;
        RECT 4.000 846.960 996.000 868.000 ;
        RECT 4.000 845.600 995.600 846.960 ;
        RECT 4.400 845.560 995.600 845.600 ;
        RECT 4.400 844.200 996.000 845.560 ;
        RECT 4.000 823.840 996.000 844.200 ;
        RECT 4.000 822.440 995.600 823.840 ;
        RECT 4.000 821.800 996.000 822.440 ;
        RECT 4.400 820.400 996.000 821.800 ;
        RECT 4.000 800.720 996.000 820.400 ;
        RECT 4.000 799.320 995.600 800.720 ;
        RECT 4.000 798.000 996.000 799.320 ;
        RECT 4.400 796.600 996.000 798.000 ;
        RECT 4.000 777.600 996.000 796.600 ;
        RECT 4.000 776.200 995.600 777.600 ;
        RECT 4.000 774.200 996.000 776.200 ;
        RECT 4.400 772.800 996.000 774.200 ;
        RECT 4.000 754.480 996.000 772.800 ;
        RECT 4.000 753.080 995.600 754.480 ;
        RECT 4.000 750.400 996.000 753.080 ;
        RECT 4.400 749.000 996.000 750.400 ;
        RECT 4.000 731.360 996.000 749.000 ;
        RECT 4.000 729.960 995.600 731.360 ;
        RECT 4.000 726.600 996.000 729.960 ;
        RECT 4.400 725.200 996.000 726.600 ;
        RECT 4.000 708.240 996.000 725.200 ;
        RECT 4.000 706.840 995.600 708.240 ;
        RECT 4.000 702.800 996.000 706.840 ;
        RECT 4.400 701.400 996.000 702.800 ;
        RECT 4.000 685.120 996.000 701.400 ;
        RECT 4.000 683.720 995.600 685.120 ;
        RECT 4.000 679.000 996.000 683.720 ;
        RECT 4.400 677.600 996.000 679.000 ;
        RECT 4.000 662.000 996.000 677.600 ;
        RECT 4.000 660.600 995.600 662.000 ;
        RECT 4.000 655.200 996.000 660.600 ;
        RECT 4.400 653.800 996.000 655.200 ;
        RECT 4.000 638.880 996.000 653.800 ;
        RECT 4.000 637.480 995.600 638.880 ;
        RECT 4.000 631.400 996.000 637.480 ;
        RECT 4.400 630.000 996.000 631.400 ;
        RECT 4.000 615.760 996.000 630.000 ;
        RECT 4.000 614.360 995.600 615.760 ;
        RECT 4.000 607.600 996.000 614.360 ;
        RECT 4.400 606.200 996.000 607.600 ;
        RECT 4.000 592.640 996.000 606.200 ;
        RECT 4.000 591.240 995.600 592.640 ;
        RECT 4.000 583.800 996.000 591.240 ;
        RECT 4.400 582.400 996.000 583.800 ;
        RECT 4.000 569.520 996.000 582.400 ;
        RECT 4.000 568.120 995.600 569.520 ;
        RECT 4.000 560.000 996.000 568.120 ;
        RECT 4.400 558.600 996.000 560.000 ;
        RECT 4.000 546.400 996.000 558.600 ;
        RECT 4.000 545.000 995.600 546.400 ;
        RECT 4.000 536.200 996.000 545.000 ;
        RECT 4.400 534.800 996.000 536.200 ;
        RECT 4.000 523.280 996.000 534.800 ;
        RECT 4.000 521.880 995.600 523.280 ;
        RECT 4.000 512.400 996.000 521.880 ;
        RECT 4.400 511.000 996.000 512.400 ;
        RECT 4.000 500.160 996.000 511.000 ;
        RECT 4.000 498.760 995.600 500.160 ;
        RECT 4.000 488.600 996.000 498.760 ;
        RECT 4.400 487.200 996.000 488.600 ;
        RECT 4.000 477.040 996.000 487.200 ;
        RECT 4.000 475.640 995.600 477.040 ;
        RECT 4.000 464.800 996.000 475.640 ;
        RECT 4.400 463.400 996.000 464.800 ;
        RECT 4.000 453.920 996.000 463.400 ;
        RECT 4.000 452.520 995.600 453.920 ;
        RECT 4.000 441.000 996.000 452.520 ;
        RECT 4.400 439.600 996.000 441.000 ;
        RECT 4.000 430.800 996.000 439.600 ;
        RECT 4.000 429.400 995.600 430.800 ;
        RECT 4.000 417.200 996.000 429.400 ;
        RECT 4.400 415.800 996.000 417.200 ;
        RECT 4.000 407.680 996.000 415.800 ;
        RECT 4.000 406.280 995.600 407.680 ;
        RECT 4.000 393.400 996.000 406.280 ;
        RECT 4.400 392.000 996.000 393.400 ;
        RECT 4.000 384.560 996.000 392.000 ;
        RECT 4.000 383.160 995.600 384.560 ;
        RECT 4.000 369.600 996.000 383.160 ;
        RECT 4.400 368.200 996.000 369.600 ;
        RECT 4.000 361.440 996.000 368.200 ;
        RECT 4.000 360.040 995.600 361.440 ;
        RECT 4.000 345.800 996.000 360.040 ;
        RECT 4.400 344.400 996.000 345.800 ;
        RECT 4.000 338.320 996.000 344.400 ;
        RECT 4.000 336.920 995.600 338.320 ;
        RECT 4.000 322.000 996.000 336.920 ;
        RECT 4.400 320.600 996.000 322.000 ;
        RECT 4.000 315.200 996.000 320.600 ;
        RECT 4.000 313.800 995.600 315.200 ;
        RECT 4.000 298.200 996.000 313.800 ;
        RECT 4.400 296.800 996.000 298.200 ;
        RECT 4.000 292.080 996.000 296.800 ;
        RECT 4.000 290.680 995.600 292.080 ;
        RECT 4.000 274.400 996.000 290.680 ;
        RECT 4.400 273.000 996.000 274.400 ;
        RECT 4.000 268.960 996.000 273.000 ;
        RECT 4.000 267.560 995.600 268.960 ;
        RECT 4.000 250.600 996.000 267.560 ;
        RECT 4.400 249.200 996.000 250.600 ;
        RECT 4.000 245.840 996.000 249.200 ;
        RECT 4.000 244.440 995.600 245.840 ;
        RECT 4.000 226.800 996.000 244.440 ;
        RECT 4.400 225.400 996.000 226.800 ;
        RECT 4.000 222.720 996.000 225.400 ;
        RECT 4.000 221.320 995.600 222.720 ;
        RECT 4.000 203.000 996.000 221.320 ;
        RECT 4.400 201.600 996.000 203.000 ;
        RECT 4.000 199.600 996.000 201.600 ;
        RECT 4.000 198.200 995.600 199.600 ;
        RECT 4.000 179.200 996.000 198.200 ;
        RECT 4.400 177.800 996.000 179.200 ;
        RECT 4.000 176.480 996.000 177.800 ;
        RECT 4.000 175.080 995.600 176.480 ;
        RECT 4.000 155.400 996.000 175.080 ;
        RECT 4.400 154.000 996.000 155.400 ;
        RECT 4.000 153.360 996.000 154.000 ;
        RECT 4.000 151.960 995.600 153.360 ;
        RECT 4.000 131.600 996.000 151.960 ;
        RECT 4.400 130.240 996.000 131.600 ;
        RECT 4.400 130.200 995.600 130.240 ;
        RECT 4.000 128.840 995.600 130.200 ;
        RECT 4.000 107.800 996.000 128.840 ;
        RECT 4.400 107.120 996.000 107.800 ;
        RECT 4.400 106.400 995.600 107.120 ;
        RECT 4.000 105.720 995.600 106.400 ;
        RECT 4.000 84.000 996.000 105.720 ;
        RECT 4.400 82.600 995.600 84.000 ;
        RECT 4.000 60.880 996.000 82.600 ;
        RECT 4.000 60.200 995.600 60.880 ;
        RECT 4.400 59.480 995.600 60.200 ;
        RECT 4.400 58.800 996.000 59.480 ;
        RECT 4.000 37.760 996.000 58.800 ;
        RECT 4.000 36.400 995.600 37.760 ;
        RECT 4.400 36.360 995.600 36.400 ;
        RECT 4.400 35.000 996.000 36.360 ;
        RECT 4.000 14.640 996.000 35.000 ;
        RECT 4.000 13.240 995.600 14.640 ;
        RECT 4.000 12.600 996.000 13.240 ;
        RECT 4.400 11.200 996.000 12.600 ;
        RECT 4.000 0.175 996.000 11.200 ;
      LAYER met4 ;
        RECT 8.575 10.240 20.640 986.505 ;
        RECT 23.040 10.240 97.440 986.505 ;
        RECT 99.840 10.240 174.240 986.505 ;
        RECT 176.640 10.240 251.040 986.505 ;
        RECT 253.440 10.240 327.840 986.505 ;
        RECT 330.240 10.240 404.640 986.505 ;
        RECT 407.040 10.240 481.440 986.505 ;
        RECT 483.840 10.240 558.240 986.505 ;
        RECT 560.640 10.240 635.040 986.505 ;
        RECT 637.440 10.240 711.840 986.505 ;
        RECT 714.240 10.240 788.640 986.505 ;
        RECT 791.040 10.240 807.465 986.505 ;
        RECT 8.575 0.175 807.465 10.240 ;
  END
END wrapped_tms1x00
END LIBRARY

