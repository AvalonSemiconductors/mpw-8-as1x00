* NGSPICE file created from wrapped_tms1x00.ext - technology: sky130B

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_4 abstract view
.subckt sky130_fd_sc_hd__nor4b_4 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

.subckt wrapped_tms1x00 io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ oram_addr[0] oram_addr[1] oram_addr[2] oram_addr[3] oram_addr[4] oram_addr[5] oram_addr[6]
+ oram_addr[7] oram_addr[8] oram_csb oram_value[0] oram_value[10] oram_value[11] oram_value[12]
+ oram_value[13] oram_value[14] oram_value[15] oram_value[16] oram_value[17] oram_value[18]
+ oram_value[19] oram_value[1] oram_value[20] oram_value[21] oram_value[22] oram_value[23]
+ oram_value[24] oram_value[25] oram_value[26] oram_value[27] oram_value[28] oram_value[29]
+ oram_value[2] oram_value[30] oram_value[31] oram_value[3] oram_value[4] oram_value[5]
+ oram_value[6] oram_value[7] oram_value[8] oram_value[9] ram_adrb[0] ram_adrb[1]
+ ram_adrb[2] ram_adrb[3] ram_adrb[4] ram_adrb[5] ram_adrb[6] ram_adrb[7] ram_adrb[8]
+ ram_csb ram_val[0] ram_val[10] ram_val[11] ram_val[12] ram_val[13] ram_val[14] ram_val[15]
+ ram_val[16] ram_val[17] ram_val[18] ram_val[19] ram_val[1] ram_val[20] ram_val[21]
+ ram_val[22] ram_val[23] ram_val[24] ram_val[25] ram_val[26] ram_val[27] ram_val[28]
+ ram_val[29] ram_val[2] ram_val[30] ram_val[31] ram_val[3] ram_val[4] ram_val[5]
+ ram_val[6] ram_val[7] ram_val[8] ram_val[9] ram_web vccd1 vssd1 wb_clk_i wb_rst_i
+ wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14]
+ wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1]
+ wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25]
+ wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30]
+ wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8]
+ wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13]
+ wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19]
+ wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24]
+ wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2]
+ wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6]
+ wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11]
+ wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17]
+ wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22]
+ wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28]
+ wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4]
+ wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_stb_i wbs_we_i
XFILLER_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2574__S0 _0799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2479__B1 _0813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3155_ tms1x00.RAM\[105\]\[1\] _1328_ _1425_ vssd1 vssd1 vccd1 vccd1 _1427_ sky130_fd_sc_hd__mux2_1
X_3086_ _1361_ tms1x00.RAM\[112\]\[0\] _1386_ vssd1 vssd1 vccd1 vccd1 _1387_ sky130_fd_sc_hd__mux2_1
XFILLER_54_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3985__S _0724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3988_ net12 _1899_ vssd1 vssd1 vccd1 vccd1 _1906_ sky130_fd_sc_hd__or2_1
XFILLER_10_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4878__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2939_ _1294_ vssd1 vssd1 vccd1 vccd1 _0088_ sky130_fd_sc_hd__clkbuf_1
XFILLER_22_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3903__A0 _1821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4609_ clknet_leaf_3_wb_clk_i _0230_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[24\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_77_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2565__S0 _0955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5033__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3122__A1 _1334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4960_ clknet_leaf_9_wb_clk_i _0570_ vssd1 vssd1 vccd1 vccd1 tms1x00.P\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_33_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3911_ _1862_ vssd1 vssd1 vccd1 vccd1 _0492_ sky130_fd_sc_hd__clkbuf_1
X_4891_ clknet_leaf_2_wb_clk_i _0505_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[90\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_3842_ _1823_ tms1x00.RAM\[83\]\[3\] _1817_ vssd1 vssd1 vccd1 vccd1 _1824_ sky130_fd_sc_hd__mux2_1
X_3773_ tms1x00.RAM\[73\]\[2\] _1777_ _1781_ vssd1 vssd1 vccd1 vccd1 _1784_ sky130_fd_sc_hd__mux2_1
XANTENNA__2722__B _1112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2724_ _0944_ _1108_ _1110_ _0804_ _1114_ vssd1 vssd1 vccd1 vccd1 _1115_ sky130_fd_sc_hd__a311o_1
X_2655_ _0975_ tms1x00.RAM\[54\]\[2\] _0977_ vssd1 vssd1 vccd1 vccd1 _1046_ sky130_fd_sc_hd__o21a_1
X_4325_ _2143_ vssd1 vssd1 vccd1 vccd1 _0625_ sky130_fd_sc_hd__clkbuf_1
X_2586_ _0975_ tms1x00.RAM\[118\]\[1\] _0977_ vssd1 vssd1 vccd1 vccd1 _0978_ sky130_fd_sc_hd__o21a_1
X_4256_ tms1x00.RAM\[119\]\[3\] _1333_ _2101_ vssd1 vssd1 vccd1 vccd1 _2105_ sky130_fd_sc_hd__mux2_1
XFILLER_74_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4187_ tms1x00.PC\[4\] _2048_ _2054_ vssd1 vssd1 vccd1 vccd1 _2055_ sky130_fd_sc_hd__a21oi_1
X_3207_ _1323_ vssd1 vssd1 vccd1 vccd1 _1456_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__2872__A0 _0912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4550__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3138_ _1417_ vssd1 vssd1 vccd1 vccd1 _0164_ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4074__C1 _1966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3069_ _1377_ vssd1 vssd1 vccd1 vccd1 _0135_ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4377__A0 tms1x00.PC\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3728__B _1337_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2927__A1 _1235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2786__S0 _0924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4301__A0 _1823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4294__B _1345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3040__A0 _1130_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4423__CLK clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2440_ _0825_ _0829_ _0832_ _0807_ _0775_ vssd1 vssd1 vccd1 vccd1 _0833_ sky130_fd_sc_hd__o221a_1
XFILLER_5_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2371_ _0718_ vssd1 vssd1 vccd1 vccd1 _0766_ sky130_fd_sc_hd__clkbuf_4
XFILLER_69_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4110_ _1992_ vssd1 vssd1 vccd1 vccd1 _0561_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4573__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2551__C1 _0942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4041_ _0732_ _0763_ _1922_ net88 vssd1 vssd1 vccd1 vccd1 _1944_ sky130_fd_sc_hd__a31o_1
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_4_wb_clk_i_A clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__2209__S _0668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4943_ clknet_leaf_7_wb_clk_i _0553_ vssd1 vssd1 vccd1 vccd1 tms1x00.SR\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_32_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4874_ clknet_leaf_15_wb_clk_i _0488_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[94\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_3825_ tms1x00.RAM\[84\]\[1\] _1775_ _1811_ vssd1 vssd1 vccd1 vccd1 _1813_ sky130_fd_sc_hd__mux2_1
XANTENNA__3031__A0 _1130_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3756_ _1237_ _1403_ vssd1 vssd1 vccd1 vccd1 _1773_ sky130_fd_sc_hd__nor2_2
X_2707_ tms1x00.RAM\[79\]\[2\] _0830_ vssd1 vssd1 vccd1 vccd1 _1098_ sky130_fd_sc_hd__or2b_1
X_3687_ _1734_ vssd1 vssd1 vccd1 vccd1 _0396_ sky130_fd_sc_hd__clkbuf_1
X_2638_ _0960_ _0983_ _1029_ vssd1 vssd1 vccd1 vccd1 _1030_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2569_ tms1x00.RAM\[100\]\[1\] tms1x00.RAM\[101\]\[1\] tms1x00.RAM\[102\]\[1\] tms1x00.RAM\[103\]\[1\]
+ _0945_ _0791_ vssd1 vssd1 vccd1 vccd1 _0961_ sky130_fd_sc_hd__mux4_1
X_4308_ tms1x00.RAM\[20\]\[2\] _1330_ _2131_ vssd1 vssd1 vccd1 vccd1 _2134_ sky130_fd_sc_hd__mux2_1
XFILLER_75_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4239_ _2095_ vssd1 vssd1 vccd1 vccd1 _0587_ sky130_fd_sc_hd__clkbuf_1
XFILLER_47_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2643__A _1034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3270__A0 _1485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2362__B tms1x00.ins_in\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4446__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3022__A0 _1130_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4596__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input55_A wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2836__A0 _1225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3261__A0 _1488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2553__A _0808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4590_ clknet_leaf_14_wb_clk_i _0211_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[115\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_3610_ tms1x00.RAM\[55\]\[1\] _1672_ _1688_ vssd1 vssd1 vccd1 vccd1 _1690_ sky130_fd_sc_hd__mux2_1
X_3541_ tms1x00.RAM\[53\]\[0\] _1571_ _1649_ vssd1 vssd1 vccd1 vccd1 _1650_ sky130_fd_sc_hd__mux2_1
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3472_ _1611_ vssd1 vssd1 vccd1 vccd1 _0304_ sky130_fd_sc_hd__clkbuf_1
X_2423_ _0815_ vssd1 vssd1 vccd1 vccd1 _0816_ sky130_fd_sc_hd__buf_6
X_2354_ _0747_ _0748_ tms1x00.ins_in\[5\] vssd1 vssd1 vccd1 vccd1 _0749_ sky130_fd_sc_hd__or3_1
XFILLER_69_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2728__A _0921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2285_ _0699_ vssd1 vssd1 vccd1 vccd1 _0704_ sky130_fd_sc_hd__buf_2
XFILLER_65_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4024_ tms1x00.Y\[2\] _1918_ vssd1 vssd1 vccd1 vccd1 _1932_ sky130_fd_sc_hd__nand2_1
XFILLER_49_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4469__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3252__A0 _1366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4926_ clknet_leaf_14_wb_clk_i _0536_ vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__dfxtp_2
XFILLER_61_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3278__B _1261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4857_ clknet_leaf_23_wb_clk_i _0471_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[86\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3808_ _1803_ vssd1 vssd1 vccd1 vccd1 _0448_ sky130_fd_sc_hd__clkbuf_1
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4788_ clknet_leaf_24_wb_clk_i _0402_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[72\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3739_ _1763_ vssd1 vssd1 vccd1 vccd1 _0419_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__2763__C1 _0802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2357__B _0742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2818__B1 _0821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3491__A0 _1590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3916__B _1409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2548__A _0819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3379__A _1229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4761__CLK clknet_leaf_20_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2972_ _1314_ vssd1 vssd1 vccd1 vccd1 _0101_ sky130_fd_sc_hd__clkbuf_1
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4711_ clknet_leaf_5_wb_clk_i _0325_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[47\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_4642_ clknet_leaf_1_wb_clk_i _0263_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[36\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_4573_ clknet_leaf_32_wb_clk_i _0194_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[120\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_3524_ _1640_ vssd1 vssd1 vccd1 vccd1 _0327_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__2745__C1 _0776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3455_ _1590_ tms1x00.RAM\[45\]\[2\] _1599_ vssd1 vssd1 vccd1 vccd1 _1602_ sky130_fd_sc_hd__mux2_1
X_2406_ _0777_ vssd1 vssd1 vccd1 vccd1 _0799_ sky130_fd_sc_hd__clkbuf_16
XFILLER_69_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3386_ _1492_ tms1x00.RAM\[35\]\[3\] _1556_ vssd1 vssd1 vccd1 vccd1 _1560_ sky130_fd_sc_hd__mux2_1
XFILLER_57_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2337_ tms1x00.X\[0\] tms1x00.ram_addr_buff\[5\] _0726_ vssd1 vssd1 vccd1 vccd1 _0736_
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2268_ _0701_ _0698_ _0700_ wbs_o_buff\[5\] vssd1 vssd1 vccd1 vccd1 _0030_ sky130_fd_sc_hd__a22o_1
X_4007_ _0755_ _0739_ _0763_ _1918_ vssd1 vssd1 vccd1 vccd1 _1919_ sky130_fd_sc_hd__and4_1
XANTENNA__2276__A1 net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2199_ _0666_ vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__clkbuf_1
XFILLER_25_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4017__A2 _0730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2905__B _1273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4909_ clknet_leaf_8_wb_clk_i _0523_ vssd1 vssd1 vccd1 vccd1 tms1x00.ins_in\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2200__A1 wbs_o_buff\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4634__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input18_A ram_val[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3464__A0 _1590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_14_wb_clk_i clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output86_A net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3240_ _1476_ vssd1 vssd1 vccd1 vccd1 _0207_ sky130_fd_sc_hd__clkbuf_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3171_ _1286_ _1430_ vssd1 vssd1 vccd1 vccd1 _1436_ sky130_fd_sc_hd__nor2_2
XFILLER_67_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3455__A0 _1590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2217__S _0668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2955_ _0914_ _1303_ vssd1 vssd1 vccd1 vccd1 _1304_ sky130_fd_sc_hd__nor2_2
XANTENNA__4507__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2886_ tms1x00.RAM\[89\]\[0\] _1235_ _1262_ vssd1 vssd1 vccd1 vccd1 _1263_ sky130_fd_sc_hd__mux2_1
X_4625_ clknet_leaf_6_wb_clk_i _0246_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[32\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_4556_ clknet_leaf_9_wb_clk_i _0177_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[124\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4657__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3507_ _1588_ tms1x00.RAM\[48\]\[1\] _1629_ vssd1 vssd1 vccd1 vccd1 _1631_ sky130_fd_sc_hd__mux2_1
XANTENNA__2194__A0 net42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3930__A1 _1777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4487_ clknet_leaf_30_wb_clk_i _0108_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[101\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_3438_ _1224_ vssd1 vssd1 vccd1 vccd1 _1592_ sky130_fd_sc_hd__buf_2
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2497__A1 _0798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3369_ _1550_ vssd1 vssd1 vccd1 vccd1 _0262_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__2592__S1 _0791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5039_ clknet_leaf_4_wb_clk_i _0649_ vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__dfxtp_1
XANTENNA__3446__A0 tms1x00.RAM\[38\]\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2354__C tms1x00.ins_in\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3749__A1 _1672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2421__A1 _0789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4174__A1 tms1x00.ins_in\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2724__A2 _1108_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput75 net75 vssd1 vssd1 vccd1 vccd1 io_out[16] sky130_fd_sc_hd__buf_2
Xoutput86 net86 vssd1 vssd1 vccd1 vccd1 io_out[27] sky130_fd_sc_hd__buf_2
XFILLER_1_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput97 net97 vssd1 vssd1 vccd1 vccd1 oram_addr[2] sky130_fd_sc_hd__buf_2
XFILLER_49_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2488__B2 _0807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2740_ _1130_ tms1x00.RAM\[109\]\[2\] _0918_ vssd1 vssd1 vccd1 vccd1 _1131_ sky130_fd_sc_hd__mux2_1
XANTENNA__2561__A _0794_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2412__A1 _0776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2671_ _0932_ _1061_ vssd1 vssd1 vccd1 vccd1 _1062_ sky130_fd_sc_hd__and2_1
XFILLER_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4410_ clknet_leaf_28_wb_clk_i _0008_ vssd1 vssd1 vccd1 vccd1 wbs_o_buff\[14\] sky130_fd_sc_hd__dfxtp_1
X_4341_ _2152_ vssd1 vssd1 vccd1 vccd1 _0632_ sky130_fd_sc_hd__clkbuf_1
X_4272_ tms1x00.RAM\[22\]\[2\] _1330_ _2111_ vssd1 vssd1 vccd1 vccd1 _2114_ sky130_fd_sc_hd__mux2_1
XANTENNA__2479__A1 _0789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3223_ tms1x00.RAM\[118\]\[1\] _1459_ _1465_ vssd1 vssd1 vccd1 vccd1 _1467_ sky130_fd_sc_hd__mux2_1
XTAP_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3154_ _1426_ vssd1 vssd1 vccd1 vccd1 _0171_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__2574__S1 _0813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2736__A _0748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3085_ _1345_ _1375_ vssd1 vssd1 vccd1 vccd1 _1386_ sky130_fd_sc_hd__or2_2
XFILLER_39_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3987_ _1905_ vssd1 vssd1 vccd1 vccd1 _0525_ sky130_fd_sc_hd__clkbuf_1
XFILLER_50_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3567__A _1240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2938_ _1035_ tms1x00.RAM\[49\]\[1\] _1292_ vssd1 vssd1 vccd1 vccd1 _1294_ sky130_fd_sc_hd__mux2_1
XFILLER_31_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2403__A1 _0787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4156__A1 _0768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2869_ _1249_ vssd1 vssd1 vccd1 vccd1 _1250_ sky130_fd_sc_hd__buf_4
X_4608_ clknet_leaf_4_wb_clk_i _0229_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[24\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_4539_ clknet_leaf_14_wb_clk_i _0160_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[108\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2565__S1 _0956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2890__A1 _1245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4822__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2381__A _0038_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3477__A _1403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4972__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2556__A _0783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3910_ _1819_ tms1x00.RAM\[93\]\[1\] _1860_ vssd1 vssd1 vccd1 vccd1 _1862_ sky130_fd_sc_hd__mux2_1
XANTENNA__2633__A1 tms1x00.RAM\[49\]\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4890_ clknet_leaf_30_wb_clk_i _0504_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[90\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_3841_ _1224_ vssd1 vssd1 vccd1 vccd1 _1823_ sky130_fd_sc_hd__clkbuf_4
XFILLER_32_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3772_ _1783_ vssd1 vssd1 vccd1 vccd1 _0432_ sky130_fd_sc_hd__clkbuf_1
X_2723_ _0996_ _1111_ _1113_ _0806_ vssd1 vssd1 vccd1 vccd1 _1114_ sky130_fd_sc_hd__o211a_1
XFILLER_9_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2654_ tms1x00.RAM\[55\]\[2\] _0975_ vssd1 vssd1 vccd1 vccd1 _1045_ sky130_fd_sc_hd__or2b_1
X_2585_ _0850_ vssd1 vssd1 vccd1 vccd1 _0977_ sky130_fd_sc_hd__buf_6
XANTENNA__4011__A tms1x00.Y\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4324_ _1819_ tms1x00.RAM\[127\]\[1\] _2141_ vssd1 vssd1 vccd1 vccd1 _2143_ sky130_fd_sc_hd__mux2_1
XFILLER_68_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4255_ _2104_ vssd1 vssd1 vccd1 vccd1 _0594_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4186_ tms1x00.PC\[5\] _2030_ _2053_ vssd1 vssd1 vccd1 vccd1 _2054_ sky130_fd_sc_hd__o21ai_1
XFILLER_28_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3206_ _1455_ vssd1 vssd1 vccd1 vccd1 _0194_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4310__A1 _1333_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3137_ tms1x00.RAM\[107\]\[1\] _1328_ _1415_ vssd1 vssd1 vccd1 vccd1 _1417_ sky130_fd_sc_hd__mux2_1
XFILLER_82_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3068_ _1361_ tms1x00.RAM\[114\]\[0\] _1376_ vssd1 vssd1 vccd1 vccd1 _1377_ sky130_fd_sc_hd__mux2_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4377__A1 net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4995__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2786__S1 _0928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2863__A1 _1245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3000__A _1333_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5000__CLK clknet_leaf_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2370_ _0755_ _0756_ _0764_ net77 vssd1 vssd1 vccd1 vccd1 _0765_ sky130_fd_sc_hd__a31o_1
XFILLER_69_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4040_ _0753_ _1942_ _1943_ _1931_ vssd1 vssd1 vccd1 vccd1 _0540_ sky130_fd_sc_hd__o211a_1
XFILLER_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4868__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4056__B1 net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4942_ clknet_leaf_7_wb_clk_i _0552_ vssd1 vssd1 vccd1 vccd1 tms1x00.status sky130_fd_sc_hd__dfxtp_1
XANTENNA__2606__A1 _0787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4873_ clknet_leaf_15_wb_clk_i _0487_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[94\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3824_ _1812_ vssd1 vssd1 vccd1 vccd1 _0455_ sky130_fd_sc_hd__clkbuf_1
X_3755_ _0911_ vssd1 vssd1 vccd1 vccd1 _1772_ sky130_fd_sc_hd__clkbuf_4
X_3686_ _1706_ tms1x00.RAM\[64\]\[1\] _1732_ vssd1 vssd1 vccd1 vccd1 _1734_ sky130_fd_sc_hd__mux2_1
X_2706_ tms1x00.RAM\[72\]\[2\] tms1x00.RAM\[73\]\[2\] tms1x00.RAM\[74\]\[2\] tms1x00.RAM\[75\]\[2\]
+ _0873_ _0822_ vssd1 vssd1 vccd1 vccd1 _1097_ sky130_fd_sc_hd__mux4_1
X_2637_ _0040_ _0993_ _1007_ _1028_ _0835_ vssd1 vssd1 vccd1 vccd1 _1029_ sky130_fd_sc_hd__o311a_1
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2542__B1 _0776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2568_ _0920_ _0935_ _0943_ _0040_ _0959_ vssd1 vssd1 vccd1 vccd1 _0960_ sky130_fd_sc_hd__a311o_1
XFILLER_59_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2499_ _0797_ _0891_ vssd1 vssd1 vccd1 vccd1 _0892_ sky130_fd_sc_hd__or2_1
XANTENNA__3580__A _1034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4307_ _2133_ vssd1 vssd1 vccd1 vccd1 _0617_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4295__A0 _1816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4238_ tms1x00.N\[3\] _2007_ vssd1 vssd1 vccd1 vccd1 _2095_ sky130_fd_sc_hd__or2_1
XFILLER_59_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4169_ tms1x00.PC\[2\] _2030_ _2039_ _1971_ vssd1 vssd1 vccd1 vccd1 _2040_ sky130_fd_sc_hd__o22a_1
XANTENNA__4047__B1 net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3755__A _0911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input48_A wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3665__A _1237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3540_ _1240_ _1284_ vssd1 vssd1 vccd1 vccd1 _1649_ sky130_fd_sc_hd__nor2_2
XFILLER_6_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3471_ tms1x00.RAM\[43\]\[1\] _1574_ _1609_ vssd1 vssd1 vccd1 vccd1 _1611_ sky130_fd_sc_hd__mux2_1
X_2422_ _0035_ vssd1 vssd1 vccd1 vccd1 _0815_ sky130_fd_sc_hd__buf_8
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2353_ tms1x00.ins_in\[6\] vssd1 vssd1 vccd1 vccd1 _0748_ sky130_fd_sc_hd__clkbuf_4
X_4023_ net82 _1929_ _1930_ _1931_ vssd1 vssd1 vccd1 vccd1 _0535_ sky130_fd_sc_hd__o211a_1
XANTENNA__2728__B _1118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4277__A0 _1816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2284_ net88 _0702_ _0703_ wbs_o_buff\[19\] vssd1 vssd1 vccd1 vccd1 _0013_ sky130_fd_sc_hd__a22o_1
XANTENNA__4029__B1 net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2744__A _0953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4925_ clknet_leaf_14_wb_clk_i _0535_ vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__dfxtp_2
XFILLER_40_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4856_ clknet_leaf_16_wb_clk_i _0470_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[81\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2460__C1 _0828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3807_ _1706_ tms1x00.RAM\[77\]\[1\] _1801_ vssd1 vssd1 vccd1 vccd1 _1803_ sky130_fd_sc_hd__mux2_1
XFILLER_20_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4787_ clknet_leaf_24_wb_clk_i _0401_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[72\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_3738_ _1703_ tms1x00.RAM\[76\]\[0\] _1762_ vssd1 vssd1 vccd1 vccd1 _1763_ sky130_fd_sc_hd__mux2_1
XFILLER_69_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3669_ _1724_ vssd1 vssd1 vccd1 vccd1 _0388_ sky130_fd_sc_hd__clkbuf_1
XFILLER_76_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3514__S _1634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2818__A1 _0944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4413__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3243__A1 _1461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2451__C1 _0775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2809__A1 _0920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2564__A _0800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3482__A1 _1576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3379__B _1525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2971_ tms1x00.RAM\[103\]\[2\] _1245_ _1311_ vssd1 vssd1 vccd1 vccd1 _1314_ sky130_fd_sc_hd__mux2_1
XANTENNA__3234__A1 _1461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4710_ clknet_leaf_4_wb_clk_i _0324_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[47\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4641_ clknet_leaf_1_wb_clk_i _0262_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[37\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_4572_ clknet_leaf_32_wb_clk_i _0193_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[120\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_3523_ _1585_ tms1x00.RAM\[46\]\[0\] _1639_ vssd1 vssd1 vccd1 vccd1 _1640_ sky130_fd_sc_hd__mux2_1
XFILLER_6_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3454_ _1601_ vssd1 vssd1 vccd1 vccd1 _0296_ sky130_fd_sc_hd__clkbuf_1
X_2405_ _0797_ vssd1 vssd1 vccd1 vccd1 _0798_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__2739__A _1129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3385_ _1559_ vssd1 vssd1 vccd1 vccd1 _0269_ sky130_fd_sc_hd__clkbuf_1
XFILLER_69_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4436__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2336_ _0735_ vssd1 vssd1 vccd1 vccd1 _0046_ sky130_fd_sc_hd__clkbuf_1
XFILLER_29_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2267_ net74 vssd1 vssd1 vccd1 vccd1 _0701_ sky130_fd_sc_hd__clkbuf_4
XFILLER_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4006_ tms1x00.Y\[0\] tms1x00.Y\[1\] vssd1 vssd1 vccd1 vccd1 _1918_ sky130_fd_sc_hd__and2b_1
XANTENNA__3473__A1 _1576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2198_ net44 wbs_o_buff\[8\] _0657_ vssd1 vssd1 vccd1 vccd1 _0666_ sky130_fd_sc_hd__mux2_1
XFILLER_52_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4586__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3225__A1 _1461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4908_ clknet_leaf_8_wb_clk_i _0522_ vssd1 vssd1 vccd1 vccd1 tms1x00.ins_in\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_40_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4839_ clknet_leaf_23_wb_clk_i _0453_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[85\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4929__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_28_wb_clk_i_A clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_71_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2323__S _0726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3943__A _1250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output79_A net79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2559__A _0818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3170_ _1435_ vssd1 vssd1 vccd1 vccd1 _0178_ sky130_fd_sc_hd__clkbuf_1
XFILLER_66_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2663__C1 _0802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2954_ _1302_ vssd1 vssd1 vccd1 vccd1 _1303_ sky130_fd_sc_hd__buf_6
XFILLER_31_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2885_ _1258_ _1261_ vssd1 vssd1 vccd1 vccd1 _1262_ sky130_fd_sc_hd__nor2_2
XANTENNA__4014__A _0732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4624_ clknet_leaf_6_wb_clk_i _0245_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[32\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_4555_ clknet_leaf_13_wb_clk_i _0176_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[124\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3853__A _1251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3391__A0 _1488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3506_ _1630_ vssd1 vssd1 vccd1 vccd1 _0319_ sky130_fd_sc_hd__clkbuf_1
X_4486_ clknet_leaf_30_wb_clk_i _0107_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[101\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_3437_ _1591_ vssd1 vssd1 vccd1 vccd1 _0289_ sky130_fd_sc_hd__clkbuf_1
XFILLER_66_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2497__A2 _0887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3368_ tms1x00.RAM\[37\]\[3\] _1463_ _1546_ vssd1 vssd1 vccd1 vccd1 _1550_ sky130_fd_sc_hd__mux2_1
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2319_ _0701_ _0720_ _0722_ vssd1 vssd1 vccd1 vccd1 _0723_ sky130_fd_sc_hd__and3b_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3299_ _1488_ tms1x00.RAM\[28\]\[1\] _1509_ vssd1 vssd1 vccd1 vccd1 _1511_ sky130_fd_sc_hd__mux2_1
X_5038_ clknet_leaf_5_wb_clk_i _0648_ vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__dfxtp_1
XANTENNA__3446__A1 _1576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4601__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3382__A0 _1488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2724__A3 _1110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput76 net76 vssd1 vssd1 vccd1 vccd1 io_out[17] sky130_fd_sc_hd__buf_2
XANTENNA__2379__A _0747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput87 net87 vssd1 vssd1 vccd1 vccd1 io_out[28] sky130_fd_sc_hd__buf_2
XFILLER_0_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput98 net98 vssd1 vssd1 vccd1 vccd1 oram_addr[3] sky130_fd_sc_hd__buf_2
XANTENNA__4751__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input30_A ram_val[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2660__A2 tms1x00.RAM\[62\]\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2670_ tms1x00.RAM\[30\]\[2\] tms1x00.RAM\[31\]\[2\] _0923_ vssd1 vssd1 vccd1 vccd1
+ _1061_ sky130_fd_sc_hd__mux2_1
XFILLER_9_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4340_ _1235_ tms1x00.RAM\[1\]\[0\] _2151_ vssd1 vssd1 vccd1 vccd1 _2152_ sky130_fd_sc_hd__mux2_1
X_4271_ _2113_ vssd1 vssd1 vccd1 vccd1 _0601_ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3222_ _1466_ vssd1 vssd1 vccd1 vccd1 _0199_ sky130_fd_sc_hd__clkbuf_1
XFILLER_79_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3153_ tms1x00.RAM\[105\]\[0\] _1324_ _1425_ vssd1 vssd1 vccd1 vccd1 _1426_ sky130_fd_sc_hd__mux2_1
XFILLER_39_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3084_ _1385_ vssd1 vssd1 vccd1 vccd1 _0142_ sky130_fd_sc_hd__clkbuf_1
XFILLER_82_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2651__A2 tms1x00.RAM\[38\]\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3986_ net103 _1904_ vssd1 vssd1 vccd1 vccd1 _1905_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout148_A net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4624__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2937_ _1293_ vssd1 vssd1 vccd1 vccd1 _0087_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__3567__B _1344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2868_ tms1x00.ram_addr_buff\[5\] tms1x00.ram_addr_buff\[6\] tms1x00.ram_addr_buff\[4\]
+ vssd1 vssd1 vccd1 vccd1 _1249_ sky130_fd_sc_hd__or3b_4
X_4607_ clknet_leaf_4_wb_clk_i _0228_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[24\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_2799_ _0818_ _1188_ _0794_ vssd1 vssd1 vccd1 vccd1 _1189_ sky130_fd_sc_hd__a21o_1
XANTENNA__3583__A _1129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4774__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4538_ clknet_leaf_14_wb_clk_i _0159_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[108\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4469_ clknet_leaf_10_wb_clk_i _0090_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[49\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3477__B _1525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3355__A0 _1488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3107__A0 _1364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4647__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3840_ _1822_ vssd1 vssd1 vccd1 vccd1 _0461_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__2572__A _0948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4263__S _2106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3771_ tms1x00.RAM\[73\]\[1\] _1775_ _1781_ vssd1 vssd1 vccd1 vccd1 _1783_ sky130_fd_sc_hd__mux2_1
X_2722_ _0783_ _1112_ vssd1 vssd1 vccd1 vccd1 _1113_ sky130_fd_sc_hd__or2_1
XFILLER_9_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4797__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4138__A2 _2007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3346__A0 _1488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2653_ _0948_ _1041_ _1043_ _0776_ vssd1 vssd1 vccd1 vccd1 _1044_ sky130_fd_sc_hd__o211a_1
X_2584_ tms1x00.RAM\[119\]\[1\] _0975_ vssd1 vssd1 vccd1 vccd1 _0976_ sky130_fd_sc_hd__or2b_1
X_4323_ _2142_ vssd1 vssd1 vccd1 vccd1 _0624_ sky130_fd_sc_hd__clkbuf_1
X_4254_ tms1x00.RAM\[119\]\[2\] _1330_ _2101_ vssd1 vssd1 vccd1 vccd1 _2104_ sky130_fd_sc_hd__mux2_1
XFILLER_68_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2747__A _0928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4185_ tms1x00.SR\[5\] _1971_ _2027_ vssd1 vssd1 vccd1 vccd1 _2053_ sky130_fd_sc_hd__or3_1
X_3205_ tms1x00.RAM\[120\]\[3\] _1334_ _1451_ vssd1 vssd1 vccd1 vccd1 _1455_ sky130_fd_sc_hd__mux2_1
XFILLER_82_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3136_ _1416_ vssd1 vssd1 vccd1 vccd1 _0163_ sky130_fd_sc_hd__clkbuf_1
XFILLER_82_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3067_ _1273_ _1375_ vssd1 vssd1 vccd1 vccd1 _1376_ sky130_fd_sc_hd__or2_2
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3969_ net93 _1893_ _0738_ vssd1 vssd1 vccd1 vccd1 _1894_ sky130_fd_sc_hd__mux2_1
XFILLER_6_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3337__A0 _1488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2376__B tms1x00.ins_in\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3328__A0 _1488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4112__A net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2551__A1 _0922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2362__C_N _0742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4941_ clknet_leaf_6_wb_clk_i _0551_ vssd1 vssd1 vccd1 vccd1 tms1x00.CL sky130_fd_sc_hd__dfxtp_1
XFILLER_32_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4872_ clknet_leaf_23_wb_clk_i _0486_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[87\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3823_ tms1x00.RAM\[84\]\[0\] _1772_ _1811_ vssd1 vssd1 vccd1 vccd1 _1812_ sky130_fd_sc_hd__mux2_1
XANTENNA__4006__B tms1x00.Y\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_9_wb_clk_i clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_3754_ _1771_ vssd1 vssd1 vccd1 vccd1 _0426_ sky130_fd_sc_hd__clkbuf_1
X_3685_ _1733_ vssd1 vssd1 vccd1 vccd1 _0395_ sky130_fd_sc_hd__clkbuf_1
X_2705_ _1092_ _1094_ _1095_ _0798_ _0775_ vssd1 vssd1 vccd1 vccd1 _1096_ sky130_fd_sc_hd__o221a_1
XANTENNA__4022__A _0718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2636_ _0773_ _1016_ _1027_ vssd1 vssd1 vccd1 vccd1 _1028_ sky130_fd_sc_hd__or3b_1
XANTENNA__2542__A1 _0922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2567_ _0944_ _0949_ _0958_ _0920_ vssd1 vssd1 vccd1 vccd1 _0959_ sky130_fd_sc_hd__a211oi_1
X_2498_ tms1x00.RAM\[56\]\[0\] tms1x00.RAM\[57\]\[0\] tms1x00.RAM\[58\]\[0\] tms1x00.RAM\[59\]\[0\]
+ _0777_ _0779_ vssd1 vssd1 vccd1 vccd1 _0891_ sky130_fd_sc_hd__mux4_1
X_4306_ tms1x00.RAM\[20\]\[1\] _1327_ _2131_ vssd1 vssd1 vccd1 vccd1 _2133_ sky130_fd_sc_hd__mux2_1
XFILLER_75_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4237_ _2094_ vssd1 vssd1 vccd1 vccd1 _0586_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4812__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2477__A _0807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4168_ tms1x00.ins_in\[4\] _1995_ _2027_ tms1x00.SR\[2\] vssd1 vssd1 vccd1 vccd1
+ _2039_ sky130_fd_sc_hd__o22a_1
XFILLER_56_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4099_ tms1x00.SR\[5\] tms1x00.PC\[5\] _1979_ vssd1 vssd1 vccd1 vccd1 _1985_ sky130_fd_sc_hd__mux2_1
XFILLER_56_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3119_ _1406_ vssd1 vssd1 vccd1 vccd1 _0156_ sky130_fd_sc_hd__clkbuf_1
XFILLER_70_325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2230__A0 net29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2387__A _0779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4286__A1 _1323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2326__S _0726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2850__A _0911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3665__B _1273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3470_ _1610_ vssd1 vssd1 vccd1 vccd1 _0303_ sky130_fd_sc_hd__clkbuf_1
X_2421_ _0789_ tms1x00.RAM\[78\]\[0\] _0813_ vssd1 vssd1 vccd1 vccd1 _0814_ sky130_fd_sc_hd__o21a_1
XFILLER_69_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2352_ tms1x00.ins_in\[7\] vssd1 vssd1 vccd1 vccd1 _0747_ sky130_fd_sc_hd__clkbuf_4
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2283_ net87 _0702_ _0703_ wbs_o_buff\[18\] vssd1 vssd1 vccd1 vccd1 _0012_ sky130_fd_sc_hd__a22o_1
X_4022_ _0718_ vssd1 vssd1 vccd1 vccd1 _1931_ sky130_fd_sc_hd__clkbuf_4
XFILLER_56_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4985__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2288__B1 _0704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4924_ clknet_leaf_13_wb_clk_i _0534_ vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__dfxtp_2
XFILLER_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4855_ clknet_leaf_16_wb_clk_i _0469_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[81\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3806_ _1802_ vssd1 vssd1 vccd1 vccd1 _0447_ sky130_fd_sc_hd__clkbuf_1
X_4786_ clknet_leaf_23_wb_clk_i _0400_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[72\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_3737_ _1236_ _1409_ vssd1 vssd1 vccd1 vccd1 _1762_ sky130_fd_sc_hd__or2_2
XANTENNA__2763__A1 _0798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4072__A_N _0742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3668_ _1706_ tms1x00.RAM\[66\]\[1\] _1722_ vssd1 vssd1 vccd1 vccd1 _1724_ sky130_fd_sc_hd__mux2_1
X_3599_ tms1x00.RAM\[56\]\[0\] _1669_ _1683_ vssd1 vssd1 vccd1 vccd1 _1684_ sky130_fd_sc_hd__mux2_1
X_2619_ _0807_ _1010_ _0802_ vssd1 vssd1 vccd1 vccd1 _1011_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4268__A1 _1323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2279__B1 _0703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_18_wb_clk_i_A clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__2935__A _1251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4708__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2203__A0 net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input60_A wbs_dat_i[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4259__A1 _1323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2970_ _1313_ vssd1 vssd1 vccd1 vccd1 _0100_ sky130_fd_sc_hd__clkbuf_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2993__A1 _1328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2580__A _0807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4640_ clknet_leaf_0_wb_clk_i _0261_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[37\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2745__A1 _0922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4571_ clknet_leaf_33_wb_clk_i _0192_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[120\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_3522_ _1396_ _1524_ vssd1 vssd1 vccd1 vccd1 _1639_ sky130_fd_sc_hd__or2_2
X_3453_ _1588_ tms1x00.RAM\[45\]\[1\] _1599_ vssd1 vssd1 vccd1 vccd1 _1601_ sky130_fd_sc_hd__mux2_1
XFILLER_6_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5013__CLK clknet_leaf_20_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2404_ _0037_ vssd1 vssd1 vccd1 vccd1 _0797_ sky130_fd_sc_hd__buf_2
XFILLER_69_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3384_ _1490_ tms1x00.RAM\[35\]\[2\] _1556_ vssd1 vssd1 vccd1 vccd1 _1559_ sky130_fd_sc_hd__mux2_1
XFILLER_58_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2335_ tms1x00.X\[2\] tms1x00.ram_addr_buff\[4\] _0726_ vssd1 vssd1 vccd1 vccd1 _0735_
+ sky130_fd_sc_hd__mux2_1
X_2266_ net73 _0698_ _0700_ wbs_o_buff\[4\] vssd1 vssd1 vccd1 vccd1 _0029_ sky130_fd_sc_hd__a22o_1
X_4005_ net78 _1916_ _1917_ _1901_ vssd1 vssd1 vccd1 vccd1 _0531_ sky130_fd_sc_hd__o211a_1
X_2197_ _0665_ vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__clkbuf_1
XFILLER_81_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4907_ clknet_leaf_8_wb_clk_i _0521_ vssd1 vssd1 vccd1 vccd1 tms1x00.ins_in\[1\]
+ sky130_fd_sc_hd__dfxtp_2
X_4838_ clknet_leaf_23_wb_clk_i _0452_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[85\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2984__A1 _1247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3586__A _1224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4769_ clknet_leaf_18_wb_clk_i _0383_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[67\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3525__S _1639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4680__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5036__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3943__B _1310_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4120__A net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_23_wb_clk_i clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__2575__A _0798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2294__B _0704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2953_ tms1x00.ram_addr_buff\[0\] tms1x00.ram_addr_buff\[1\] _1259_ vssd1 vssd1 vccd1
+ vccd1 _1302_ sky130_fd_sc_hd__or3_1
XFILLER_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2884_ _1260_ vssd1 vssd1 vccd1 vccd1 _1261_ sky130_fd_sc_hd__buf_6
X_4623_ clknet_leaf_8_wb_clk_i _0244_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[32\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_4554_ clknet_leaf_12_wb_clk_i _0175_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[124\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3853__B _1257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3505_ _1585_ tms1x00.RAM\[48\]\[0\] _1629_ vssd1 vssd1 vccd1 vccd1 _1630_ sky130_fd_sc_hd__mux2_1
X_4485_ clknet_leaf_29_wb_clk_i _0106_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[102\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_3436_ _1590_ tms1x00.RAM\[3\]\[2\] _1586_ vssd1 vssd1 vccd1 vccd1 _1591_ sky130_fd_sc_hd__mux2_1
XANTENNA__4340__A0 _1235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3367_ _1549_ vssd1 vssd1 vccd1 vccd1 _0261_ sky130_fd_sc_hd__clkbuf_1
XFILLER_57_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2318_ net148 _0721_ vssd1 vssd1 vccd1 vccd1 _0722_ sky130_fd_sc_hd__nand2_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3298_ _1510_ vssd1 vssd1 vccd1 vccd1 _0231_ sky130_fd_sc_hd__clkbuf_1
X_5037_ clknet_leaf_2_wb_clk_i _0647_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[9\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_73_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2249_ _0692_ vssd1 vssd1 vccd1 vccd1 tms1x00.K_in\[0\] sky130_fd_sc_hd__clkbuf_1
XFILLER_54_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2424__S _0816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2379__B _0748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4331__A0 _1235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput88 net88 vssd1 vssd1 vccd1 vccd1 io_out[29] sky130_fd_sc_hd__buf_2
Xoutput77 net77 vssd1 vssd1 vccd1 vccd1 io_out[18] sky130_fd_sc_hd__buf_2
XFILLER_76_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput99 net99 vssd1 vssd1 vccd1 vccd1 oram_addr[4] sky130_fd_sc_hd__buf_2
XFILLER_49_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input23_A ram_val[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2395__A _0777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2660__A3 tms1x00.RAM\[63\]\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3070__A0 _1364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output91_A net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3373__A1 _1459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2581__C1 _0806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4576__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4270_ tms1x00.RAM\[22\]\[1\] _1327_ _2111_ vssd1 vssd1 vccd1 vccd1 _2113_ sky130_fd_sc_hd__mux2_1
XFILLER_79_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4322__A0 _1816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3221_ tms1x00.RAM\[118\]\[0\] _1456_ _1465_ vssd1 vssd1 vccd1 vccd1 _1466_ sky130_fd_sc_hd__mux2_1
XFILLER_67_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3152_ _0914_ _1261_ vssd1 vssd1 vccd1 vccd1 _1425_ sky130_fd_sc_hd__nor2_2
X_3083_ _1368_ tms1x00.RAM\[113\]\[3\] _1381_ vssd1 vssd1 vccd1 vccd1 _1385_ sky130_fd_sc_hd__mux2_1
XFILLER_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3985_ tms1x00.ins_in\[5\] net11 _0724_ vssd1 vssd1 vccd1 vccd1 _1904_ sky130_fd_sc_hd__mux2_1
XFILLER_22_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2936_ _0912_ tms1x00.RAM\[49\]\[0\] _1292_ vssd1 vssd1 vccd1 vccd1 _1293_ sky130_fd_sc_hd__mux2_1
XANTENNA__2244__S net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2867_ _1248_ vssd1 vssd1 vccd1 vccd1 _0062_ sky130_fd_sc_hd__clkbuf_1
X_4606_ clknet_leaf_4_wb_clk_i _0227_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[24\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4919__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2798_ tms1x00.RAM\[4\]\[3\] tms1x00.RAM\[5\]\[3\] _0778_ vssd1 vssd1 vccd1 vccd1
+ _1188_ sky130_fd_sc_hd__mux2_1
XANTENNA__3364__A1 _1459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4537_ clknet_leaf_30_wb_clk_i _0158_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[10\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_4468_ clknet_leaf_10_wb_clk_i _0089_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[49\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4313__A0 _1816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3116__A1 _1324_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3419_ _1303_ _1525_ vssd1 vssd1 vccd1 vccd1 _1580_ sky130_fd_sc_hd__nor2_2
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4399_ clknet_leaf_35_wb_clk_i _0028_ vssd1 vssd1 vccd1 vccd1 wbs_o_buff\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3104__A _0913_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4077__C1 _1966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4006__A_N tms1x00.Y\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4449__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3052__A0 _1366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2329__S _0726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2853__A tms1x00.ram_addr_buff\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2572__B _0963_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3770_ _1782_ vssd1 vssd1 vccd1 vccd1 _0431_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__3594__A1 _1674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2721_ tms1x00.RAM\[120\]\[2\] tms1x00.RAM\[121\]\[2\] tms1x00.RAM\[122\]\[2\] tms1x00.RAM\[123\]\[2\]
+ _0823_ _0850_ vssd1 vssd1 vccd1 vccd1 _1112_ sky130_fd_sc_hd__mux4_1
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2652_ _0819_ _1042_ vssd1 vssd1 vccd1 vccd1 _1043_ sky130_fd_sc_hd__or2_1
XFILLER_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2583_ _0778_ vssd1 vssd1 vccd1 vccd1 _0975_ sky130_fd_sc_hd__clkbuf_8
X_4322_ _1816_ tms1x00.RAM\[127\]\[0\] _2141_ vssd1 vssd1 vccd1 vccd1 _2142_ sky130_fd_sc_hd__mux2_1
X_4253_ _2103_ vssd1 vssd1 vccd1 vccd1 _0593_ sky130_fd_sc_hd__clkbuf_1
X_3204_ _1454_ vssd1 vssd1 vccd1 vccd1 _0193_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4184_ _0760_ _2051_ _2052_ _1966_ vssd1 vssd1 vccd1 vccd1 _0575_ sky130_fd_sc_hd__o211a_1
XFILLER_67_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3135_ tms1x00.RAM\[107\]\[0\] _1324_ _1415_ vssd1 vssd1 vccd1 vccd1 _1416_ sky130_fd_sc_hd__mux2_1
XFILLER_67_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3066_ tms1x00.ram_addr_buff\[4\] tms1x00.ram_addr_buff\[5\] tms1x00.ram_addr_buff\[6\]
+ vssd1 vssd1 vccd1 vccd1 _1375_ sky130_fd_sc_hd__nand3_2
XANTENNA__2704__S0 _0840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3968_ net1 chip_sel_override net148 vssd1 vssd1 vccd1 vccd1 _1893_ sky130_fd_sc_hd__mux2_1
XFILLER_51_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4231__C1 _0766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2919_ _1281_ vssd1 vssd1 vccd1 vccd1 _0081_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4741__CLK clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3899_ _1816_ tms1x00.RAM\[94\]\[0\] _1855_ vssd1 vssd1 vccd1 vccd1 _1856_ sky130_fd_sc_hd__mux2_1
XANTENNA__2702__S _0788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4891__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2848__A0 _1225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2312__A2 net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4614__CLK clknet_leaf_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3500__A1 _1576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4940_ clknet_leaf_7_wb_clk_i _0550_ vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__dfxtp_2
XANTENNA__3264__A0 _1490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4764__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2583__A _0778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4274__S _2111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4871_ clknet_leaf_23_wb_clk_i _0485_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[87\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_60_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3822_ _1258_ _1337_ vssd1 vssd1 vccd1 vccd1 _1811_ sky130_fd_sc_hd__nor2_2
XFILLER_21_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3753_ tms1x00.RAM\[75\]\[3\] _1676_ _1767_ vssd1 vssd1 vccd1 vccd1 _1771_ sky130_fd_sc_hd__mux2_1
X_2704_ tms1x00.RAM\[64\]\[2\] tms1x00.RAM\[65\]\[2\] tms1x00.RAM\[66\]\[2\] tms1x00.RAM\[67\]\[2\]
+ _0840_ _0813_ vssd1 vssd1 vccd1 vccd1 _1095_ sky130_fd_sc_hd__mux4_1
X_3684_ _1703_ tms1x00.RAM\[64\]\[0\] _1732_ vssd1 vssd1 vccd1 vccd1 _1733_ sky130_fd_sc_hd__mux2_1
XFILLER_9_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4303__A _1250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2635_ _1018_ _1020_ _1024_ _1026_ _0804_ vssd1 vssd1 vccd1 vccd1 _1027_ sky130_fd_sc_hd__a221o_1
XANTENNA__3319__A1 _1461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2566_ _0951_ _0954_ _0957_ _0948_ _0942_ vssd1 vssd1 vccd1 vccd1 _0958_ sky130_fd_sc_hd__o221a_1
X_4305_ _2132_ vssd1 vssd1 vccd1 vccd1 _0616_ sky130_fd_sc_hd__clkbuf_1
X_2497_ _0798_ _0887_ _0889_ _0775_ vssd1 vssd1 vccd1 vccd1 _0890_ sky130_fd_sc_hd__o211a_1
XFILLER_68_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4236_ tms1x00.N\[2\] _2007_ vssd1 vssd1 vccd1 vccd1 _2094_ sky130_fd_sc_hd__or2_1
XFILLER_74_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4167_ tms1x00.PC\[1\] _2025_ vssd1 vssd1 vccd1 vccd1 _2038_ sky130_fd_sc_hd__nand2_1
XFILLER_56_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3118_ tms1x00.RAM\[10\]\[1\] _1328_ _1404_ vssd1 vssd1 vccd1 vccd1 _1406_ sky130_fd_sc_hd__mux2_1
XFILLER_82_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4098_ _1984_ vssd1 vssd1 vccd1 vccd1 _0557_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__3589__A _1261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3049_ _1364_ tms1x00.RAM\[96\]\[1\] _1362_ vssd1 vssd1 vccd1 vccd1 _1365_ sky130_fd_sc_hd__mux2_1
XFILLER_43_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4637__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2668__A _0819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4787__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4123__A _0738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2757__C1 _0775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2420_ _0812_ vssd1 vssd1 vccd1 vccd1 _0813_ sky130_fd_sc_hd__buf_6
XANTENNA__2509__C1 _0040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2351_ net148 _0721_ _0745_ vssd1 vssd1 vccd1 vccd1 _0746_ sky130_fd_sc_hd__a21o_2
X_2282_ net86 _0702_ _0703_ wbs_o_buff\[17\] vssd1 vssd1 vccd1 vccd1 _0011_ sky130_fd_sc_hd__a22o_1
X_4021_ _0732_ _0753_ _1928_ vssd1 vssd1 vccd1 vccd1 _1930_ sky130_fd_sc_hd__or3_1
XFILLER_38_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2288__A1 net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4029__A2 _0763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4923_ clknet_leaf_13_wb_clk_i _0533_ vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__dfxtp_2
XFILLER_33_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4854_ clknet_leaf_17_wb_clk_i _0468_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[81\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2460__B2 _0786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3805_ _1703_ tms1x00.RAM\[77\]\[0\] _1801_ vssd1 vssd1 vccd1 vccd1 _1802_ sky130_fd_sc_hd__mux2_1
X_4785_ clknet_leaf_24_wb_clk_i _0399_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[72\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2252__S net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3736_ _1761_ vssd1 vssd1 vccd1 vccd1 _0418_ sky130_fd_sc_hd__clkbuf_1
X_3667_ _1723_ vssd1 vssd1 vccd1 vccd1 _0387_ sky130_fd_sc_hd__clkbuf_1
X_2618_ tms1x00.RAM\[40\]\[1\] tms1x00.RAM\[41\]\[1\] tms1x00.RAM\[42\]\[1\] tms1x00.RAM\[43\]\[1\]
+ _0808_ _0780_ vssd1 vssd1 vccd1 vccd1 _1010_ sky130_fd_sc_hd__mux4_1
X_3598_ _1284_ _1303_ vssd1 vssd1 vccd1 vccd1 _1683_ sky130_fd_sc_hd__nor2_2
X_2549_ _0937_ _0938_ _0939_ _0787_ _0940_ vssd1 vssd1 vccd1 vccd1 _0941_ sky130_fd_sc_hd__a221o_1
XFILLER_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4219_ _0732_ _2082_ _2063_ vssd1 vssd1 vccd1 vccd1 _2083_ sky130_fd_sc_hd__mux2_1
XFILLER_75_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2279__A1 net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2935__B _1283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2451__A1 _0798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3400__A0 _1488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_3_wb_clk_i_A clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_3_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2398__A _0780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input53_A wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2337__S _0726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2580__B _0971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4802__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4570_ clknet_leaf_31_wb_clk_i _0191_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[120\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_3521_ _1638_ vssd1 vssd1 vccd1 vccd1 _0326_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__2745__A2 _1132_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3692__A _1237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4952__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3452_ _1600_ vssd1 vssd1 vccd1 vccd1 _0295_ sky130_fd_sc_hd__clkbuf_1
X_3383_ _1558_ vssd1 vssd1 vccd1 vccd1 _0268_ sky130_fd_sc_hd__clkbuf_1
X_2403_ _0787_ _0790_ _0795_ vssd1 vssd1 vccd1 vccd1 _0796_ sky130_fd_sc_hd__a21o_1
XFILLER_69_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2334_ _0734_ vssd1 vssd1 vccd1 vccd1 _0045_ sky130_fd_sc_hd__clkbuf_1
XFILLER_69_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2265_ net72 _0698_ _0700_ wbs_o_buff\[3\] vssd1 vssd1 vccd1 vccd1 _0028_ sky130_fd_sc_hd__a22o_1
X_4004_ _0732_ _0730_ _0752_ _1915_ vssd1 vssd1 vccd1 vccd1 _1917_ sky130_fd_sc_hd__or4b_1
X_2196_ net43 wbs_o_buff\[7\] _0657_ vssd1 vssd1 vccd1 vccd1 _0665_ sky130_fd_sc_hd__mux2_1
XFILLER_38_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2681__B2 _0807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4906_ clknet_leaf_7_wb_clk_i _0520_ vssd1 vssd1 vccd1 vccd1 tms1x00.ins_in\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3630__A0 _1590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4837_ clknet_leaf_23_wb_clk_i _0451_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[85\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4186__A1 tms1x00.PC\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4768_ clknet_leaf_12_wb_clk_i _0382_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[60\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_4699_ clknet_leaf_3_wb_clk_i _0313_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[50\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_3719_ _1317_ _1344_ vssd1 vssd1 vccd1 vccd1 _1752_ sky130_fd_sc_hd__nor2_2
XFILLER_76_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3777__A _1258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4825__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3621__A0 _1590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4975__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2188__A0 net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3688__A0 _1708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3017__A _1344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3451__S _1599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2856__A _1237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3860__A0 _1823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2663__A1 _0953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2952_ _1301_ vssd1 vssd1 vccd1 vccd1 _0094_ sky130_fd_sc_hd__clkbuf_1
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4168__A1 tms1x00.ins_in\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2883_ tms1x00.ram_addr_buff\[1\] _1259_ tms1x00.ram_addr_buff\[0\] vssd1 vssd1 vccd1
+ vccd1 _1260_ sky130_fd_sc_hd__or3b_1
XFILLER_30_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4622_ clknet_leaf_5_wb_clk_i _0243_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[32\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_4553_ clknet_leaf_30_wb_clk_i _0174_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[105\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_3504_ _1284_ _1345_ vssd1 vssd1 vccd1 vccd1 _1629_ sky130_fd_sc_hd__or2_2
X_4484_ clknet_leaf_30_wb_clk_i _0105_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[102\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_3435_ _1129_ vssd1 vssd1 vccd1 vccd1 _1590_ sky130_fd_sc_hd__buf_2
XANTENNA__4030__B _0752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3679__A0 _1708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3366_ tms1x00.RAM\[37\]\[2\] _1461_ _1546_ vssd1 vssd1 vccd1 vccd1 _1549_ sky130_fd_sc_hd__mux2_1
X_2317_ tms1x00.wb_step tms1x00.wb_step_state vssd1 vssd1 vccd1 vccd1 _0721_ sky130_fd_sc_hd__xnor2_2
XFILLER_58_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3297_ _1485_ tms1x00.RAM\[28\]\[0\] _1509_ vssd1 vssd1 vccd1 vccd1 _1510_ sky130_fd_sc_hd__mux2_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5105_ net47 vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__clkbuf_2
X_2248_ net2 K_override\[0\] net148 vssd1 vssd1 vccd1 vccd1 _0692_ sky130_fd_sc_hd__mux2_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5036_ clknet_leaf_2_wb_clk_i _0646_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[9\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_66_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4848__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3851__A0 _1823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2179_ net67 net58 vssd1 vssd1 vccd1 vccd1 _0656_ sky130_fd_sc_hd__and2_1
XFILLER_25_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4998__CLK clknet_leaf_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2590__B1 _0040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput89 net89 vssd1 vssd1 vccd1 vccd1 io_out[30] sky130_fd_sc_hd__buf_2
Xoutput78 net78 vssd1 vssd1 vccd1 vccd1 io_out[19] sky130_fd_sc_hd__buf_2
XFILLER_1_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input16_A ram_val[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3842__A0 _1823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5003__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4131__A _0858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output84_A net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3220_ _1317_ _1430_ vssd1 vssd1 vccd1 vccd1 _1465_ sky130_fd_sc_hd__nor2_2
XFILLER_79_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3151_ _1424_ vssd1 vssd1 vccd1 vccd1 _0170_ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3082_ _1384_ vssd1 vssd1 vccd1 vccd1 _0141_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2545__B_N _0924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3833__A0 _1816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3984_ tms1x00.ins_in\[4\] _0724_ _1903_ _1901_ vssd1 vssd1 vccd1 vccd1 _0524_ sky130_fd_sc_hd__o211a_1
XFILLER_16_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2935_ _1251_ _1283_ vssd1 vssd1 vccd1 vccd1 _1292_ sky130_fd_sc_hd__or2_2
XFILLER_31_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2495__S0 _0777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2866_ tms1x00.RAM\[69\]\[3\] _1247_ _1241_ vssd1 vssd1 vccd1 vccd1 _1248_ sky130_fd_sc_hd__mux2_1
X_4605_ clknet_leaf_4_wb_clk_i _0226_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[25\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_2797_ _0927_ _1186_ vssd1 vssd1 vccd1 vccd1 _1187_ sky130_fd_sc_hd__and2_1
XANTENNA__4520__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4536_ clknet_leaf_30_wb_clk_i _0157_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[10\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_4467_ clknet_leaf_10_wb_clk_i _0088_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[49\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3880__A _1258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3418_ _1579_ vssd1 vssd1 vccd1 vccd1 _0282_ sky130_fd_sc_hd__clkbuf_1
X_4398_ clknet_leaf_35_wb_clk_i _0025_ vssd1 vssd1 vccd1 vccd1 wbs_o_buff\[2\] sky130_fd_sc_hd__dfxtp_1
X_3349_ _1539_ vssd1 vssd1 vccd1 vccd1 _0253_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4670__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input8_A oram_value[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2496__A _0828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3104__B _1396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5019_ clknet_leaf_21_wb_clk_i _0629_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[15\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__5026__CLK clknet_leaf_20_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2418__B_N _0789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4304__A1 _1323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2866__A1 _1247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4126__A _0738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2720_ tms1x00.RAM\[124\]\[2\] tms1x00.RAM\[125\]\[2\] tms1x00.RAM\[126\]\[2\] tms1x00.RAM\[127\]\[2\]
+ _0816_ _0977_ vssd1 vssd1 vccd1 vccd1 _1111_ sky130_fd_sc_hd__mux4_1
XANTENNA__4543__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2651_ tms1x00.RAM\[36\]\[2\] tms1x00.RAM\[37\]\[2\] tms1x00.RAM\[38\]\[2\] tms1x00.RAM\[39\]\[2\]
+ _0799_ _0800_ vssd1 vssd1 vccd1 vccd1 _1042_ sky130_fd_sc_hd__mux4_2
X_2582_ tms1x00.RAM\[112\]\[1\] tms1x00.RAM\[113\]\[1\] tms1x00.RAM\[114\]\[1\] tms1x00.RAM\[115\]\[1\]
+ _0955_ _0956_ vssd1 vssd1 vccd1 vccd1 _0974_ sky130_fd_sc_hd__mux4_2
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4321_ _1267_ _1375_ vssd1 vssd1 vccd1 vccd1 _2141_ sky130_fd_sc_hd__or2_2
XANTENNA__4693__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4252_ tms1x00.RAM\[119\]\[1\] _1327_ _2101_ vssd1 vssd1 vccd1 vccd1 _2103_ sky130_fd_sc_hd__mux2_1
XFILLER_68_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3203_ tms1x00.RAM\[120\]\[2\] _1331_ _1451_ vssd1 vssd1 vccd1 vccd1 _1454_ sky130_fd_sc_hd__mux2_1
XFILLER_79_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4183_ tms1x00.PC\[4\] _1908_ vssd1 vssd1 vccd1 vccd1 _2052_ sky130_fd_sc_hd__or2_1
XANTENNA__2857__A1 _1235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3134_ _0914_ _1286_ vssd1 vssd1 vccd1 vccd1 _1415_ sky130_fd_sc_hd__nor2_2
XFILLER_82_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3065_ _1374_ vssd1 vssd1 vccd1 vccd1 _0134_ sky130_fd_sc_hd__clkbuf_1
XFILLER_82_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2704__S1 _0813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3967_ _1892_ vssd1 vssd1 vccd1 vccd1 _0518_ sky130_fd_sc_hd__clkbuf_1
X_2918_ K_override\[2\] net60 _0715_ vssd1 vssd1 vccd1 vccd1 _1281_ sky130_fd_sc_hd__mux2_1
XANTENNA__2793__B1 _0940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3898_ _1257_ _1396_ vssd1 vssd1 vccd1 vccd1 _1855_ sky130_fd_sc_hd__or2_2
X_2849_ _1234_ vssd1 vssd1 vccd1 vccd1 _0058_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4519_ clknet_leaf_15_wb_clk_i _0140_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[113\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3814__S _1806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3115__A _1344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4566__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2784__B1 _0804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4909__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2698__S0 _0931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4870_ clknet_leaf_19_wb_clk_i _0484_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[87\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4213__A0 tms1x00.Y\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3821_ _1810_ vssd1 vssd1 vccd1 vccd1 _0454_ sky130_fd_sc_hd__clkbuf_1
XFILLER_20_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2775__B1 _0927_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3752_ _1770_ vssd1 vssd1 vccd1 vccd1 _0425_ sky130_fd_sc_hd__clkbuf_1
X_3683_ _1236_ _1345_ vssd1 vssd1 vccd1 vccd1 _1732_ sky130_fd_sc_hd__or2_2
X_2703_ _0786_ _1093_ _0794_ vssd1 vssd1 vccd1 vccd1 _1094_ sky130_fd_sc_hd__a21o_1
XANTENNA__4303__B _1337_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2634_ _0783_ _1025_ _0774_ vssd1 vssd1 vccd1 vccd1 _1026_ sky130_fd_sc_hd__o21a_1
X_2565_ tms1x00.RAM\[88\]\[1\] tms1x00.RAM\[89\]\[1\] tms1x00.RAM\[90\]\[1\] tms1x00.RAM\[91\]\[1\]
+ _0955_ _0956_ vssd1 vssd1 vccd1 vccd1 _0957_ sky130_fd_sc_hd__mux4_1
XANTENNA__2622__S0 _0808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4304_ tms1x00.RAM\[20\]\[0\] _1323_ _2131_ vssd1 vssd1 vccd1 vccd1 _2132_ sky130_fd_sc_hd__mux2_1
X_2496_ _0828_ _0888_ vssd1 vssd1 vccd1 vccd1 _0889_ sky130_fd_sc_hd__or2_1
XANTENNA__4439__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4235_ _2093_ vssd1 vssd1 vccd1 vccd1 _0585_ sky130_fd_sc_hd__clkbuf_1
X_4166_ _0760_ _2036_ _2037_ _1966_ vssd1 vssd1 vccd1 vccd1 _0572_ sky130_fd_sc_hd__o211a_1
XFILLER_67_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3117_ _1405_ vssd1 vssd1 vccd1 vccd1 _0155_ sky130_fd_sc_hd__clkbuf_1
X_4097_ tms1x00.SR\[4\] tms1x00.PC\[4\] _1979_ vssd1 vssd1 vccd1 vccd1 _1984_ sky130_fd_sc_hd__mux2_1
XFILLER_56_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3589__B _1284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4589__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3048_ _1034_ vssd1 vssd1 vccd1 vccd1 _1364_ sky130_fd_sc_hd__clkbuf_4
XFILLER_70_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2463__C1 _0804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4999_ clknet_leaf_1_wb_clk_i _0609_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[21\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2613__S0 _0931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2668__B _1058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4375__S _2006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_17_wb_clk_i clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_6_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2859__A _1034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2350_ net76 net75 net74 vssd1 vssd1 vccd1 vccd1 _0745_ sky130_fd_sc_hd__nand3b_1
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2281_ net85 _0702_ _0703_ wbs_o_buff\[16\] vssd1 vssd1 vccd1 vccd1 _0010_ sky130_fd_sc_hd__a22o_1
X_4020_ _1928_ _0755_ _0764_ vssd1 vssd1 vccd1 vccd1 _1929_ sky130_fd_sc_hd__and3b_1
XANTENNA__4731__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2288__A2 _0697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2693__C1 _0944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4922_ clknet_leaf_13_wb_clk_i _0532_ vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__dfxtp_2
XANTENNA__4881__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4853_ clknet_leaf_17_wb_clk_i _0467_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[81\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3804_ _0917_ _1236_ vssd1 vssd1 vccd1 vccd1 _1801_ sky130_fd_sc_hd__or2_2
X_4784_ clknet_leaf_18_wb_clk_i _0398_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[64\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2533__S _0924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3735_ tms1x00.RAM\[68\]\[3\] _1676_ _1757_ vssd1 vssd1 vccd1 vccd1 _1761_ sky130_fd_sc_hd__mux2_1
X_3666_ _1703_ tms1x00.RAM\[66\]\[0\] _1722_ vssd1 vssd1 vccd1 vccd1 _1723_ sky130_fd_sc_hd__mux2_1
X_2617_ _0953_ _1008_ vssd1 vssd1 vccd1 vccd1 _1009_ sky130_fd_sc_hd__nor2_1
X_3597_ _1682_ vssd1 vssd1 vccd1 vccd1 _0358_ sky130_fd_sc_hd__clkbuf_1
X_2548_ _0819_ vssd1 vssd1 vccd1 vccd1 _0940_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__2920__A0 K_override\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4218_ _2080_ _2081_ vssd1 vssd1 vccd1 vccd1 _2082_ sky130_fd_sc_hd__xnor2_1
X_2479_ _0789_ tms1x00.RAM\[14\]\[0\] _0813_ vssd1 vssd1 vccd1 vccd1 _0872_ sky130_fd_sc_hd__o21a_1
XANTENNA__2629__B_N _0873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4149_ _2011_ _2022_ vssd1 vssd1 vccd1 vccd1 _2023_ sky130_fd_sc_hd__or2_1
XFILLER_56_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2451__A2 _0841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4604__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4754__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input46_A wb_rst_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2675__C1 _0942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2427__C1 _0819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4134__A _0701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3520_ _1592_ tms1x00.RAM\[47\]\[3\] _1634_ vssd1 vssd1 vccd1 vccd1 _1638_ sky130_fd_sc_hd__mux2_1
XANTENNA__2825__S0 _0923_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3692__B _1303_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3451_ _1585_ tms1x00.RAM\[45\]\[0\] _1599_ vssd1 vssd1 vccd1 vccd1 _1600_ sky130_fd_sc_hd__mux2_1
XFILLER_69_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3382_ _1488_ tms1x00.RAM\[35\]\[1\] _1556_ vssd1 vssd1 vccd1 vccd1 _1558_ sky130_fd_sc_hd__mux2_1
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2402_ _0791_ _0792_ _0794_ vssd1 vssd1 vccd1 vccd1 _0795_ sky130_fd_sc_hd__a21o_1
XFILLER_69_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2902__A0 _1225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2333_ _0733_ tms1x00.ram_addr_buff\[3\] _0726_ vssd1 vssd1 vccd1 vccd1 _0734_ sky130_fd_sc_hd__mux2_1
X_2264_ net71 _0698_ _0700_ wbs_o_buff\[2\] vssd1 vssd1 vccd1 vccd1 _0025_ sky130_fd_sc_hd__a22o_1
X_4003_ _0755_ _0739_ _0764_ _1915_ vssd1 vssd1 vccd1 vccd1 _1916_ sky130_fd_sc_hd__and4_1
XFILLER_37_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2195_ _0664_ vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__clkbuf_1
XFILLER_53_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4905_ clknet_leaf_8_wb_clk_i _0519_ vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__dfxtp_2
XANTENNA__4627__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3630__A1 tms1x00.RAM\[62\]\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4836_ clknet_leaf_18_wb_clk_i _0450_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[77\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4767_ clknet_leaf_20_wb_clk_i _0381_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[60\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_4698_ clknet_leaf_3_wb_clk_i _0312_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[50\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_3718_ _1751_ vssd1 vssd1 vccd1 vccd1 _0410_ sky130_fd_sc_hd__clkbuf_1
X_3649_ _1713_ vssd1 vssd1 vccd1 vccd1 _0379_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__3697__A1 _1674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2657__C1 _0953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3777__B _1345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3621__A1 tms1x00.RAM\[63\]\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2202__A net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3017__B _1345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2856__B _1240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2951_ _1225_ tms1x00.RAM\[19\]\[3\] _1297_ vssd1 vssd1 vccd1 vccd1 _1301_ sky130_fd_sc_hd__mux2_1
XANTENNA__3612__A1 _1674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_32_wb_clk_i clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_32_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2882_ tms1x00.ram_addr_buff\[2\] _0915_ tms1x00.ram_addr_buff\[3\] vssd1 vssd1 vccd1
+ vccd1 _1259_ sky130_fd_sc_hd__or3b_1
X_4621_ clknet_leaf_4_wb_clk_i _0242_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[26\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4552_ clknet_leaf_31_wb_clk_i _0173_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[105\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_3503_ _1628_ vssd1 vssd1 vccd1 vccd1 _0318_ sky130_fd_sc_hd__clkbuf_1
X_4483_ clknet_leaf_30_wb_clk_i _0104_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[102\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3128__A0 _1364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3434_ _1589_ vssd1 vssd1 vccd1 vccd1 _0288_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__3208__A _1286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2351__A1 net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3365_ _1548_ vssd1 vssd1 vccd1 vccd1 _0260_ sky130_fd_sc_hd__clkbuf_1
X_2316_ _0719_ net75 vssd1 vssd1 vccd1 vccd1 _0720_ sky130_fd_sc_hd__nor2_2
X_3296_ _1249_ _1409_ vssd1 vssd1 vccd1 vccd1 _1509_ sky130_fd_sc_hd__or2_2
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5104_ net57 vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__clkbuf_2
XFILLER_73_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2247_ _0691_ vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__clkbuf_1
X_5035_ clknet_leaf_30_wb_clk_i _0645_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[9\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_66_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2782__A _0783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3603__A1 _1674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4159__A2 net75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4819_ clknet_leaf_23_wb_clk_i _0433_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[73\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2590__A1 _0920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput79 net79 vssd1 vssd1 vccd1 vccd1 io_out[20] sky130_fd_sc_hd__buf_2
XFILLER_0_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4095__A1 tms1x00.PC\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4383__S _2006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2692__A _0953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2631__S _0778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4131__B _0903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2581__A1 _0940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output77_A net77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2333__A1 tms1x00.ram_addr_buff\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3150_ tms1x00.RAM\[106\]\[3\] _1334_ _1420_ vssd1 vssd1 vccd1 vccd1 _1424_ sky130_fd_sc_hd__mux2_1
XANTENNA__4472__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3081_ _1366_ tms1x00.RAM\[113\]\[2\] _1381_ vssd1 vssd1 vccd1 vccd1 _1384_ sky130_fd_sc_hd__mux2_1
XFILLER_67_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3983_ net10 _1899_ vssd1 vssd1 vccd1 vccd1 _1903_ sky130_fd_sc_hd__or2_1
XFILLER_22_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2495__S1 _0779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2934_ _1291_ vssd1 vssd1 vccd1 vccd1 _0086_ sky130_fd_sc_hd__clkbuf_1
X_2865_ _1224_ vssd1 vssd1 vccd1 vccd1 _1247_ sky130_fd_sc_hd__buf_4
X_4604_ clknet_leaf_4_wb_clk_i _0225_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[25\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4535_ clknet_leaf_30_wb_clk_i _0156_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[10\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_2796_ tms1x00.RAM\[6\]\[3\] tms1x00.RAM\[7\]\[3\] _0788_ vssd1 vssd1 vccd1 vccd1
+ _1186_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_27_wb_clk_i_A clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_4466_ clknet_leaf_10_wb_clk_i _0087_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[49\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_3417_ tms1x00.RAM\[41\]\[3\] _1578_ _1572_ vssd1 vssd1 vccd1 vccd1 _1579_ sky130_fd_sc_hd__mux2_1
XANTENNA__4815__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4397_ clknet_leaf_35_wb_clk_i _0014_ vssd1 vssd1 vccd1 vccd1 wbs_o_buff\[1\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__3880__B _1303_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3348_ _1490_ tms1x00.RAM\[30\]\[2\] _1536_ vssd1 vssd1 vccd1 vccd1 _1539_ sky130_fd_sc_hd__mux2_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3279_ tms1x00.RAM\[25\]\[0\] _1456_ _1499_ vssd1 vssd1 vccd1 vccd1 _1500_ sky130_fd_sc_hd__mux2_1
XFILLER_27_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4965__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5018_ clknet_leaf_21_wb_clk_i _0628_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[15\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2627__A2 tms1x00.RAM\[62\]\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2716__S _0789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output115_A net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2650_ tms1x00.RAM\[32\]\[2\] tms1x00.RAM\[33\]\[2\] tms1x00.RAM\[34\]\[2\] tms1x00.RAM\[35\]\[2\]
+ _0955_ _0956_ vssd1 vssd1 vccd1 vccd1 _1041_ sky130_fd_sc_hd__mux4_2
XANTENNA__3457__S _1599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3981__A net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2581_ _0940_ _0970_ _0972_ _0806_ vssd1 vssd1 vccd1 vccd1 _0973_ sky130_fd_sc_hd__o211a_1
X_4320_ _2140_ vssd1 vssd1 vccd1 vccd1 _0623_ sky130_fd_sc_hd__clkbuf_1
XFILLER_4_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4251_ _2102_ vssd1 vssd1 vccd1 vccd1 _0592_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3202_ _1453_ vssd1 vssd1 vccd1 vccd1 _0192_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4988__CLK clknet_leaf_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4182_ _2048_ _2050_ vssd1 vssd1 vccd1 vccd1 _2051_ sky130_fd_sc_hd__xor2_1
X_3133_ _1414_ vssd1 vssd1 vccd1 vccd1 _0162_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3064_ _1368_ tms1x00.RAM\[95\]\[3\] _1370_ vssd1 vssd1 vccd1 vccd1 _1374_ sky130_fd_sc_hd__mux2_1
XFILLER_36_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3966_ tms1x00.wb_step _0766_ vssd1 vssd1 vccd1 vccd1 _1892_ sky130_fd_sc_hd__and2_1
X_2917_ _1280_ vssd1 vssd1 vccd1 vccd1 _0080_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4075__A_N _0742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2793__A1 _0787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3897_ _1854_ vssd1 vssd1 vccd1 vccd1 _0486_ sky130_fd_sc_hd__clkbuf_1
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2848_ _1225_ tms1x00.RAM\[99\]\[3\] _1230_ vssd1 vssd1 vccd1 vccd1 _1234_ sky130_fd_sc_hd__mux2_1
XANTENNA__3742__A0 _1708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2779_ _0921_ _1168_ vssd1 vssd1 vccd1 vccd1 _1169_ sky130_fd_sc_hd__or2_1
XFILLER_3_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4518_ clknet_leaf_15_wb_clk_i _0139_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[113\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_4449_ clknet_leaf_22_wb_clk_i _0070_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[89\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_59_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3115__B _1403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2784__A1 _0944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2210__A _0672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2698__S1 _0932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2472__B1 _0828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3820_ tms1x00.RAM\[85\]\[3\] _1779_ _1806_ vssd1 vssd1 vccd1 vccd1 _1810_ sky130_fd_sc_hd__mux2_1
XFILLER_60_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2224__A0 net26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3751_ tms1x00.RAM\[75\]\[2\] _1674_ _1767_ vssd1 vssd1 vccd1 vccd1 _1770_ sky130_fd_sc_hd__mux2_1
XANTENNA__4660__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2775__A1 _0955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2702_ tms1x00.RAM\[68\]\[2\] tms1x00.RAM\[69\]\[2\] _0788_ vssd1 vssd1 vccd1 vccd1
+ _1093_ sky130_fd_sc_hd__mux2_1
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3682_ _1731_ vssd1 vssd1 vccd1 vccd1 _0394_ sky130_fd_sc_hd__clkbuf_1
X_2633_ tms1x00.RAM\[48\]\[1\] tms1x00.RAM\[49\]\[1\] tms1x00.RAM\[50\]\[1\] tms1x00.RAM\[51\]\[1\]
+ _0788_ _0780_ vssd1 vssd1 vccd1 vccd1 _1025_ sky130_fd_sc_hd__mux4_1
X_2564_ _0800_ vssd1 vssd1 vccd1 vccd1 _0956_ sky130_fd_sc_hd__buf_6
XFILLER_5_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2622__S1 _0831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4303_ _1250_ _1337_ vssd1 vssd1 vccd1 vccd1 _2131_ sky130_fd_sc_hd__nor2_2
XFILLER_59_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2495_ tms1x00.RAM\[36\]\[0\] tms1x00.RAM\[37\]\[0\] tms1x00.RAM\[38\]\[0\] tms1x00.RAM\[39\]\[0\]
+ _0777_ _0779_ vssd1 vssd1 vccd1 vccd1 _0888_ sky130_fd_sc_hd__mux4_1
X_4234_ tms1x00.N\[1\] _2007_ vssd1 vssd1 vccd1 vccd1 _2093_ sky130_fd_sc_hd__or2_1
X_4165_ tms1x00.PC\[1\] _1908_ vssd1 vssd1 vccd1 vccd1 _2037_ sky130_fd_sc_hd__or2_1
XFILLER_56_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3116_ tms1x00.RAM\[10\]\[0\] _1324_ _1404_ vssd1 vssd1 vccd1 vccd1 _1405_ sky130_fd_sc_hd__mux2_1
X_4096_ _1983_ vssd1 vssd1 vccd1 vccd1 _0556_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3047_ _1363_ vssd1 vssd1 vccd1 vccd1 _0127_ sky130_fd_sc_hd__clkbuf_1
XFILLER_24_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4998_ clknet_leaf_0_wb_clk_i _0608_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[21\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_3949_ _1883_ vssd1 vssd1 vccd1 vccd1 _0509_ sky130_fd_sc_hd__clkbuf_1
XFILLER_23_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3825__S _1811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2613__S1 _0956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4683__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3954__A0 tms1x00.Y\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5039__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2757__B2 _0807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2509__A1 _0039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2280_ net84 _0702_ _0703_ wbs_o_buff\[15\] vssd1 vssd1 vccd1 vccd1 _0009_ sky130_fd_sc_hd__a22o_1
XFILLER_77_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4921_ clknet_leaf_9_wb_clk_i _0531_ vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__dfxtp_2
XFILLER_52_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4852_ clknet_leaf_16_wb_clk_i _0466_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[82\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_3803_ _1800_ vssd1 vssd1 vccd1 vccd1 _0446_ sky130_fd_sc_hd__clkbuf_1
XFILLER_20_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4783_ clknet_leaf_18_wb_clk_i _0397_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[64\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_3734_ _1760_ vssd1 vssd1 vccd1 vccd1 _0417_ sky130_fd_sc_hd__clkbuf_1
X_3665_ _1237_ _1273_ vssd1 vssd1 vccd1 vccd1 _1722_ sky130_fd_sc_hd__or2_2
XANTENNA__4406__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2616_ tms1x00.RAM\[44\]\[1\] tms1x00.RAM\[45\]\[1\] tms1x00.RAM\[46\]\[1\] tms1x00.RAM\[47\]\[1\]
+ _0799_ _0800_ vssd1 vssd1 vccd1 vccd1 _1008_ sky130_fd_sc_hd__mux4_1
XANTENNA__4330__A _1267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3596_ tms1x00.RAM\[57\]\[3\] _1676_ _1678_ vssd1 vssd1 vccd1 vccd1 _1682_ sky130_fd_sc_hd__mux2_1
X_2547_ tms1x00.RAM\[76\]\[1\] tms1x00.RAM\[77\]\[1\] _0924_ vssd1 vssd1 vccd1 vccd1
+ _0939_ sky130_fd_sc_hd__mux2_1
XFILLER_69_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4556__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2478_ tms1x00.RAM\[15\]\[0\] _0789_ vssd1 vssd1 vccd1 vccd1 _0871_ sky130_fd_sc_hd__or2b_1
X_4217_ tms1x00.P\[3\] tms1x00.N\[3\] vssd1 vssd1 vccd1 vccd1 _2081_ sky130_fd_sc_hd__xor2_1
XFILLER_68_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4148_ _0743_ tms1x00.K_latch\[3\] _1956_ _2012_ _0732_ vssd1 vssd1 vccd1 vccd1 _2022_
+ sky130_fd_sc_hd__a32o_1
XFILLER_56_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2684__B1 _0812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4079_ _0760_ _1971_ vssd1 vssd1 vccd1 vccd1 _1972_ sky130_fd_sc_hd__nor2_1
XFILLER_55_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2436__B1 _0828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4189__B1 _0766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2372__C1 _0766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2695__A _0928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input39_A ram_val[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2675__B1 _1065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2770__S0 _0931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2978__A1 _1235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4134__B _2006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4429__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2825__S1 _0927_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4579__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3450_ _0917_ _1524_ vssd1 vssd1 vccd1 vccd1 _1599_ sky130_fd_sc_hd__or2_2
XANTENNA__3155__A1 _1328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3381_ _1557_ vssd1 vssd1 vccd1 vccd1 _0267_ sky130_fd_sc_hd__clkbuf_1
X_2401_ _0793_ vssd1 vssd1 vccd1 vccd1 _0794_ sky130_fd_sc_hd__clkbuf_4
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2332_ _0732_ vssd1 vssd1 vccd1 vccd1 _0733_ sky130_fd_sc_hd__buf_2
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4002_ tms1x00.Y\[1\] tms1x00.Y\[0\] vssd1 vssd1 vccd1 vccd1 _1915_ sky130_fd_sc_hd__and2b_1
X_2263_ net70 _0698_ _0700_ wbs_o_buff\[1\] vssd1 vssd1 vccd1 vccd1 _0014_ sky130_fd_sc_hd__a22o_1
XFILLER_65_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2194_ net42 wbs_o_buff\[6\] _0657_ vssd1 vssd1 vccd1 vccd1 _0664_ sky130_fd_sc_hd__mux2_1
XFILLER_80_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2969__A1 _1243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4904_ clknet_leaf_7_wb_clk_i _0518_ vssd1 vssd1 vccd1 vccd1 tms1x00.wb_step_state
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4835_ clknet_leaf_18_wb_clk_i _0449_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[77\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_4766_ clknet_leaf_21_wb_clk_i _0380_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[60\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4040__C1 _1931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3717_ tms1x00.RAM\[70\]\[3\] _1676_ _1747_ vssd1 vssd1 vccd1 vccd1 _1751_ sky130_fd_sc_hd__mux2_1
X_4697_ clknet_leaf_4_wb_clk_i _0311_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[50\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3648_ _1703_ tms1x00.RAM\[60\]\[0\] _1712_ vssd1 vssd1 vccd1 vccd1 _1713_ sky130_fd_sc_hd__mux2_1
XANTENNA__3146__A1 _1328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3579_ _1671_ vssd1 vssd1 vccd1 vccd1 _0351_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_2_wb_clk_i clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_29_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4721__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3137__A1 _1328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2896__A0 _0912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3314__A _1250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2743__S0 _0840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2950_ _1300_ vssd1 vssd1 vccd1 vccd1 _0093_ sky130_fd_sc_hd__clkbuf_1
XFILLER_15_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2881_ _1257_ vssd1 vssd1 vccd1 vccd1 _1258_ sky130_fd_sc_hd__buf_6
XFILLER_42_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2820__B1 _0791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4620_ clknet_leaf_4_wb_clk_i _0241_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[26\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_17_wb_clk_i_A clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_4551_ clknet_leaf_31_wb_clk_i _0172_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[105\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_3502_ tms1x00.RAM\[4\]\[3\] _1578_ _1624_ vssd1 vssd1 vccd1 vccd1 _1628_ sky130_fd_sc_hd__mux2_1
X_4482_ clknet_leaf_30_wb_clk_i _0103_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[102\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_3433_ _1588_ tms1x00.RAM\[3\]\[1\] _1586_ vssd1 vssd1 vccd1 vccd1 _1589_ sky130_fd_sc_hd__mux2_1
XANTENNA__3208__B _1344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5103_ net56 vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__clkbuf_2
X_3364_ tms1x00.RAM\[37\]\[1\] _1459_ _1546_ vssd1 vssd1 vccd1 vccd1 _1548_ sky130_fd_sc_hd__mux2_1
XFILLER_58_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2315_ net76 vssd1 vssd1 vccd1 vccd1 _0719_ sky130_fd_sc_hd__inv_2
XFILLER_57_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3295_ _1508_ vssd1 vssd1 vccd1 vccd1 _0230_ sky130_fd_sc_hd__clkbuf_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2246_ net38 wbs_o_buff\[31\] net49 vssd1 vssd1 vccd1 vccd1 _0691_ sky130_fd_sc_hd__mux2_1
X_5034_ clknet_leaf_30_wb_clk_i _0644_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[9\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_72_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2782__B _1171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3064__A0 _1368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4744__CLK clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4818_ clknet_leaf_23_wb_clk_i _0432_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[73\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4894__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4749_ clknet_leaf_22_wb_clk_i _0363_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[55\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput69 net69 vssd1 vssd1 vccd1 vccd1 io_out[10] sky130_fd_sc_hd__buf_2
XANTENNA__2878__A0 _1225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3134__A _0914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2725__S0 _0873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3055__A0 _1368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2566__C1 _0942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4617__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3044__A _0911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3080_ _1383_ vssd1 vssd1 vccd1 vccd1 _0140_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__3979__A _0718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4767__CLK clknet_leaf_20_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3046__A0 _1361_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3982_ _0743_ _0724_ _1902_ _1901_ vssd1 vssd1 vccd1 vccd1 _0523_ sky130_fd_sc_hd__o211a_1
XFILLER_50_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2933_ tms1x00.RAM\[59\]\[3\] _1247_ _1287_ vssd1 vssd1 vccd1 vccd1 _1291_ sky130_fd_sc_hd__mux2_1
XFILLER_22_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2864_ _1246_ vssd1 vssd1 vccd1 vccd1 _0061_ sky130_fd_sc_hd__clkbuf_1
X_2795_ _1181_ _1183_ _1184_ _0922_ _0942_ vssd1 vssd1 vccd1 vccd1 _1185_ sky130_fd_sc_hd__o221a_1
X_4603_ clknet_leaf_4_wb_clk_i _0224_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[25\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_891 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4534_ clknet_leaf_30_wb_clk_i _0155_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[10\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4465_ clknet_leaf_24_wb_clk_i _0086_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[59\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_4396_ clknet_leaf_35_wb_clk_i _0003_ vssd1 vssd1 vccd1 vccd1 wbs_o_buff\[0\] sky130_fd_sc_hd__dfxtp_1
X_3416_ _1224_ vssd1 vssd1 vccd1 vccd1 _1578_ sky130_fd_sc_hd__clkbuf_4
X_3347_ _1538_ vssd1 vssd1 vccd1 vccd1 _0252_ sky130_fd_sc_hd__clkbuf_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5017_ clknet_leaf_12_wb_clk_i _0627_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[127\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_3278_ _1250_ _1261_ vssd1 vssd1 vccd1 vccd1 _1499_ sky130_fd_sc_hd__nor2_2
XANTENNA__3889__A _1258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2627__A3 tms1x00.RAM\[63\]\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2229_ _0682_ vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__clkbuf_1
XFILLER_27_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4232__B _2007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3760__A1 _1775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input21_A ram_val[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3276__A0 _1492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output108_A net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2319__A_N _0701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2580_ _0807_ _0971_ vssd1 vssd1 vccd1 vccd1 _0972_ sky130_fd_sc_hd__or2_1
XANTENNA__3751__A1 _1674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4250_ tms1x00.RAM\[119\]\[0\] _1323_ _2101_ vssd1 vssd1 vccd1 vccd1 _2102_ sky130_fd_sc_hd__mux2_1
XFILLER_4_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4181_ tms1x00.PC\[4\] _2030_ _2049_ _1971_ vssd1 vssd1 vccd1 vccd1 _2050_ sky130_fd_sc_hd__o22a_1
X_3201_ tms1x00.RAM\[120\]\[1\] _1328_ _1451_ vssd1 vssd1 vccd1 vccd1 _1453_ sky130_fd_sc_hd__mux2_1
XFILLER_79_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3132_ _1368_ tms1x00.RAM\[108\]\[3\] _1410_ vssd1 vssd1 vccd1 vccd1 _1414_ sky130_fd_sc_hd__mux2_1
XANTENNA__2711__C1 _0802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3063_ _1373_ vssd1 vssd1 vccd1 vccd1 _0133_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__3267__A0 _1492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3965_ _1891_ vssd1 vssd1 vccd1 vccd1 _0517_ sky130_fd_sc_hd__clkbuf_1
X_3896_ tms1x00.RAM\[87\]\[3\] _1779_ _1850_ vssd1 vssd1 vccd1 vccd1 _1854_ sky130_fd_sc_hd__mux2_1
X_2916_ K_override\[1\] net66 _0715_ vssd1 vssd1 vccd1 vccd1 _1280_ sky130_fd_sc_hd__mux2_1
XFILLER_10_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4052__B _0730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2847_ _1233_ vssd1 vssd1 vccd1 vccd1 _0057_ sky130_fd_sc_hd__clkbuf_1
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2778_ tms1x00.RAM\[112\]\[3\] tms1x00.RAM\[113\]\[3\] tms1x00.RAM\[114\]\[3\] tms1x00.RAM\[115\]\[3\]
+ _0873_ _0977_ vssd1 vssd1 vccd1 vccd1 _1168_ sky130_fd_sc_hd__mux4_1
X_4517_ clknet_leaf_14_wb_clk_i _0138_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[114\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2788__A _0996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4448_ clknet_leaf_22_wb_clk_i _0069_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[89\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_59_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4379_ tms1x00.PC\[4\] net97 _2006_ vssd1 vssd1 vccd1 vccd1 _2173_ sky130_fd_sc_hd__mux2_1
XANTENNA__2300__B _0704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3258__A0 _1485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2769__C1 _0942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3430__A0 _1585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4462__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2784__A2 _1167_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4389__S _2006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3733__A1 _1674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2472__A1 _0786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4805__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3750_ _1769_ vssd1 vssd1 vccd1 vccd1 _0424_ sky130_fd_sc_hd__clkbuf_1
X_2701_ _0977_ _1091_ vssd1 vssd1 vccd1 vccd1 _1092_ sky130_fd_sc_hd__and2_1
X_3681_ _1710_ tms1x00.RAM\[65\]\[3\] _1727_ vssd1 vssd1 vccd1 vccd1 _1731_ sky130_fd_sc_hd__mux2_1
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4955__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2632_ _1021_ _1022_ _1023_ _0818_ _0794_ vssd1 vssd1 vccd1 vccd1 _1024_ sky130_fd_sc_hd__a221o_1
X_2563_ _0799_ vssd1 vssd1 vccd1 vccd1 _0955_ sky130_fd_sc_hd__buf_8
XANTENNA__3724__A1 _1674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4302_ _2130_ vssd1 vssd1 vccd1 vccd1 _0615_ sky130_fd_sc_hd__clkbuf_1
X_4233_ _2092_ vssd1 vssd1 vccd1 vccd1 _0584_ sky130_fd_sc_hd__clkbuf_1
X_2494_ tms1x00.RAM\[32\]\[0\] tms1x00.RAM\[33\]\[0\] tms1x00.RAM\[34\]\[0\] tms1x00.RAM\[35\]\[0\]
+ _0799_ _0800_ vssd1 vssd1 vccd1 vccd1 _0887_ sky130_fd_sc_hd__mux4_2
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4164_ _2025_ _2035_ vssd1 vssd1 vccd1 vccd1 _2036_ sky130_fd_sc_hd__xor2_1
XFILLER_68_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4095_ tms1x00.SR\[3\] tms1x00.PC\[3\] _1979_ vssd1 vssd1 vccd1 vccd1 _1983_ sky130_fd_sc_hd__mux2_1
XANTENNA__2547__S _0924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3115_ _1344_ _1403_ vssd1 vssd1 vccd1 vccd1 _1404_ sky130_fd_sc_hd__nor2_2
X_3046_ _1361_ tms1x00.RAM\[96\]\[0\] _1362_ vssd1 vssd1 vccd1 vccd1 _1363_ sky130_fd_sc_hd__mux2_1
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4063__A net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4997_ clknet_leaf_12_wb_clk_i _0607_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[29\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_3948_ tms1x00.RAM\[23\]\[2\] _1330_ _1880_ vssd1 vssd1 vccd1 vccd1 _1883_ sky130_fd_sc_hd__mux2_1
XFILLER_20_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3879_ _1844_ vssd1 vssd1 vccd1 vccd1 _0478_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3715__A1 _1674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3407__A _1261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4140__B2 tms1x00.Y\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4828__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2502__B_N _0778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4978__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2920__S _0715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3706__A1 _1674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_26_wb_clk_i clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__4065__A_N _0742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2693__A1 _0922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4920_ clknet_leaf_8_wb_clk_i tms1x00.K_in\[3\] vssd1 vssd1 vccd1 vccd1 tms1x00.K_latch\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3642__A0 _1708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4851_ clknet_leaf_16_wb_clk_i _0465_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[82\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_60_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3802_ _1710_ tms1x00.RAM\[78\]\[3\] _1796_ vssd1 vssd1 vccd1 vccd1 _1800_ sky130_fd_sc_hd__mux2_1
XFILLER_33_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4782_ clknet_leaf_18_wb_clk_i _0396_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[64\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_3733_ tms1x00.RAM\[68\]\[2\] _1674_ _1757_ vssd1 vssd1 vccd1 vccd1 _1760_ sky130_fd_sc_hd__mux2_1
X_3664_ _1721_ vssd1 vssd1 vccd1 vccd1 _0386_ sky130_fd_sc_hd__clkbuf_1
X_2615_ _0998_ _1000_ _1004_ _1006_ _0920_ vssd1 vssd1 vccd1 vccd1 _1007_ sky130_fd_sc_hd__o221a_1
XANTENNA__4330__B _1343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3595_ _1681_ vssd1 vssd1 vccd1 vccd1 _0357_ sky130_fd_sc_hd__clkbuf_1
X_2546_ _0924_ tms1x00.RAM\[78\]\[1\] _0932_ vssd1 vssd1 vccd1 vccd1 _0938_ sky130_fd_sc_hd__o21a_1
X_2477_ _0807_ _0869_ vssd1 vssd1 vccd1 vccd1 _0870_ sky130_fd_sc_hd__or2_1
X_4216_ _2074_ _2076_ _2073_ vssd1 vssd1 vccd1 vccd1 _2080_ sky130_fd_sc_hd__o21ba_1
XFILLER_68_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4147_ _2009_ _1221_ vssd1 vssd1 vccd1 vccd1 _2021_ sky130_fd_sc_hd__and2b_1
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4058__A tms1x00.ins_in\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2684__A1 _0788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4078_ net74 _0720_ vssd1 vssd1 vccd1 vccd1 _1971_ sky130_fd_sc_hd__nand2_4
X_3029_ _1035_ tms1x00.RAM\[98\]\[1\] _1351_ vssd1 vssd1 vccd1 vccd1 _1353_ sky130_fd_sc_hd__mux2_1
XFILLER_37_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2436__A1 _0786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4189__A1 tms1x00.PC\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4240__B _0738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4500__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4650__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2675__B2 _0948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2770__S1 _0932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2427__B2 _0818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5006__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2216__A _0675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2400_ _0037_ vssd1 vssd1 vccd1 vccd1 _0793_ sky130_fd_sc_hd__inv_2
X_3380_ _1485_ tms1x00.RAM\[35\]\[0\] _1556_ vssd1 vssd1 vccd1 vccd1 _1557_ sky130_fd_sc_hd__mux2_1
X_2331_ tms1x00.Y\[3\] vssd1 vssd1 vccd1 vccd1 _0732_ sky130_fd_sc_hd__buf_2
XFILLER_69_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4104__A1 tms1x00.PA\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2262_ net69 _0698_ _0700_ wbs_o_buff\[0\] vssd1 vssd1 vccd1 vccd1 _0003_ sky130_fd_sc_hd__a22o_1
XFILLER_66_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4001_ net103 _1914_ vssd1 vssd1 vccd1 vccd1 _0530_ sky130_fd_sc_hd__nor2_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2193_ _0663_ vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__clkbuf_1
XFILLER_37_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4903_ clknet_leaf_10_wb_clk_i _0517_ vssd1 vssd1 vccd1 vccd1 tms1x00.ram_addr_buff\[6\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_52_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4834_ clknet_leaf_17_wb_clk_i _0448_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[77\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4765_ clknet_leaf_20_wb_clk_i _0379_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[60\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2560__S _0923_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3716_ _1750_ vssd1 vssd1 vccd1 vccd1 _0409_ sky130_fd_sc_hd__clkbuf_1
X_4696_ clknet_leaf_32_wb_clk_i _0310_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[42\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_3647_ _1283_ _1409_ vssd1 vssd1 vccd1 vccd1 _1712_ sky130_fd_sc_hd__or2_2
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_918 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3578_ tms1x00.RAM\[58\]\[0\] _1669_ _1670_ vssd1 vssd1 vccd1 vccd1 _1671_ sky130_fd_sc_hd__mux2_1
XANTENNA__4673__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2529_ _0797_ vssd1 vssd1 vccd1 vccd1 _0921_ sky130_fd_sc_hd__clkbuf_4
XFILLER_29_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3854__A0 _1816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2657__B2 _0818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5029__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input51_A wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3845__A0 _1816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3314__B _1403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2743__S1 _0813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2880_ tms1x00.ram_addr_buff\[5\] tms1x00.ram_addr_buff\[6\] tms1x00.ram_addr_buff\[4\]
+ vssd1 vssd1 vccd1 vccd1 _1257_ sky130_fd_sc_hd__nand3b_4
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4546__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2820__A1 _0931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4550_ clknet_leaf_31_wb_clk_i _0171_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[105\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4696__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3501_ _1627_ vssd1 vssd1 vccd1 vccd1 _0317_ sky130_fd_sc_hd__clkbuf_1
X_4481_ clknet_leaf_29_wb_clk_i _0102_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[103\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_3432_ _1034_ vssd1 vssd1 vccd1 vccd1 _1588_ sky130_fd_sc_hd__buf_2
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3363_ _1547_ vssd1 vssd1 vccd1 vccd1 _0259_ sky130_fd_sc_hd__clkbuf_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5102_ net55 vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__clkbuf_2
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3294_ tms1x00.RAM\[24\]\[3\] _1463_ _1504_ vssd1 vssd1 vccd1 vccd1 _1508_ sky130_fd_sc_hd__mux2_1
X_2314_ wb_rst_override net46 vssd1 vssd1 vccd1 vccd1 _0718_ sky130_fd_sc_hd__nor2_8
XANTENNA__3836__A0 _1819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5033_ clknet_leaf_21_wb_clk_i _0643_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[14\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_2245_ _0690_ vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__clkbuf_1
XFILLER_66_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_2_wb_clk_i_A clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_25_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2498__S0 _0777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4817_ clknet_leaf_24_wb_clk_i _0431_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[73\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4748_ clknet_leaf_26_wb_clk_i _0362_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[56\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_4679_ clknet_leaf_1_wb_clk_i _0293_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[38\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4419__CLK clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3134__B _1286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2725__S1 _0822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2661__S0 _0815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3325__A _1345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3294__A1 _1463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3981_ net9 _1899_ vssd1 vssd1 vccd1 vccd1 _1902_ sky130_fd_sc_hd__or2_1
XFILLER_51_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3995__A _0718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2932_ _1290_ vssd1 vssd1 vccd1 vccd1 _0085_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__2736__B_N _0747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2863_ tms1x00.RAM\[69\]\[2\] _1245_ _1241_ vssd1 vssd1 vccd1 vccd1 _1246_ sky130_fd_sc_hd__mux2_1
X_2794_ tms1x00.RAM\[24\]\[3\] tms1x00.RAM\[25\]\[3\] tms1x00.RAM\[26\]\[3\] tms1x00.RAM\[27\]\[3\]
+ _0924_ _0928_ vssd1 vssd1 vccd1 vccd1 _1184_ sky130_fd_sc_hd__mux4_2
X_4602_ clknet_leaf_4_wb_clk_i _0223_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[25\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4533_ clknet_leaf_14_wb_clk_i _0154_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[110\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_4464_ clknet_leaf_28_wb_clk_i _0085_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[59\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_4395_ clknet_leaf_34_wb_clk_i _0050_ vssd1 vssd1 vccd1 vccd1 chip_sel_override sky130_fd_sc_hd__dfxtp_1
X_3415_ _1577_ vssd1 vssd1 vccd1 vccd1 _0281_ sky130_fd_sc_hd__clkbuf_1
X_3346_ _1488_ tms1x00.RAM\[30\]\[1\] _1536_ vssd1 vssd1 vccd1 vccd1 _1538_ sky130_fd_sc_hd__mux2_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3809__A0 _1708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5016_ clknet_leaf_14_wb_clk_i _0626_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[127\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_3277_ _1498_ vssd1 vssd1 vccd1 vccd1 _0222_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4711__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3889__B _1310_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3285__A1 _1463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2228_ net28 wbs_o_buff\[22\] _0679_ vssd1 vssd1 vccd1 vccd1 _0682_ sky130_fd_sc_hd__mux2_1
XFILLER_26_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4066__A net70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2493__C1 _0802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4391__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input14_A ram_val[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2759__B_N _0778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3984__C1 _1901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output82_A net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4161__C1 _1966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4180_ _0748_ _1995_ _2027_ tms1x00.SR\[4\] vssd1 vssd1 vccd1 vccd1 _2049_ sky130_fd_sc_hd__o22a_1
XANTENNA__4734__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3200_ _1452_ vssd1 vssd1 vccd1 vccd1 _0191_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3131_ _1413_ vssd1 vssd1 vccd1 vccd1 _0161_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3062_ _1366_ tms1x00.RAM\[95\]\[2\] _1370_ vssd1 vssd1 vccd1 vccd1 _1373_ sky130_fd_sc_hd__mux2_1
XANTENNA__4884__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2475__C1 _0804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3964_ tms1x00.X\[1\] tms1x00.ram_addr_buff\[6\] _0725_ vssd1 vssd1 vccd1 vccd1 _1891_
+ sky130_fd_sc_hd__mux2_1
XFILLER_50_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3895_ _1853_ vssd1 vssd1 vccd1 vccd1 _0485_ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2915_ _1279_ vssd1 vssd1 vccd1 vccd1 _0079_ sky130_fd_sc_hd__clkbuf_1
X_2846_ _1130_ tms1x00.RAM\[99\]\[2\] _1230_ vssd1 vssd1 vccd1 vccd1 _1233_ sky130_fd_sc_hd__mux2_1
XANTENNA__4052__C _0763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2777_ _1164_ _1165_ _1166_ _0787_ _0996_ vssd1 vssd1 vccd1 vccd1 _1167_ sky130_fd_sc_hd__a221o_1
XANTENNA__2625__S0 _0823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4516_ clknet_leaf_15_wb_clk_i _0137_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[114\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2788__B _1177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4447_ clknet_leaf_21_wb_clk_i _0068_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[89\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_59_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4378_ _2172_ vssd1 vssd1 vccd1 vccd1 _0649_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_input6_A oram_value[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3329_ _1528_ vssd1 vssd1 vccd1 vccd1 _0244_ sky130_fd_sc_hd__clkbuf_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4607__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2616__S0 _0799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4757__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2918__S _0715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2700_ tms1x00.RAM\[70\]\[2\] tms1x00.RAM\[71\]\[2\] _0788_ vssd1 vssd1 vccd1 vccd1
+ _1091_ sky130_fd_sc_hd__mux2_1
X_3680_ _1730_ vssd1 vssd1 vccd1 vccd1 _0393_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__2607__S0 _0955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2631_ tms1x00.RAM\[52\]\[1\] tms1x00.RAM\[53\]\[1\] _0778_ vssd1 vssd1 vccd1 vccd1
+ _1023_ sky130_fd_sc_hd__mux2_1
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2562_ _0928_ _0952_ _0953_ vssd1 vssd1 vccd1 vccd1 _0954_ sky130_fd_sc_hd__a21o_1
X_4301_ _1823_ tms1x00.RAM\[16\]\[3\] _2126_ vssd1 vssd1 vccd1 vccd1 _2130_ sky130_fd_sc_hd__mux2_1
XFILLER_5_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4232_ tms1x00.N\[0\] _2007_ vssd1 vssd1 vccd1 vccd1 _2092_ sky130_fd_sc_hd__or2_1
X_2493_ _0819_ _0883_ _0885_ _0802_ vssd1 vssd1 vccd1 vccd1 _0886_ sky130_fd_sc_hd__o211a_1
XFILLER_68_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4163_ tms1x00.PC\[1\] _2030_ _2034_ _1971_ vssd1 vssd1 vccd1 vccd1 _2035_ sky130_fd_sc_hd__o22a_1
XANTENNA__3513__A _1267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4094_ _1982_ vssd1 vssd1 vccd1 vccd1 _0555_ sky130_fd_sc_hd__clkbuf_1
XFILLER_56_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3114_ _1402_ vssd1 vssd1 vccd1 vccd1 _1403_ sky130_fd_sc_hd__buf_6
XFILLER_82_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3045_ _0913_ _1345_ vssd1 vssd1 vccd1 vccd1 _1362_ sky130_fd_sc_hd__or2_2
XFILLER_36_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4996_ clknet_leaf_11_wb_clk_i _0606_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[29\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3947_ _1882_ vssd1 vssd1 vccd1 vccd1 _0508_ sky130_fd_sc_hd__clkbuf_1
X_3878_ tms1x00.RAM\[8\]\[3\] _1779_ _1840_ vssd1 vssd1 vccd1 vccd1 _1844_ sky130_fd_sc_hd__mux2_1
X_2829_ _0944_ _1212_ _1214_ _0920_ _1218_ vssd1 vssd1 vccd1 vccd1 _1219_ sky130_fd_sc_hd__a311o_1
XANTENNA__3407__B _1525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2687__C1 _0802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4238__B _2007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3167__A0 _1366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2914__A0 K_override\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3890__A1 _1772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2693__A2 _1081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4850_ clknet_leaf_17_wb_clk_i _0464_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[82\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3801_ _1799_ vssd1 vssd1 vccd1 vccd1 _0445_ sky130_fd_sc_hd__clkbuf_1
X_4781_ clknet_leaf_19_wb_clk_i _0395_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[64\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3732_ _1759_ vssd1 vssd1 vccd1 vccd1 _0416_ sky130_fd_sc_hd__clkbuf_1
X_3663_ _1710_ tms1x00.RAM\[67\]\[3\] _1717_ vssd1 vssd1 vccd1 vccd1 _1721_ sky130_fd_sc_hd__mux2_1
XFILLER_9_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2614_ _0948_ _1005_ _0942_ vssd1 vssd1 vccd1 vccd1 _1006_ sky130_fd_sc_hd__o21ai_1
X_3594_ tms1x00.RAM\[57\]\[2\] _1674_ _1678_ vssd1 vssd1 vccd1 vccd1 _1681_ sky130_fd_sc_hd__mux2_1
X_2545_ tms1x00.RAM\[79\]\[1\] _0924_ vssd1 vssd1 vccd1 vccd1 _0937_ sky130_fd_sc_hd__or2b_1
X_2476_ tms1x00.RAM\[8\]\[0\] tms1x00.RAM\[9\]\[0\] tms1x00.RAM\[10\]\[0\] tms1x00.RAM\[11\]\[0\]
+ _0808_ _0780_ vssd1 vssd1 vccd1 vccd1 _0869_ sky130_fd_sc_hd__mux4_1
XANTENNA__2558__S _0816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4215_ _2079_ vssd1 vssd1 vccd1 vccd1 _0579_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4339__A _1251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2669__C1 _0776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3330__A0 _1490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4146_ tms1x00.P\[2\] _2007_ _2018_ _2020_ vssd1 vssd1 vccd1 vccd1 _0569_ sky130_fd_sc_hd__o22a_1
XFILLER_55_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4452__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3881__A1 _1772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4077_ _1958_ _1969_ _1970_ _1966_ vssd1 vssd1 vccd1 vccd1 _0550_ sky130_fd_sc_hd__o211a_1
XFILLER_28_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3028_ _1352_ vssd1 vssd1 vccd1 vccd1 _0119_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4979_ clknet_leaf_8_wb_clk_i _0589_ vssd1 vssd1 vccd1 vccd1 tms1x00.A\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_50_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4249__A _1310_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2468__S _0783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3872__A1 _1772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2992__A _1327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2330_ _0731_ vssd1 vssd1 vccd1 vccd1 _0044_ sky130_fd_sc_hd__clkbuf_1
XFILLER_69_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2261_ _0699_ vssd1 vssd1 vccd1 vccd1 _0700_ sky130_fd_sc_hd__buf_2
XFILLER_66_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4000_ net76 _1909_ _0761_ vssd1 vssd1 vccd1 vccd1 _1914_ sky130_fd_sc_hd__a21oi_1
XFILLER_65_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2192_ net41 wbs_o_buff\[5\] _0657_ vssd1 vssd1 vccd1 vccd1 _0663_ sky130_fd_sc_hd__mux2_1
XANTENNA__3863__A1 _1772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4902_ clknet_leaf_10_wb_clk_i _0516_ vssd1 vssd1 vccd1 vccd1 tms1x00.ram_addr_buff\[5\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_52_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2407__A _0779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4833_ clknet_leaf_17_wb_clk_i _0447_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[77\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_4764_ clknet_leaf_12_wb_clk_i _0378_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[61\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3715_ tms1x00.RAM\[70\]\[2\] _1674_ _1747_ vssd1 vssd1 vccd1 vccd1 _1750_ sky130_fd_sc_hd__mux2_1
X_4695_ clknet_leaf_31_wb_clk_i _0309_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[42\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3238__A _1337_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3646_ _1711_ vssd1 vssd1 vccd1 vccd1 _0378_ sky130_fd_sc_hd__clkbuf_1
X_3577_ _1284_ _1403_ vssd1 vssd1 vccd1 vccd1 _1670_ sky130_fd_sc_hd__nor2_2
X_2528_ _0804_ vssd1 vssd1 vccd1 vccd1 _0920_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4069__A net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4968__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3303__A0 _1492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2459_ tms1x00.RAM\[116\]\[0\] tms1x00.RAM\[117\]\[0\] _0788_ vssd1 vssd1 vccd1 vccd1
+ _0852_ sky130_fd_sc_hd__mux2_1
XFILLER_29_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4129_ _2005_ vssd1 vssd1 vccd1 vccd1 _2006_ sky130_fd_sc_hd__buf_4
XFILLER_44_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3701__A _1237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2317__A tms1x00.wb_step vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4498__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2987__A _1323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input44_A ram_val[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4270__A1 _1327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2281__B1 _0703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3757__S _1773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3500_ tms1x00.RAM\[4\]\[2\] _1576_ _1624_ vssd1 vssd1 vccd1 vccd1 _1627_ sky130_fd_sc_hd__mux2_1
X_4480_ clknet_leaf_30_wb_clk_i _0101_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[103\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_3431_ _1587_ vssd1 vssd1 vccd1 vccd1 _0287_ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3362_ tms1x00.RAM\[37\]\[0\] _1456_ _1546_ vssd1 vssd1 vccd1 vccd1 _1547_ sky130_fd_sc_hd__mux2_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2313_ tms1x00.ram_addr_buff\[0\] vssd1 vssd1 vccd1 vccd1 _0717_ sky130_fd_sc_hd__clkbuf_4
X_5101_ net54 vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__clkbuf_2
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3293_ _1507_ vssd1 vssd1 vccd1 vccd1 _0229_ sky130_fd_sc_hd__clkbuf_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5032_ clknet_leaf_21_wb_clk_i _0642_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[14\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_2244_ net37 wbs_o_buff\[30\] net49 vssd1 vssd1 vccd1 vccd1 _0690_ sky130_fd_sc_hd__mux2_1
XFILLER_65_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_10_wb_clk_i clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_38_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2498__S1 _0779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4261__A1 _1327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4816_ clknet_leaf_23_wb_clk_i _0430_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[74\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_4747_ clknet_leaf_24_wb_clk_i _0361_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[56\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4640__CLK clknet_leaf_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4678_ clknet_leaf_1_wb_clk_i _0292_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[38\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_3629_ _1700_ vssd1 vssd1 vccd1 vccd1 _0372_ sky130_fd_sc_hd__clkbuf_1
XFILLER_1_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4790__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3827__A1 _1777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2746__S _0923_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4252__A1 _1327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2481__S _0873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2566__B2 _0948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2661__S1 _0812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3325__B _1525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3818__A1 _1777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2656__S _0923_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4513__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3980_ tms1x00.ins_in\[2\] _0724_ _1900_ _1901_ vssd1 vssd1 vccd1 vccd1 _0522_ sky130_fd_sc_hd__o211a_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2931_ tms1x00.RAM\[59\]\[2\] _1245_ _1287_ vssd1 vssd1 vccd1 vccd1 _1290_ sky130_fd_sc_hd__mux2_1
XANTENNA__2391__S _0783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4601_ clknet_leaf_12_wb_clk_i _0222_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[125\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_2862_ _1129_ vssd1 vssd1 vccd1 vccd1 _1245_ sky130_fd_sc_hd__buf_4
XFILLER_31_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2793_ _0787_ _1182_ _0940_ vssd1 vssd1 vccd1 vccd1 _1183_ sky130_fd_sc_hd__a21o_1
X_4532_ clknet_leaf_14_wb_clk_i _0153_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[110\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5019__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4463_ clknet_leaf_22_wb_clk_i _0084_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[59\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2420__A _0812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3414_ tms1x00.RAM\[41\]\[2\] _1576_ _1572_ vssd1 vssd1 vccd1 vccd1 _1577_ sky130_fd_sc_hd__mux2_1
X_4394_ clknet_leaf_34_wb_clk_i _0001_ vssd1 vssd1 vccd1 vccd1 wb_rst_override sky130_fd_sc_hd__dfxtp_1
X_3345_ _1537_ vssd1 vssd1 vccd1 vccd1 _0251_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__3950__S _1880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3276_ _1492_ tms1x00.RAM\[125\]\[3\] _1494_ vssd1 vssd1 vccd1 vccd1 _1498_ sky130_fd_sc_hd__mux2_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5015_ clknet_leaf_14_wb_clk_i _0625_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[127\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2227_ _0681_ vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__clkbuf_1
XFILLER_66_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4082__A tms1x00.ins_in\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3161__A _1375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4686__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2236__A0 net32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3984__B1 _1903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output75_A net75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3130_ _1366_ tms1x00.RAM\[108\]\[2\] _1410_ vssd1 vssd1 vccd1 vccd1 _1413_ sky130_fd_sc_hd__mux2_1
XANTENNA__2711__A1 _0921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3061_ _1372_ vssd1 vssd1 vccd1 vccd1 _0132_ sky130_fd_sc_hd__clkbuf_1
XFILLER_36_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3963_ _1890_ vssd1 vssd1 vccd1 vccd1 _0516_ sky130_fd_sc_hd__clkbuf_1
XFILLER_50_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3894_ tms1x00.RAM\[87\]\[2\] _1777_ _1850_ vssd1 vssd1 vccd1 vccd1 _1853_ sky130_fd_sc_hd__mux2_1
XANTENNA__2415__A _0777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2914_ K_override\[0\] net65 _0715_ vssd1 vssd1 vccd1 vccd1 _1279_ sky130_fd_sc_hd__mux2_1
X_2845_ _1232_ vssd1 vssd1 vccd1 vccd1 _0056_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4409__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4515_ clknet_leaf_14_wb_clk_i _0136_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[114\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_2776_ tms1x00.RAM\[116\]\[3\] tms1x00.RAM\[117\]\[3\] _0789_ vssd1 vssd1 vccd1 vccd1
+ _1166_ sky130_fd_sc_hd__mux2_1
XANTENNA__2625__S1 _0850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4446_ clknet_leaf_21_wb_clk_i _0067_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[89\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_4377_ tms1x00.PC\[3\] net96 _2006_ vssd1 vssd1 vccd1 vccd1 _2172_ sky130_fd_sc_hd__mux2_1
XANTENNA__2389__S0 _0778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3328_ _1488_ tms1x00.RAM\[32\]\[1\] _1526_ vssd1 vssd1 vccd1 vccd1 _1528_ sky130_fd_sc_hd__mux2_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3259_ _1487_ vssd1 vssd1 vccd1 vccd1 _0215_ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2309__B _0715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2769__A1 _0940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2616__S1 _0800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3194__A1 _1331_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output113_A net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_26_wb_clk_i_A clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_17_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2630_ _0840_ tms1x00.RAM\[54\]\[1\] _0780_ vssd1 vssd1 vccd1 vccd1 _1022_ sky130_fd_sc_hd__o21a_1
XANTENNA__2607__S1 _0956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3185__A1 _1331_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2561_ _0794_ vssd1 vssd1 vccd1 vccd1 _0953_ sky130_fd_sc_hd__buf_4
X_4300_ _2129_ vssd1 vssd1 vccd1 vccd1 _0614_ sky130_fd_sc_hd__clkbuf_1
X_2492_ _0797_ _0884_ vssd1 vssd1 vccd1 vccd1 _0885_ sky130_fd_sc_hd__or2_1
XANTENNA__4851__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4231_ tms1x00.X\[2\] _2088_ _2091_ _0766_ vssd1 vssd1 vccd1 vccd1 _0583_ sky130_fd_sc_hd__o211a_1
XFILLER_4_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4162_ _0743_ _1995_ _2027_ tms1x00.SR\[1\] vssd1 vssd1 vccd1 vccd1 _2034_ sky130_fd_sc_hd__o22a_1
XFILLER_68_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4093_ tms1x00.SR\[2\] tms1x00.PC\[2\] _1979_ vssd1 vssd1 vccd1 vccd1 _1982_ sky130_fd_sc_hd__mux2_1
XFILLER_56_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3113_ _1259_ tms1x00.ram_addr_buff\[0\] tms1x00.ram_addr_buff\[1\] vssd1 vssd1 vccd1
+ vccd1 _1402_ sky130_fd_sc_hd__or3b_1
XFILLER_67_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3044_ _0911_ vssd1 vssd1 vccd1 vccd1 _1361_ sky130_fd_sc_hd__buf_2
XFILLER_82_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4995_ clknet_leaf_12_wb_clk_i _0605_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[29\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3946_ tms1x00.RAM\[23\]\[1\] _1327_ _1880_ vssd1 vssd1 vccd1 vccd1 _1882_ sky130_fd_sc_hd__mux2_1
X_3877_ _1843_ vssd1 vssd1 vccd1 vccd1 _0477_ sky130_fd_sc_hd__clkbuf_1
X_2828_ _0940_ _1215_ _1217_ _0806_ vssd1 vssd1 vccd1 vccd1 _1218_ sky130_fd_sc_hd__o211a_1
XANTENNA__3176__A1 _1331_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2759_ tms1x00.RAM\[79\]\[3\] _0778_ vssd1 vssd1 vccd1 vccd1 _1149_ sky130_fd_sc_hd__or2b_1
XFILLER_3_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4429_ clknet_leaf_32_wb_clk_i valid vssd1 vssd1 vccd1 vccd1 feedback_delay sky130_fd_sc_hd__dfxtp_1
XFILLER_58_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2754__S _0826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3939__A0 tms1x00.RAM\[90\]\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4724__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2611__B1 _0996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4364__A0 _1247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3800_ _1708_ tms1x00.RAM\[78\]\[2\] _1796_ vssd1 vssd1 vccd1 vccd1 _1799_ sky130_fd_sc_hd__mux2_1
X_4780_ clknet_leaf_18_wb_clk_i _0394_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[65\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3731_ tms1x00.RAM\[68\]\[1\] _1672_ _1757_ vssd1 vssd1 vccd1 vccd1 _1759_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_35_wb_clk_i clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_35_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_3662_ _1720_ vssd1 vssd1 vccd1 vccd1 _0385_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4355__A0 _1247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2613_ tms1x00.RAM\[8\]\[1\] tms1x00.RAM\[9\]\[1\] tms1x00.RAM\[10\]\[1\] tms1x00.RAM\[11\]\[1\]
+ _0931_ _0956_ vssd1 vssd1 vccd1 vccd1 _1005_ sky130_fd_sc_hd__mux4_1
X_3593_ _1680_ vssd1 vssd1 vccd1 vccd1 _0356_ sky130_fd_sc_hd__clkbuf_1
X_2544_ tms1x00.RAM\[72\]\[1\] tms1x00.RAM\[73\]\[1\] tms1x00.RAM\[74\]\[1\] tms1x00.RAM\[75\]\[1\]
+ _0924_ _0928_ vssd1 vssd1 vccd1 vccd1 _0936_ sky130_fd_sc_hd__mux4_1
XFILLER_5_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2475_ _0776_ _0861_ _0867_ _0804_ vssd1 vssd1 vccd1 vccd1 _0868_ sky130_fd_sc_hd__a211o_1
X_4214_ _0766_ _2078_ vssd1 vssd1 vccd1 vccd1 _2079_ sky130_fd_sc_hd__and2_1
XANTENNA__4339__B _1343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4145_ _0730_ _2012_ _2019_ _2011_ vssd1 vssd1 vccd1 vccd1 _2020_ sky130_fd_sc_hd__a211o_1
XFILLER_55_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4076_ net73 _1960_ vssd1 vssd1 vccd1 vccd1 _1970_ sky130_fd_sc_hd__or2_1
XFILLER_55_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3027_ _0912_ tms1x00.RAM\[98\]\[0\] _1351_ vssd1 vssd1 vccd1 vccd1 _1352_ sky130_fd_sc_hd__mux2_1
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4747__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4978_ clknet_leaf_8_wb_clk_i _0588_ vssd1 vssd1 vccd1 vccd1 tms1x00.A\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_52_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4897__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3929_ _1872_ vssd1 vssd1 vccd1 vccd1 _0500_ sky130_fd_sc_hd__clkbuf_1
XFILLER_50_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4346__A0 _1247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4249__B _1430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3321__A1 _1463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4034__C1 _0766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4337__A0 _1247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2260_ net46 _0697_ vssd1 vssd1 vccd1 vccd1 _0699_ sky130_fd_sc_hd__nor2_4
XANTENNA__3312__A1 _1463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2191_ _0662_ vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__clkbuf_1
XFILLER_37_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4901_ clknet_leaf_9_wb_clk_i _0515_ vssd1 vssd1 vccd1 vccd1 tms1x00.ram_addr_buff\[4\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_45_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4832_ clknet_leaf_20_wb_clk_i _0446_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[78\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_60_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4763_ clknet_leaf_20_wb_clk_i _0377_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[61\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2423__A _0815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4694_ clknet_leaf_32_wb_clk_i _0308_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[42\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_3714_ _1749_ vssd1 vssd1 vccd1 vccd1 _0408_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4328__A0 _1823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3238__B _1430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3645_ _1710_ tms1x00.RAM\[61\]\[3\] _1704_ vssd1 vssd1 vccd1 vccd1 _1711_ sky130_fd_sc_hd__mux2_1
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3576_ _0911_ vssd1 vssd1 vccd1 vccd1 _1669_ sky130_fd_sc_hd__clkbuf_4
X_2527_ _0919_ vssd1 vssd1 vccd1 vccd1 _0051_ sky130_fd_sc_hd__clkbuf_1
X_2458_ _0808_ tms1x00.RAM\[118\]\[0\] _0850_ vssd1 vssd1 vccd1 vccd1 _0851_ sky130_fd_sc_hd__o21a_1
XFILLER_68_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2389_ tms1x00.RAM\[84\]\[0\] tms1x00.RAM\[85\]\[0\] tms1x00.RAM\[86\]\[0\] tms1x00.RAM\[87\]\[0\]
+ _0778_ _0780_ vssd1 vssd1 vccd1 vccd1 _0782_ sky130_fd_sc_hd__mux4_1
XFILLER_72_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4128_ _0738_ _0760_ _1912_ vssd1 vssd1 vccd1 vccd1 _2005_ sky130_fd_sc_hd__or3b_1
XFILLER_56_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4059_ _0743_ _0768_ tms1x00.ins_in\[1\] _1956_ vssd1 vssd1 vccd1 vccd1 _1957_ sky130_fd_sc_hd__and4_1
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3701__B _1310_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3429__A _1229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4319__A0 _1823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4912__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input37_A ram_val[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3058__A0 _1361_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2281__A1 net85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4442__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3430_ _1585_ tms1x00.RAM\[3\]\[0\] _1586_ vssd1 vssd1 vccd1 vccd1 _1587_ sky130_fd_sc_hd__mux2_1
X_3361_ _1240_ _1525_ vssd1 vssd1 vccd1 vccd1 _1546_ sky130_fd_sc_hd__nor2_2
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2312_ _0713_ net148 _0714_ _0716_ vssd1 vssd1 vccd1 vccd1 _0000_ sky130_fd_sc_hd__a31o_1
X_5100_ net53 vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__clkbuf_2
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3292_ tms1x00.RAM\[24\]\[2\] _1461_ _1504_ vssd1 vssd1 vccd1 vccd1 _1507_ sky130_fd_sc_hd__mux2_1
X_5031_ clknet_leaf_21_wb_clk_i _0641_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[14\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_78_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3297__A0 _1485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2243_ _0689_ vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__clkbuf_1
XFILLER_66_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3049__A0 _1364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3948__S _1880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2272__A1 net78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2272__B2 wbs_o_buff\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4815_ clknet_leaf_22_wb_clk_i _0429_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[74\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4746_ clknet_leaf_25_wb_clk_i _0360_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[56\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_4677_ clknet_leaf_1_wb_clk_i _0291_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[38\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_3628_ _1588_ tms1x00.RAM\[62\]\[1\] _1698_ vssd1 vssd1 vccd1 vccd1 _1700_ sky130_fd_sc_hd__mux2_1
XANTENNA__2732__C1 _0806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3559_ _1585_ tms1x00.RAM\[51\]\[0\] _1659_ vssd1 vssd1 vccd1 vccd1 _1660_ sky130_fd_sc_hd__mux2_1
XFILLER_72_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2328__A tms1x00.Y\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3460__A0 _1585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2263__A1 net70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4465__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3763__A1 _1777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2723__C1 _0806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4808__CLK clknet_leaf_20_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2254__A1 K_override\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2672__S _0789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3451__A0 _1585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2930_ _1289_ vssd1 vssd1 vccd1 vccd1 _0084_ sky130_fd_sc_hd__clkbuf_1
XFILLER_22_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4600_ clknet_leaf_13_wb_clk_i _0221_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[125\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2861_ _1244_ vssd1 vssd1 vccd1 vccd1 _0060_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4958__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2792_ tms1x00.RAM\[28\]\[3\] tms1x00.RAM\[29\]\[3\] _0945_ vssd1 vssd1 vccd1 vccd1
+ _1182_ sky130_fd_sc_hd__mux2_1
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4531_ clknet_leaf_13_wb_clk_i _0152_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[110\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4462_ clknet_leaf_28_wb_clk_i _0083_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[59\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2701__A _0977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3413_ _1129_ vssd1 vssd1 vccd1 vccd1 _1576_ sky130_fd_sc_hd__clkbuf_4
X_4393_ clknet_leaf_34_wb_clk_i _0002_ vssd1 vssd1 vccd1 vccd1 tms1x00.wb_step sky130_fd_sc_hd__dfxtp_2
X_3344_ _1485_ tms1x00.RAM\[30\]\[0\] _1536_ vssd1 vssd1 vccd1 vccd1 _1537_ sky130_fd_sc_hd__mux2_1
XANTENNA__2190__A0 net40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3275_ _1497_ vssd1 vssd1 vccd1 vccd1 _0221_ sky130_fd_sc_hd__clkbuf_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5014_ clknet_leaf_12_wb_clk_i _0624_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[127\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_39_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2226_ net27 wbs_o_buff\[21\] _0679_ vssd1 vssd1 vccd1 vccd1 _0681_ sky130_fd_sc_hd__mux2_1
XFILLER_54_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3690__A0 _1710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2493__A1 _0819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4729_ clknet_leaf_3_wb_clk_i _0343_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[51\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2705__C1 _0775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_16_wb_clk_i_A clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_29_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3681__A0 _1710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3433__A0 _1588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3984__A1 tms1x00.ins_in\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2521__A _0913_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4068__A_N _0742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3060_ _1364_ tms1x00.RAM\[95\]\[1\] _1370_ vssd1 vssd1 vccd1 vccd1 _1372_ sky130_fd_sc_hd__mux2_1
XANTENNA__3352__A _1273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4630__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2475__A1 _0776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3672__A0 _1710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4183__A tms1x00.PC\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3962_ tms1x00.X\[0\] tms1x00.ram_addr_buff\[5\] _0725_ vssd1 vssd1 vccd1 vccd1 _1890_
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2913_ _1278_ vssd1 vssd1 vccd1 vccd1 _0078_ sky130_fd_sc_hd__clkbuf_1
X_3893_ _1852_ vssd1 vssd1 vccd1 vccd1 _0484_ sky130_fd_sc_hd__clkbuf_1
X_2844_ _1035_ tms1x00.RAM\[99\]\[1\] _1230_ vssd1 vssd1 vccd1 vccd1 _1232_ sky130_fd_sc_hd__mux2_1
X_4514_ clknet_leaf_14_wb_clk_i _0135_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[114\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_2775_ _0955_ tms1x00.RAM\[118\]\[3\] _0927_ vssd1 vssd1 vccd1 vccd1 _1165_ sky130_fd_sc_hd__o21a_1
XFILLER_8_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4445_ clknet_leaf_12_wb_clk_i _0066_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[17\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_4376_ _2171_ vssd1 vssd1 vccd1 vccd1 _0648_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__2389__S1 _0780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3327_ _1527_ vssd1 vssd1 vccd1 vccd1 _0243_ sky130_fd_sc_hd__clkbuf_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3258_ _1485_ tms1x00.RAM\[126\]\[0\] _1486_ vssd1 vssd1 vccd1 vccd1 _1487_ sky130_fd_sc_hd__mux2_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2209_ net18 wbs_o_buff\[13\] _0668_ vssd1 vssd1 vccd1 vccd1 _0672_ sky130_fd_sc_hd__mux2_1
XANTENNA__3663__A0 _1710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3189_ _1261_ _1430_ vssd1 vssd1 vccd1 vccd1 _1446_ sky130_fd_sc_hd__nor2_2
XFILLER_82_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2341__A _0718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4503__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4653__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3654__A0 _1710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5009__CLK clknet_leaf_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5099__A net52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output106_A net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2560_ tms1x00.RAM\[94\]\[1\] tms1x00.RAM\[95\]\[1\] _0923_ vssd1 vssd1 vccd1 vccd1
+ _0952_ sky130_fd_sc_hd__mux2_1
X_2491_ tms1x00.RAM\[40\]\[0\] tms1x00.RAM\[41\]\[0\] tms1x00.RAM\[42\]\[0\] tms1x00.RAM\[43\]\[0\]
+ _0777_ _0779_ vssd1 vssd1 vccd1 vccd1 _0884_ sky130_fd_sc_hd__mux4_1
X_4230_ tms1x00.X\[2\] _2087_ vssd1 vssd1 vccd1 vccd1 _2091_ sky130_fd_sc_hd__nand2_1
X_4161_ tms1x00.PC\[0\] _1908_ _2033_ _1966_ vssd1 vssd1 vccd1 vccd1 _0571_ sky130_fd_sc_hd__o211a_1
XANTENNA__2397__S _0789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4092_ _1981_ vssd1 vssd1 vccd1 vccd1 _0554_ sky130_fd_sc_hd__clkbuf_1
X_3112_ _1401_ vssd1 vssd1 vccd1 vccd1 _0154_ sky130_fd_sc_hd__clkbuf_1
XFILLER_56_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3043_ _1360_ vssd1 vssd1 vccd1 vccd1 _0126_ sky130_fd_sc_hd__clkbuf_1
XFILLER_49_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3645__A0 _1710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4994_ clknet_leaf_11_wb_clk_i _0604_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[29\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_36_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3948__A1 _1330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3945_ _1881_ vssd1 vssd1 vccd1 vccd1 _0507_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__3956__S _0726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3876_ tms1x00.RAM\[8\]\[2\] _1777_ _1840_ vssd1 vssd1 vccd1 vccd1 _1843_ sky130_fd_sc_hd__mux2_1
XANTENNA__3257__A _1430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2827_ _0783_ _1216_ vssd1 vssd1 vccd1 vccd1 _1217_ sky130_fd_sc_hd__or2_1
XANTENNA__4373__A1 _1333_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2758_ tms1x00.RAM\[72\]\[3\] tms1x00.RAM\[73\]\[3\] tms1x00.RAM\[74\]\[3\] tms1x00.RAM\[75\]\[3\]
+ _0799_ _0813_ vssd1 vssd1 vccd1 vccd1 _1148_ sky130_fd_sc_hd__mux4_1
X_2689_ _0920_ _1060_ _1066_ _1079_ _0773_ vssd1 vssd1 vccd1 vccd1 _1080_ sky130_fd_sc_hd__o311a_1
X_4428_ clknet_leaf_32_wb_clk_i net200 vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__dfxtp_1
XFILLER_59_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4359_ _2162_ vssd1 vssd1 vccd1 vccd1 _0640_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__2687__A1 _0807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_5_wb_clk_i clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__3636__A0 _1703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3939__A1 _1330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2611__A1 _0787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input67_A wbs_stb_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4116__A1 tms1x00.PA\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4549__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3730_ _1758_ vssd1 vssd1 vccd1 vccd1 _0415_ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4699__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3661_ _1708_ tms1x00.RAM\[67\]\[2\] _1717_ vssd1 vssd1 vccd1 vccd1 _1720_ sky130_fd_sc_hd__mux2_1
XFILLER_9_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2612_ _0928_ _1001_ _1003_ vssd1 vssd1 vccd1 vccd1 _1004_ sky130_fd_sc_hd__a21oi_1
X_3592_ tms1x00.RAM\[57\]\[1\] _1672_ _1678_ vssd1 vssd1 vccd1 vccd1 _1680_ sky130_fd_sc_hd__mux2_1
X_2543_ _0922_ _0926_ _0930_ _0934_ vssd1 vssd1 vccd1 vccd1 _0935_ sky130_fd_sc_hd__a31o_1
XANTENNA__2461__S0 _0815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2474_ _0863_ _0865_ _0866_ _0798_ _0802_ vssd1 vssd1 vccd1 vccd1 _0867_ sky130_fd_sc_hd__o221a_1
XFILLER_68_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4213_ tms1x00.Y\[2\] _2077_ _2063_ vssd1 vssd1 vccd1 vccd1 _2078_ sky130_fd_sc_hd__mux2_1
XANTENNA__2669__A1 _0948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4144_ _0743_ tms1x00.K_latch\[2\] _1956_ _1031_ vssd1 vssd1 vccd1 vccd1 _2019_ sky130_fd_sc_hd__a31o_1
XFILLER_56_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4075_ _0742_ tms1x00.status vssd1 vssd1 vccd1 vccd1 _1969_ sky130_fd_sc_hd__and2b_1
XFILLER_37_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3540__A _1240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3026_ _0913_ _1273_ vssd1 vssd1 vccd1 vccd1 _1351_ sky130_fd_sc_hd__or2_2
XFILLER_55_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4977_ clknet_leaf_9_wb_clk_i _0587_ vssd1 vssd1 vccd1 vccd1 tms1x00.N\[3\] sky130_fd_sc_hd__dfxtp_1
X_3928_ tms1x00.RAM\[91\]\[1\] _1775_ _1870_ vssd1 vssd1 vccd1 vccd1 _1872_ sky130_fd_sc_hd__mux2_1
X_3859_ _1833_ vssd1 vssd1 vccd1 vccd1 _0469_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2452__S0 _0815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3450__A _0917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2691__S0 _0873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4991__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2443__S0 _0799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3625__A _1284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2190_ net40 wbs_o_buff\[4\] _0657_ vssd1 vssd1 vccd1 vccd1 _0662_ sky130_fd_sc_hd__mux2_1
XFILLER_77_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4900_ clknet_leaf_10_wb_clk_i _0514_ vssd1 vssd1 vccd1 vccd1 tms1x00.ram_addr_buff\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_46_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4831_ clknet_leaf_19_wb_clk_i _0445_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[78\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_34_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4191__A _0748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4762_ clknet_leaf_20_wb_clk_i _0376_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[61\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_4693_ clknet_leaf_32_wb_clk_i _0307_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[42\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2682__S0 _0830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3713_ tms1x00.RAM\[70\]\[1\] _1672_ _1747_ vssd1 vssd1 vccd1 vccd1 _1749_ sky130_fd_sc_hd__mux2_1
X_3644_ _1224_ vssd1 vssd1 vccd1 vccd1 _1710_ sky130_fd_sc_hd__clkbuf_4
X_3575_ _1668_ vssd1 vssd1 vccd1 vccd1 _0350_ sky130_fd_sc_hd__clkbuf_1
X_2526_ _0912_ tms1x00.RAM\[109\]\[0\] _0918_ vssd1 vssd1 vccd1 vccd1 _0919_ sky130_fd_sc_hd__mux2_1
XANTENNA__3839__A0 _1821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2457_ _0779_ vssd1 vssd1 vccd1 vccd1 _0850_ sky130_fd_sc_hd__buf_6
XFILLER_69_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4714__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2388_ tms1x00.RAM\[80\]\[0\] tms1x00.RAM\[81\]\[0\] tms1x00.RAM\[82\]\[0\] tms1x00.RAM\[83\]\[0\]
+ _0778_ _0780_ vssd1 vssd1 vccd1 vccd1 _0781_ sky130_fd_sc_hd__mux4_1
XFILLER_29_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4127_ _2004_ vssd1 vssd1 vccd1 vccd1 _0566_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4366__A _1261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4085__B _0738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4058_ tms1x00.ins_in\[4\] _0749_ vssd1 vssd1 vccd1 vccd1 _1956_ sky130_fd_sc_hd__nor2_2
XFILLER_43_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3009_ _1340_ vssd1 vssd1 vccd1 vccd1 _0112_ sky130_fd_sc_hd__clkbuf_1
XFILLER_52_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3429__B _1343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4276__A _0917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3180__A _1430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3230__A1 _1456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2416__S0 _0808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output98_A net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3360_ _1545_ vssd1 vssd1 vccd1 vccd1 _0258_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4737__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2311_ tms1x00.wb_step _0713_ _0714_ _0716_ net63 vssd1 vssd1 vccd1 vccd1 _0002_
+ sky130_fd_sc_hd__a32o_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5030_ clknet_leaf_20_wb_clk_i _0640_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[14\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_3291_ _1506_ vssd1 vssd1 vccd1 vccd1 _0228_ sky130_fd_sc_hd__clkbuf_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2242_ net35 wbs_o_buff\[29\] _0679_ vssd1 vssd1 vccd1 vccd1 _0689_ sky130_fd_sc_hd__mux2_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4887__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4814_ clknet_leaf_22_wb_clk_i _0428_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[74\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_4745_ clknet_leaf_26_wb_clk_i _0359_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[56\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3221__A1 _1456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4676_ clknet_leaf_11_wb_clk_i _0048_ vssd1 vssd1 vccd1 vccd1 _0041_ sky130_fd_sc_hd__dfxtp_1
X_3627_ _1699_ vssd1 vssd1 vccd1 vccd1 _0371_ sky130_fd_sc_hd__clkbuf_1
X_3558_ _1229_ _1283_ vssd1 vssd1 vccd1 vccd1 _1659_ sky130_fd_sc_hd__or2_2
X_2509_ _0039_ _0886_ _0890_ _0901_ _0040_ vssd1 vssd1 vccd1 vccd1 _0902_ sky130_fd_sc_hd__o311a_1
XFILLER_1_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3489_ _1588_ tms1x00.RAM\[50\]\[1\] _1619_ vssd1 vssd1 vccd1 vccd1 _1621_ sky130_fd_sc_hd__mux2_1
XFILLER_57_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3288__A1 _1456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5042__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2799__B1 _0794_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2344__A tms1x00.Y\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2646__S0 _0955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3212__A1 _1459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2584__B_N _0975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3279__A1 _1456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2519__A _0911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2860_ tms1x00.RAM\[69\]\[1\] _1243_ _1241_ vssd1 vssd1 vccd1 vccd1 _1244_ sky130_fd_sc_hd__mux2_1
XFILLER_30_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2791_ _0928_ _1180_ vssd1 vssd1 vccd1 vccd1 _1181_ sky130_fd_sc_hd__and2_1
XANTENNA__3203__A1 _1331_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4530_ clknet_leaf_13_wb_clk_i _0151_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[110\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4461_ clknet_leaf_34_wb_clk_i _0082_ vssd1 vssd1 vccd1 vccd1 K_override\[3\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__3085__A _1345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3412_ _1575_ vssd1 vssd1 vccd1 vccd1 _0280_ sky130_fd_sc_hd__clkbuf_1
X_4392_ clknet_leaf_33_wb_clk_i _0000_ vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__dfxtp_4
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3343_ _1249_ _1396_ vssd1 vssd1 vccd1 vccd1 _1536_ sky130_fd_sc_hd__or2_2
XANTENNA__3813__A _1240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3274_ _1490_ tms1x00.RAM\[125\]\[2\] _1494_ vssd1 vssd1 vccd1 vccd1 _1497_ sky130_fd_sc_hd__mux2_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5013_ clknet_leaf_20_wb_clk_i _0623_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[12\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2429__A _0812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2225_ _0680_ vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__clkbuf_1
XANTENNA__4219__A0 _0732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2493__A2 _0883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3442__A1 _1571_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4902__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2989_ tms1x00.RAM\[101\]\[0\] _1324_ _1325_ vssd1 vssd1 vccd1 vccd1 _1326_ sky130_fd_sc_hd__mux2_1
XFILLER_21_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4728_ clknet_leaf_29_wb_clk_i _0342_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[52\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_4659_ clknet_leaf_32_wb_clk_i _0280_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[41\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2800__S0 _0816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3130__A0 _1366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3984__A2 _0724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4582__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_1_wb_clk_i_A clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_5_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3352__B _1343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_29_wb_clk_i clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_75_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3961_ _1889_ vssd1 vssd1 vccd1 vccd1 _0515_ sky130_fd_sc_hd__clkbuf_1
XFILLER_50_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3424__A1 _1576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2912_ _1225_ tms1x00.RAM\[18\]\[3\] _1274_ vssd1 vssd1 vccd1 vccd1 _1278_ sky130_fd_sc_hd__mux2_1
XFILLER_32_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3892_ tms1x00.RAM\[87\]\[1\] _1775_ _1850_ vssd1 vssd1 vccd1 vccd1 _1852_ sky130_fd_sc_hd__mux2_1
XANTENNA__2632__C1 _0794_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2843_ _1231_ vssd1 vssd1 vccd1 vccd1 _0055_ sky130_fd_sc_hd__clkbuf_1
X_2774_ tms1x00.RAM\[119\]\[3\] _0955_ vssd1 vssd1 vccd1 vccd1 _1164_ sky130_fd_sc_hd__or2b_1
XANTENNA__2712__A _0821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4513_ clknet_leaf_17_wb_clk_i _0134_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[95\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_4444_ clknet_leaf_12_wb_clk_i _0065_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[17\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_4375_ tms1x00.PC\[2\] net95 _2006_ vssd1 vssd1 vccd1 vccd1 _2171_ sky130_fd_sc_hd__mux2_1
XANTENNA__2699__C1 _0942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3326_ _1485_ tms1x00.RAM\[32\]\[0\] _1526_ vssd1 vssd1 vccd1 vccd1 _1527_ sky130_fd_sc_hd__mux2_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4455__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3257_ _1430_ _1396_ vssd1 vssd1 vccd1 vccd1 _1486_ sky130_fd_sc_hd__or2_2
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2208_ _0671_ vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__clkbuf_1
X_3188_ _1445_ vssd1 vssd1 vccd1 vccd1 _0186_ sky130_fd_sc_hd__clkbuf_1
XFILLER_66_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input12_A oram_value[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2532__A _0923_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output80_A net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2490_ tms1x00.RAM\[44\]\[0\] tms1x00.RAM\[45\]\[0\] tms1x00.RAM\[46\]\[0\] tms1x00.RAM\[47\]\[0\]
+ _0808_ _0831_ vssd1 vssd1 vccd1 vccd1 _0883_ sky130_fd_sc_hd__mux4_2
XFILLER_5_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2678__S _0823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4160_ _2025_ _2032_ _1908_ vssd1 vssd1 vccd1 vccd1 _2033_ sky130_fd_sc_hd__o21ai_1
XFILLER_4_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3111_ _1368_ tms1x00.RAM\[110\]\[3\] _1397_ vssd1 vssd1 vccd1 vccd1 _1401_ sky130_fd_sc_hd__mux2_1
XFILLER_1_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4091_ tms1x00.SR\[1\] tms1x00.PC\[1\] _1979_ vssd1 vssd1 vccd1 vccd1 _1981_ sky130_fd_sc_hd__mux2_1
X_3042_ _1225_ tms1x00.RAM\[97\]\[3\] _1356_ vssd1 vssd1 vccd1 vccd1 _1360_ sky130_fd_sc_hd__mux2_1
XFILLER_49_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4993_ clknet_leaf_0_wb_clk_i _0603_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[22\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_51_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3944_ tms1x00.RAM\[23\]\[0\] _1323_ _1880_ vssd1 vssd1 vccd1 vccd1 _1881_ sky130_fd_sc_hd__mux2_1
XFILLER_20_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3875_ _1842_ vssd1 vssd1 vccd1 vccd1 _0476_ sky130_fd_sc_hd__clkbuf_1
X_2826_ tms1x00.RAM\[56\]\[3\] tms1x00.RAM\[57\]\[3\] tms1x00.RAM\[58\]\[3\] tms1x00.RAM\[59\]\[3\]
+ _0826_ _0850_ vssd1 vssd1 vccd1 vccd1 _1216_ sky130_fd_sc_hd__mux4_1
XANTENNA__3257__B _1396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2908__A0 _1035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2757_ _1143_ _1145_ _1146_ _0807_ _0775_ vssd1 vssd1 vccd1 vccd1 _1147_ sky130_fd_sc_hd__o221a_1
X_2688_ _0039_ _1072_ _1078_ vssd1 vssd1 vccd1 vccd1 _1079_ sky130_fd_sc_hd__or3_1
X_4427_ clknet_leaf_27_wb_clk_i _0027_ vssd1 vssd1 vccd1 vccd1 wbs_o_buff\[31\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_input4_A io_in[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4358_ _1235_ tms1x00.RAM\[14\]\[0\] _2161_ vssd1 vssd1 vccd1 vccd1 _2162_ sky130_fd_sc_hd__mux2_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3309_ _1516_ vssd1 vssd1 vccd1 vccd1 _0236_ sky130_fd_sc_hd__clkbuf_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4289_ _2123_ vssd1 vssd1 vccd1 vccd1 _0609_ sky130_fd_sc_hd__clkbuf_1
XFILLER_73_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2617__A _0953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4620__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4429__D valid vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3660_ _1719_ vssd1 vssd1 vccd1 vccd1 _0384_ sky130_fd_sc_hd__clkbuf_1
X_2611_ _0787_ _1002_ _0996_ vssd1 vssd1 vccd1 vccd1 _1003_ sky130_fd_sc_hd__a21o_1
X_3591_ _1679_ vssd1 vssd1 vccd1 vccd1 _0355_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3563__A0 _1590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2542_ _0922_ _0933_ _0776_ vssd1 vssd1 vccd1 vccd1 _0934_ sky130_fd_sc_hd__o21ai_1
XANTENNA__2461__S1 _0812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4212_ _2075_ _2076_ vssd1 vssd1 vccd1 vccd1 _2077_ sky130_fd_sc_hd__xnor2_1
X_2473_ tms1x00.RAM\[24\]\[0\] tms1x00.RAM\[25\]\[0\] tms1x00.RAM\[26\]\[0\] tms1x00.RAM\[27\]\[0\]
+ _0830_ _0800_ vssd1 vssd1 vccd1 vccd1 _0866_ sky130_fd_sc_hd__mux4_2
XFILLER_68_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2669__A2 _1057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4143_ _2009_ _1126_ vssd1 vssd1 vccd1 vccd1 _2018_ sky130_fd_sc_hd__and2b_1
XFILLER_29_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4074_ _1958_ _1967_ _1968_ _1966_ vssd1 vssd1 vccd1 vccd1 _0549_ sky130_fd_sc_hd__o211a_1
XFILLER_55_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3025_ _1350_ vssd1 vssd1 vccd1 vccd1 _0118_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__3540__B _1284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2437__A _0777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4976_ clknet_leaf_9_wb_clk_i _0586_ vssd1 vssd1 vccd1 vccd1 tms1x00.N\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3927_ _1871_ vssd1 vssd1 vccd1 vccd1 _0499_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4643__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3858_ _1821_ tms1x00.RAM\[81\]\[2\] _1830_ vssd1 vssd1 vccd1 vccd1 _1833_ sky130_fd_sc_hd__mux2_1
XFILLER_50_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2809_ _0920_ _1179_ _1185_ _1198_ _0773_ vssd1 vssd1 vccd1 vccd1 _1199_ sky130_fd_sc_hd__o311a_1
X_3789_ tms1x00.RAM\[7\]\[1\] _1775_ _1791_ vssd1 vssd1 vccd1 vccd1 _1793_ sky130_fd_sc_hd__mux2_1
XANTENNA__4793__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2452__S1 _0812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2817__C1 _0806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2691__S1 _0977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2443__S1 _0800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3625__B _1396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3641__A _1129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2257__A net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4666__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2284__B1 _0703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4830_ clknet_leaf_20_wb_clk_i _0444_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[78\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_34_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4191__B tms1x00.ins_in\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3784__A0 _1710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4761_ clknet_leaf_20_wb_clk_i _0375_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[61\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_4692_ clknet_leaf_32_wb_clk_i _0306_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[43\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_3712_ _1748_ vssd1 vssd1 vccd1 vccd1 _0407_ sky130_fd_sc_hd__clkbuf_1
X_3643_ _1709_ vssd1 vssd1 vccd1 vccd1 _0377_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__2682__S1 _0800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3574_ tms1x00.RAM\[5\]\[3\] _1578_ _1664_ vssd1 vssd1 vccd1 vccd1 _1668_ sky130_fd_sc_hd__mux2_1
X_2525_ _0914_ _0917_ vssd1 vssd1 vccd1 vccd1 _0918_ sky130_fd_sc_hd__or2_2
X_2456_ tms1x00.RAM\[119\]\[0\] _0808_ vssd1 vssd1 vccd1 vccd1 _0849_ sky130_fd_sc_hd__or2b_1
XFILLER_69_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4126_ _0738_ _2003_ vssd1 vssd1 vccd1 vccd1 _2004_ sky130_fd_sc_hd__or2_1
XFILLER_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2387_ _0779_ vssd1 vssd1 vccd1 vccd1 _0780_ sky130_fd_sc_hd__buf_6
XFILLER_68_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4366__B _1344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4057_ _0753_ _1954_ _1955_ _1931_ vssd1 vssd1 vccd1 vccd1 _0545_ sky130_fd_sc_hd__o211a_1
XFILLER_71_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2275__B1 _0703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3008_ tms1x00.RAM\[100\]\[1\] _1328_ _1338_ vssd1 vssd1 vccd1 vccd1 _1340_ sky130_fd_sc_hd__mux2_1
XFILLER_61_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4959_ clknet_leaf_9_wb_clk_i _0569_ vssd1 vssd1 vccd1 vccd1 tms1x00.P\[2\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__3527__A0 _1590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_35_wb_clk_i_A clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_10_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2776__S _0789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4276__B _1249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4689__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3180__B _1403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3518__A0 _1590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2540__A _0822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2416__S1 _0780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3290_ tms1x00.RAM\[24\]\[1\] _1459_ _1504_ vssd1 vssd1 vccd1 vccd1 _1506_ sky130_fd_sc_hd__mux2_1
XFILLER_3_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2310_ wb_rst_override _0713_ _0714_ _0716_ net62 vssd1 vssd1 vccd1 vccd1 _0001_
+ sky130_fd_sc_hd__a32o_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2241_ _0688_ vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__clkbuf_1
XFILLER_66_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3310__S _1514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4813_ clknet_leaf_24_wb_clk_i _0427_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[74\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_4744_ clknet_leaf_26_wb_clk_i _0358_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[57\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3509__A0 _1590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4675_ clknet_leaf_11_wb_clk_i _0047_ vssd1 vssd1 vccd1 vccd1 _0040_ sky130_fd_sc_hd__dfxtp_4
XANTENNA__2980__A1 _1243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3626_ _1585_ tms1x00.RAM\[62\]\[0\] _1698_ vssd1 vssd1 vccd1 vccd1 _1699_ sky130_fd_sc_hd__mux2_1
XANTENNA__2450__A _0828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3557_ _1658_ vssd1 vssd1 vccd1 vccd1 _0342_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__2732__A1 _0996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2508_ _0892_ _0894_ _0898_ _0900_ _0804_ vssd1 vssd1 vccd1 vccd1 _0901_ sky130_fd_sc_hd__a221o_1
XFILLER_0_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3488_ _1620_ vssd1 vssd1 vccd1 vccd1 _0311_ sky130_fd_sc_hd__clkbuf_1
XFILLER_69_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2439_ tms1x00.RAM\[64\]\[0\] tms1x00.RAM\[65\]\[0\] tms1x00.RAM\[66\]\[0\] tms1x00.RAM\[67\]\[0\]
+ _0830_ _0831_ vssd1 vssd1 vccd1 vccd1 _0832_ sky130_fd_sc_hd__mux4_1
XFILLER_56_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4109_ net103 _1991_ vssd1 vssd1 vccd1 vccd1 _1992_ sky130_fd_sc_hd__or2_1
XFILLER_45_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4981__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2799__A1 _0818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2646__S1 _0956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2971__A1 _1245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2723__A1 _0996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input42_A ram_val[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2582__S0 _0955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2535__A _0850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2790_ tms1x00.RAM\[30\]\[3\] tms1x00.RAM\[31\]\[3\] _0945_ vssd1 vssd1 vccd1 vccd1
+ _1180_ sky130_fd_sc_hd__mux2_1
XANTENNA__4704__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2962__A1 _1247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4460_ clknet_leaf_32_wb_clk_i _0081_ vssd1 vssd1 vccd1 vccd1 K_override\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_7_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3085__B _1375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4854__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4391_ clknet_leaf_9_wb_clk_i _0049_ vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__dfxtp_2
X_3411_ tms1x00.RAM\[41\]\[1\] _1574_ _1572_ vssd1 vssd1 vccd1 vccd1 _1575_ sky130_fd_sc_hd__mux2_1
X_3342_ _1535_ vssd1 vssd1 vccd1 vccd1 _0250_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__3813__B _1258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3273_ _1496_ vssd1 vssd1 vccd1 vccd1 _0220_ sky130_fd_sc_hd__clkbuf_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5012_ clknet_leaf_20_wb_clk_i _0622_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[12\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2224_ net26 wbs_o_buff\[20\] _0679_ vssd1 vssd1 vccd1 vccd1 _0680_ sky130_fd_sc_hd__mux2_1
XANTENNA__2573__S0 _0955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2988_ _0914_ _1240_ vssd1 vssd1 vccd1 vccd1 _1325_ sky130_fd_sc_hd__nor2_2
XANTENNA__2402__B1 _0794_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4727_ clknet_leaf_29_wb_clk_i _0341_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[52\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_4658_ clknet_leaf_32_wb_clk_i _0279_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[41\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_3609_ _1689_ vssd1 vssd1 vccd1 vccd1 _0363_ sky130_fd_sc_hd__clkbuf_1
X_4589_ clknet_leaf_2_wb_clk_i _0210_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[116\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2705__B2 _0798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2800__S1 _0977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3969__A0 net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2355__A tms1x00.ins_in\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2555__S0 _0945_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3960_ tms1x00.X\[2\] tms1x00.ram_addr_buff\[4\] _0725_ vssd1 vssd1 vccd1 vccd1 _1889_
+ sky130_fd_sc_hd__mux2_1
X_2911_ _1277_ vssd1 vssd1 vccd1 vccd1 _0077_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4196__D_N tms1x00.ins_in\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3891_ _1851_ vssd1 vssd1 vccd1 vccd1 _0483_ sky130_fd_sc_hd__clkbuf_1
X_2842_ _0912_ tms1x00.RAM\[99\]\[0\] _1230_ vssd1 vssd1 vccd1 vccd1 _1231_ sky130_fd_sc_hd__mux2_1
X_2773_ _0922_ _1160_ _1162_ _0944_ vssd1 vssd1 vccd1 vccd1 _1163_ sky130_fd_sc_hd__o211a_1
X_4512_ clknet_leaf_17_wb_clk_i _0133_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[95\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4443_ clknet_leaf_12_wb_clk_i _0064_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[17\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__5032__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4374_ _2170_ vssd1 vssd1 vccd1 vccd1 _0647_ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3325_ _1345_ _1525_ vssd1 vssd1 vccd1 vccd1 _1526_ sky130_fd_sc_hd__or2_2
XANTENNA__2794__S0 _0924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3256_ _0911_ vssd1 vssd1 vccd1 vccd1 _1485_ sky130_fd_sc_hd__clkbuf_4
XFILLER_39_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2207_ net17 wbs_o_buff\[12\] _0668_ vssd1 vssd1 vccd1 vccd1 _0671_ sky130_fd_sc_hd__mux2_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3187_ tms1x00.RAM\[122\]\[3\] _1334_ _1441_ vssd1 vssd1 vccd1 vccd1 _1445_ sky130_fd_sc_hd__mux2_1
XFILLER_27_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2623__B1 _0775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4064__C1 _1931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2614__B1 _0942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2813__A _0921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3590__A1 _1669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3644__A _1224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output73_A net73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3110_ _1400_ vssd1 vssd1 vccd1 vccd1 _0153_ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4090_ _1980_ vssd1 vssd1 vccd1 vccd1 _0553_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2694__S _0789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3041_ _1359_ vssd1 vssd1 vccd1 vccd1 _0125_ sky130_fd_sc_hd__clkbuf_1
XFILLER_76_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4992_ clknet_leaf_0_wb_clk_i _0602_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[22\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_3943_ _1250_ _1310_ vssd1 vssd1 vccd1 vccd1 _1880_ sky130_fd_sc_hd__nor2_2
XANTENNA__2605__B1 _0996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3874_ tms1x00.RAM\[8\]\[1\] _1775_ _1840_ vssd1 vssd1 vccd1 vccd1 _1842_ sky130_fd_sc_hd__mux2_1
XFILLER_20_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2825_ tms1x00.RAM\[60\]\[3\] tms1x00.RAM\[61\]\[3\] tms1x00.RAM\[62\]\[3\] tms1x00.RAM\[63\]\[3\]
+ _0923_ _0927_ vssd1 vssd1 vccd1 vccd1 _1215_ sky130_fd_sc_hd__mux4_1
XANTENNA__4358__A0 _1235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2756_ tms1x00.RAM\[64\]\[3\] tms1x00.RAM\[65\]\[3\] tms1x00.RAM\[66\]\[3\] tms1x00.RAM\[67\]\[3\]
+ _0830_ _0831_ vssd1 vssd1 vccd1 vccd1 _1146_ sky130_fd_sc_hd__mux4_1
X_2687_ _0807_ _1073_ _1077_ _0802_ vssd1 vssd1 vccd1 vccd1 _1078_ sky130_fd_sc_hd__o211a_1
XANTENNA__3581__A1 _1672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4426_ clknet_leaf_27_wb_clk_i _0026_ vssd1 vssd1 vccd1 vccd1 wbs_o_buff\[30\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__2767__S0 _0840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4357_ _1343_ _1396_ vssd1 vssd1 vccd1 vccd1 _2161_ sky130_fd_sc_hd__or2_2
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4572__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3308_ tms1x00.RAM\[27\]\[1\] _1459_ _1514_ vssd1 vssd1 vccd1 vccd1 _1516_ sky130_fd_sc_hd__mux2_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4288_ tms1x00.RAM\[21\]\[1\] _1327_ _2121_ vssd1 vssd1 vccd1 vccd1 _2123_ sky130_fd_sc_hd__mux2_1
XANTENNA__3097__A0 _1364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3239_ tms1x00.RAM\[116\]\[0\] _1456_ _1475_ vssd1 vssd1 vccd1 vccd1 _1476_ sky130_fd_sc_hd__mux2_1
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2844__A0 _1035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2617__B _1008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4349__A0 _1235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3572__A1 _1576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4915__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2758__S0 _0799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3088__A0 _1364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2808__A _0821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4037__C1 _1931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output111_A net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4002__A_N tms1x00.Y\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4445__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2610_ tms1x00.RAM\[12\]\[1\] tms1x00.RAM\[13\]\[1\] _0975_ vssd1 vssd1 vccd1 vccd1
+ _1002_ sky130_fd_sc_hd__mux2_1
X_3590_ tms1x00.RAM\[57\]\[0\] _1669_ _1678_ vssd1 vssd1 vccd1 vccd1 _1679_ sky130_fd_sc_hd__mux2_1
X_2541_ tms1x00.RAM\[64\]\[1\] tms1x00.RAM\[65\]\[1\] tms1x00.RAM\[66\]\[1\] tms1x00.RAM\[67\]\[1\]
+ _0931_ _0932_ vssd1 vssd1 vccd1 vccd1 _0933_ sky130_fd_sc_hd__mux4_1
XANTENNA__4595__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2472_ _0786_ _0864_ _0828_ vssd1 vssd1 vccd1 vccd1 _0865_ sky130_fd_sc_hd__a21o_1
XFILLER_5_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4211_ _2067_ _2069_ _2066_ vssd1 vssd1 vccd1 vccd1 _2076_ sky130_fd_sc_hd__a21boi_1
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3315__A1 _1456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4142_ tms1x00.P\[1\] _2007_ _2015_ _2017_ vssd1 vssd1 vccd1 vccd1 _0568_ sky130_fd_sc_hd__o22a_1
XANTENNA__3079__A0 _1364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4073_ net72 _1960_ vssd1 vssd1 vccd1 vccd1 _1968_ sky130_fd_sc_hd__or2_1
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3024_ _1225_ tms1x00.RAM\[0\]\[3\] _1346_ vssd1 vssd1 vccd1 vccd1 _1350_ sky130_fd_sc_hd__mux2_1
XFILLER_36_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_13_wb_clk_i clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_36_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4975_ clknet_leaf_8_wb_clk_i _0585_ vssd1 vssd1 vccd1 vccd1 tms1x00.N\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_52_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3549__A _1284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3926_ tms1x00.RAM\[91\]\[0\] _1772_ _1870_ vssd1 vssd1 vccd1 vccd1 _1871_ sky130_fd_sc_hd__mux2_1
X_3857_ _1832_ vssd1 vssd1 vccd1 vccd1 _0468_ sky130_fd_sc_hd__clkbuf_1
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2808_ _0821_ _1191_ _1197_ vssd1 vssd1 vccd1 vccd1 _1198_ sky130_fd_sc_hd__or3_1
X_3788_ _1792_ vssd1 vssd1 vccd1 vccd1 _0439_ sky130_fd_sc_hd__clkbuf_1
X_2739_ _1129_ vssd1 vssd1 vccd1 vccd1 _1130_ sky130_fd_sc_hd__buf_4
XFILLER_4_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3554__A1 _1576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_25_wb_clk_i_A clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__2762__C1 _0828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3306__A1 _1456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4409_ clknet_leaf_28_wb_clk_i _0007_ vssd1 vssd1 vccd1 vccd1 wbs_o_buff\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_75_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4468__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3459__A _1409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3793__A1 _1779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3545__A1 _1576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2505__C1 _0828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2538__A _0928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2257__B net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2284__A1 net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2273__A _0697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4760_ clknet_leaf_10_wb_clk_i _0374_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[62\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4691_ clknet_leaf_31_wb_clk_i _0305_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[43\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_3711_ tms1x00.RAM\[70\]\[0\] _1669_ _1747_ vssd1 vssd1 vccd1 vccd1 _1748_ sky130_fd_sc_hd__mux2_1
X_3642_ _1708_ tms1x00.RAM\[61\]\[2\] _1704_ vssd1 vssd1 vccd1 vccd1 _1709_ sky130_fd_sc_hd__mux2_1
XANTENNA__3536__A1 _1576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3308__S _1514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3573_ _1667_ vssd1 vssd1 vccd1 vccd1 _0349_ sky130_fd_sc_hd__clkbuf_1
X_2524_ _0728_ _0916_ _0717_ vssd1 vssd1 vccd1 vccd1 _0917_ sky130_fd_sc_hd__nand3b_4
X_2455_ _0794_ _0847_ _0038_ vssd1 vssd1 vccd1 vccd1 _0848_ sky130_fd_sc_hd__o21a_1
XANTENNA__3832__A _1229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2386_ _0036_ vssd1 vssd1 vccd1 vccd1 _0779_ sky130_fd_sc_hd__clkbuf_8
XFILLER_69_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4125_ tms1x00.PB\[3\] tms1x00.PA\[3\] _1996_ vssd1 vssd1 vccd1 vccd1 _2003_ sky130_fd_sc_hd__mux2_1
XFILLER_56_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4056_ _0733_ _0764_ _1935_ net92 vssd1 vssd1 vccd1 vccd1 _1955_ sky130_fd_sc_hd__a31o_1
XFILLER_45_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2275__A1 net79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3007_ _1339_ vssd1 vssd1 vccd1 vccd1 _0111_ sky130_fd_sc_hd__clkbuf_1
XFILLER_25_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4958_ clknet_leaf_8_wb_clk_i _0568_ vssd1 vssd1 vccd1 vccd1 tms1x00.P\[1\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__4760__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3909_ _1861_ vssd1 vssd1 vccd1 vccd1 _0491_ sky130_fd_sc_hd__clkbuf_1
X_4889_ clknet_leaf_30_wb_clk_i _0503_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[90\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3775__A1 _1779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2750__A2 tms1x00.RAM\[90\]\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2358__A _0752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_2_1__f_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2792__S _0945_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2266__A1 net73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3189__A _1261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3766__A1 _1779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2240_ net34 wbs_o_buff\[28\] _0679_ vssd1 vssd1 vccd1 vccd1 _0688_ sky130_fd_sc_hd__mux2_1
XANTENNA__4633__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2207__S _0668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4812_ clknet_leaf_24_wb_clk_i _0426_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[75\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3757__A1 _1772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4743_ clknet_leaf_28_wb_clk_i _0357_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[57\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2731__A _0783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4674_ clknet_leaf_9_wb_clk_i _0046_ vssd1 vssd1 vccd1 vccd1 _0039_ sky130_fd_sc_hd__dfxtp_1
X_3625_ _1284_ _1396_ vssd1 vssd1 vccd1 vccd1 _1698_ sky130_fd_sc_hd__or2_2
XANTENNA__2717__C1 _0953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3556_ tms1x00.RAM\[52\]\[3\] _1578_ _1654_ vssd1 vssd1 vccd1 vccd1 _1658_ sky130_fd_sc_hd__mux2_1
X_2507_ _0797_ _0899_ _0774_ vssd1 vssd1 vccd1 vccd1 _0900_ sky130_fd_sc_hd__o21a_1
X_3487_ _1585_ tms1x00.RAM\[50\]\[0\] _1619_ vssd1 vssd1 vccd1 vccd1 _1620_ sky130_fd_sc_hd__mux2_1
X_2438_ _0779_ vssd1 vssd1 vccd1 vccd1 _0831_ sky130_fd_sc_hd__buf_6
XFILLER_69_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2369_ _0763_ vssd1 vssd1 vccd1 vccd1 _0764_ sky130_fd_sc_hd__buf_2
XFILLER_57_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4108_ tms1x00.PA\[2\] _1973_ _1987_ tms1x00.PB\[2\] vssd1 vssd1 vccd1 vccd1 _1991_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__2248__A1 K_override\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4039_ _0733_ _0739_ _0764_ _1918_ net87 vssd1 vssd1 vccd1 vccd1 _1943_ sky130_fd_sc_hd__a41o_1
XFILLER_56_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4506__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3737__A _1236_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2184__A0 net25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4656__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input35_A ram_val[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3684__A0 _1703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2582__S1 _0956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3436__A0 _1590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2816__A _0783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3647__A _1283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4390_ _2178_ vssd1 vssd1 vccd1 vccd1 _0655_ sky130_fd_sc_hd__clkbuf_1
X_3410_ _1034_ vssd1 vssd1 vccd1 vccd1 _1574_ sky130_fd_sc_hd__clkbuf_4
X_3341_ _1492_ tms1x00.RAM\[31\]\[3\] _1531_ vssd1 vssd1 vccd1 vccd1 _1535_ sky130_fd_sc_hd__mux2_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3272_ _1488_ tms1x00.RAM\[125\]\[1\] _1494_ vssd1 vssd1 vccd1 vccd1 _1496_ sky130_fd_sc_hd__mux2_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5011_ clknet_leaf_12_wb_clk_i _0621_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[12\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2223_ net49 vssd1 vssd1 vccd1 vccd1 _0679_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__3675__A0 _1703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2573__S1 _0956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3321__S _1519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5102__A net55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2726__A _0953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2987_ _1323_ vssd1 vssd1 vccd1 vccd1 _1324_ sky130_fd_sc_hd__buf_2
XANTENNA__2402__A1 _0791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4726_ clknet_leaf_28_wb_clk_i _0340_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[52\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_4657_ clknet_leaf_6_wb_clk_i _0278_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[33\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4679__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3608_ tms1x00.RAM\[55\]\[0\] _1669_ _1688_ vssd1 vssd1 vccd1 vccd1 _1689_ sky130_fd_sc_hd__mux2_1
X_4588_ clknet_leaf_1_wb_clk_i _0209_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[116\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_3539_ _1648_ vssd1 vssd1 vccd1 vccd1 _0334_ sky130_fd_sc_hd__clkbuf_1
XFILLER_76_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3666__A0 _1703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2636__A _0773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2371__A _0718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3657__A0 _1703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2555__S1 _0791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2910_ _1130_ tms1x00.RAM\[18\]\[2\] _1274_ vssd1 vssd1 vccd1 vccd1 _1277_ sky130_fd_sc_hd__mux2_1
XFILLER_32_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3890_ tms1x00.RAM\[87\]\[0\] _1772_ _1850_ vssd1 vssd1 vccd1 vccd1 _1851_ sky130_fd_sc_hd__mux2_1
XANTENNA__2632__B2 _0818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2841_ _0914_ _1229_ vssd1 vssd1 vccd1 vccd1 _1230_ sky130_fd_sc_hd__or2_2
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2772_ _0996_ _1161_ vssd1 vssd1 vccd1 vccd1 _1162_ sky130_fd_sc_hd__or2_1
XFILLER_12_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4511_ clknet_leaf_15_wb_clk_i _0132_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[95\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4137__A1 tms1x00.ins_in\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4442_ clknet_leaf_12_wb_clk_i _0063_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[17\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2491__S0 _0777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4971__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4373_ tms1x00.RAM\[9\]\[3\] _1333_ _2166_ vssd1 vssd1 vccd1 vccd1 _2170_ sky130_fd_sc_hd__mux2_1
XANTENNA__2699__B2 _0922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4001__A net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3324_ _1524_ vssd1 vssd1 vccd1 vccd1 _1525_ sky130_fd_sc_hd__buf_4
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2794__S1 _0928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3255_ _1484_ vssd1 vssd1 vccd1 vccd1 _0214_ sky130_fd_sc_hd__clkbuf_1
XFILLER_58_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3648__A0 _1703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2206_ _0670_ vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__clkbuf_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3186_ _1444_ vssd1 vssd1 vccd1 vccd1 _0185_ sky130_fd_sc_hd__clkbuf_1
XFILLER_81_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2623__A1 _0819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3287__A _1250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4709_ clknet_leaf_3_wb_clk_i _0323_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[47\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3639__A0 _1706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2366__A _0760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3811__A0 _1710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2614__A1 _0948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2813__B _1202_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4367__A1 _1323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2473__S0 _0830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3925__A _1258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3040_ _1130_ tms1x00.RAM\[97\]\[2\] _1356_ vssd1 vssd1 vccd1 vccd1 _1359_ sky130_fd_sc_hd__mux2_1
XFILLER_49_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4991_ clknet_leaf_1_wb_clk_i _0601_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[22\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3802__A0 _1710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3942_ _1879_ vssd1 vssd1 vccd1 vccd1 _0506_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__2605__A1 _0928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3873_ _1841_ vssd1 vssd1 vccd1 vccd1 _0475_ sky130_fd_sc_hd__clkbuf_1
X_2824_ _0921_ _1213_ vssd1 vssd1 vccd1 vccd1 _1214_ sky130_fd_sc_hd__or2_1
XANTENNA__2215__S _0668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_15_wb_clk_i_A clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__3835__A _1034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2755_ _0786_ _1144_ _0828_ vssd1 vssd1 vccd1 vccd1 _1145_ sky130_fd_sc_hd__a21o_1
X_2686_ _1074_ _1075_ _1076_ _0785_ _0793_ vssd1 vssd1 vccd1 vccd1 _1077_ sky130_fd_sc_hd__a221o_1
X_4425_ clknet_leaf_26_wb_clk_i _0024_ vssd1 vssd1 vccd1 vccd1 wbs_o_buff\[29\] sky130_fd_sc_hd__dfxtp_1
X_4356_ _2160_ vssd1 vssd1 vccd1 vccd1 _0639_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__2767__S1 _0813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3307_ _1515_ vssd1 vssd1 vccd1 vccd1 _0235_ sky130_fd_sc_hd__clkbuf_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4287_ _2122_ vssd1 vssd1 vccd1 vccd1 _0608_ sky130_fd_sc_hd__clkbuf_1
X_3238_ _1337_ _1430_ vssd1 vssd1 vccd1 vccd1 _1475_ sky130_fd_sc_hd__nor2_2
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3169_ _1368_ tms1x00.RAM\[124\]\[3\] _1431_ vssd1 vssd1 vccd1 vccd1 _1435_ sky130_fd_sc_hd__mux2_1
XANTENNA__4867__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2758__S1 _0813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5022__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2824__A _0921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output104_A net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3012__A1 _1334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2540_ _0822_ vssd1 vssd1 vccd1 vccd1 _0932_ sky130_fd_sc_hd__clkbuf_8
X_2471_ tms1x00.RAM\[28\]\[0\] tms1x00.RAM\[29\]\[0\] _0826_ vssd1 vssd1 vccd1 vccd1
+ _0864_ sky130_fd_sc_hd__mux2_1
X_4210_ _2073_ _2074_ vssd1 vssd1 vccd1 vccd1 _2075_ sky130_fd_sc_hd__nor2_1
X_4141_ tms1x00.ins_in\[5\] _1031_ _2011_ _2016_ vssd1 vssd1 vccd1 vccd1 _2017_ sky130_fd_sc_hd__a211o_1
XFILLER_68_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4072_ _0742_ tms1x00.A\[3\] vssd1 vssd1 vccd1 vccd1 _1967_ sky130_fd_sc_hd__and2b_1
XFILLER_37_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3023_ _1349_ vssd1 vssd1 vccd1 vccd1 _0117_ sky130_fd_sc_hd__clkbuf_1
XFILLER_37_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4974_ clknet_leaf_8_wb_clk_i _0584_ vssd1 vssd1 vccd1 vccd1 tms1x00.N\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_52_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3925_ _1258_ _1286_ vssd1 vssd1 vccd1 vccd1 _1870_ sky130_fd_sc_hd__nor2_2
XANTENNA__3549__B _1337_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2453__B _0845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3856_ _1819_ tms1x00.RAM\[81\]\[1\] _1830_ vssd1 vssd1 vccd1 vccd1 _1832_ sky130_fd_sc_hd__mux2_1
X_2807_ _0921_ _1192_ _1196_ _0806_ vssd1 vssd1 vccd1 vccd1 _1197_ sky130_fd_sc_hd__o211a_1
X_3787_ tms1x00.RAM\[7\]\[0\] _1772_ _1791_ vssd1 vssd1 vccd1 vccd1 _1792_ sky130_fd_sc_hd__mux2_1
X_2738_ _1128_ vssd1 vssd1 vccd1 vccd1 _1129_ sky130_fd_sc_hd__buf_4
X_2669_ _0948_ _1057_ _1059_ _0776_ vssd1 vssd1 vccd1 vccd1 _1060_ sky130_fd_sc_hd__o211a_1
X_4408_ clknet_leaf_28_wb_clk_i _0006_ vssd1 vssd1 vccd1 vccd1 wbs_o_buff\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_59_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4339_ _1251_ _1343_ vssd1 vssd1 vccd1 vccd1 _2151_ sky130_fd_sc_hd__or2_2
XFILLER_75_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2817__A1 _0940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5045__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input65_A wbs_dat_i[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2257__C valid vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4412__CLK clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2667__S0 _0799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3710_ _1237_ _1317_ vssd1 vssd1 vccd1 vccd1 _1747_ sky130_fd_sc_hd__nor2_2
XFILLER_41_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4690_ clknet_leaf_27_wb_clk_i _0304_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[43\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_3641_ _1129_ vssd1 vssd1 vccd1 vccd1 _1708_ sky130_fd_sc_hd__buf_2
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3572_ tms1x00.RAM\[5\]\[2\] _1576_ _1664_ vssd1 vssd1 vccd1 vccd1 _1667_ sky130_fd_sc_hd__mux2_1
X_2523_ _0915_ tms1x00.ram_addr_buff\[3\] tms1x00.ram_addr_buff\[2\] vssd1 vssd1 vccd1
+ vccd1 _0916_ sky130_fd_sc_hd__and3b_2
X_2454_ tms1x00.RAM\[124\]\[0\] tms1x00.RAM\[125\]\[0\] tms1x00.RAM\[126\]\[0\] tms1x00.RAM\[127\]\[0\]
+ _0815_ _0812_ vssd1 vssd1 vccd1 vccd1 _0847_ sky130_fd_sc_hd__mux4_1
XANTENNA__3832__B _1257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2385_ _0777_ vssd1 vssd1 vccd1 vccd1 _0778_ sky130_fd_sc_hd__buf_4
XFILLER_69_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4124_ _2002_ vssd1 vssd1 vccd1 vccd1 _0565_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5105__A net47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput1 io_in[5] vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__clkbuf_1
XFILLER_68_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4055_ _0733_ _1935_ vssd1 vssd1 vccd1 vccd1 _1954_ sky130_fd_sc_hd__nand2_1
X_3006_ tms1x00.RAM\[100\]\[0\] _1324_ _1338_ vssd1 vssd1 vccd1 vccd1 _1339_ sky130_fd_sc_hd__mux2_1
XFILLER_24_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4905__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4957_ clknet_leaf_9_wb_clk_i _0567_ vssd1 vssd1 vccd1 vccd1 tms1x00.P\[0\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__2658__S0 _0799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3908_ _1816_ tms1x00.RAM\[93\]\[0\] _1860_ vssd1 vssd1 vccd1 vccd1 _1861_ sky130_fd_sc_hd__mux2_1
X_4888_ clknet_leaf_22_wb_clk_i _0502_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[91\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_3839_ _1821_ tms1x00.RAM\[83\]\[2\] _1817_ vssd1 vssd1 vccd1 vccd1 _1822_ sky130_fd_sc_hd__mux2_1
XFILLER_20_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2735__B1 _1104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4435__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3999__C1 _1901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2374__A net76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3189__B _1430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4585__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3215__A1 _1461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4928__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4811_ clknet_leaf_24_wb_clk_i _0425_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[75\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_15_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4742_ clknet_leaf_26_wb_clk_i _0356_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[57\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_4673_ clknet_leaf_10_wb_clk_i _0045_ vssd1 vssd1 vccd1 vccd1 _0038_ sky130_fd_sc_hd__dfxtp_2
XANTENNA__2731__B _1121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3624_ _1697_ vssd1 vssd1 vccd1 vccd1 _0370_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__3319__S _1519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4004__A _0732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2812__S0 _0816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3555_ _1657_ vssd1 vssd1 vccd1 vccd1 _0341_ sky130_fd_sc_hd__clkbuf_1
X_3486_ _1273_ _1283_ vssd1 vssd1 vccd1 vccd1 _1619_ sky130_fd_sc_hd__or2_2
X_2506_ tms1x00.RAM\[48\]\[0\] tms1x00.RAM\[49\]\[0\] tms1x00.RAM\[50\]\[0\] tms1x00.RAM\[51\]\[0\]
+ _0815_ _0812_ vssd1 vssd1 vccd1 vccd1 _0899_ sky130_fd_sc_hd__mux4_1
X_2437_ _0777_ vssd1 vssd1 vccd1 vccd1 _0830_ sky130_fd_sc_hd__buf_6
XFILLER_69_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2368_ _0757_ _0758_ _0761_ _0762_ vssd1 vssd1 vccd1 vccd1 _0763_ sky130_fd_sc_hd__and4b_2
XFILLER_56_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3693__A1 _1669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4107_ _1990_ vssd1 vssd1 vccd1 vccd1 _0560_ sky130_fd_sc_hd__clkbuf_1
XFILLER_38_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2299_ _0709_ vssd1 vssd1 vccd1 vccd1 _0023_ sky130_fd_sc_hd__clkbuf_1
X_4038_ _0754_ _0730_ _1918_ vssd1 vssd1 vccd1 vccd1 _1942_ sky130_fd_sc_hd__or3b_1
XFILLER_37_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2653__C1 _0776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3737__B _1409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2708__B1 _0850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2369__A _0763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input28_A ram_val[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2832__A _0747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2947__A0 _1035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3647__B _1409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output96_A net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3340_ _1534_ vssd1 vssd1 vccd1 vccd1 _0249_ sky130_fd_sc_hd__clkbuf_1
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3271_ _1495_ vssd1 vssd1 vccd1 vccd1 _0219_ sky130_fd_sc_hd__clkbuf_1
X_5010_ clknet_leaf_12_wb_clk_i _0620_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[12\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4750__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2222_ _0678_ vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__clkbuf_1
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2635__C1 _0804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3838__A _1129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2938__A0 _1035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2986_ _0910_ vssd1 vssd1 vccd1 vccd1 _1323_ sky130_fd_sc_hd__clkbuf_4
XFILLER_21_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4725_ clknet_leaf_28_wb_clk_i _0339_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[52\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_4656_ clknet_leaf_6_wb_clk_i _0277_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[33\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_4587_ clknet_leaf_0_wb_clk_i _0208_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[116\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_3607_ _1284_ _1310_ vssd1 vssd1 vccd1 vccd1 _1688_ sky130_fd_sc_hd__nor2_2
X_3538_ tms1x00.RAM\[54\]\[3\] _1578_ _1644_ vssd1 vssd1 vccd1 vccd1 _1648_ sky130_fd_sc_hd__mux2_1
XANTENNA__2511__D_N tms1x00.ins_in\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3469_ tms1x00.RAM\[43\]\[0\] _1571_ _1609_ vssd1 vssd1 vccd1 vccd1 _1610_ sky130_fd_sc_hd__mux2_1
XFILLER_69_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_8_wb_clk_i clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_38_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2641__A2 _1030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2652__A _0819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4623__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4146__A2 _2007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2798__S _0778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2827__A _0783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2840_ _1227_ _1228_ vssd1 vssd1 vccd1 vccd1 _1229_ sky130_fd_sc_hd__or2_4
XFILLER_31_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2771_ tms1x00.RAM\[100\]\[3\] tms1x00.RAM\[101\]\[3\] tms1x00.RAM\[102\]\[3\] tms1x00.RAM\[103\]\[3\]
+ _0873_ _0977_ vssd1 vssd1 vccd1 vccd1 _1161_ sky130_fd_sc_hd__mux4_1
X_4510_ clknet_leaf_15_wb_clk_i _0131_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[95\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2491__S1 _0779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4441_ clknet_leaf_24_wb_clk_i _0062_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[69\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3896__A1 _1779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4372_ _2169_ vssd1 vssd1 vccd1 vccd1 _0646_ sky130_fd_sc_hd__clkbuf_1
X_3323_ tms1x00.ram_addr_buff\[4\] tms1x00.ram_addr_buff\[6\] tms1x00.ram_addr_buff\[5\]
+ vssd1 vssd1 vccd1 vccd1 _1524_ sky130_fd_sc_hd__or3b_2
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3254_ _1368_ tms1x00.RAM\[115\]\[3\] _1480_ vssd1 vssd1 vccd1 vccd1 _1484_ sky130_fd_sc_hd__mux2_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2205_ net16 wbs_o_buff\[11\] _0668_ vssd1 vssd1 vccd1 vccd1 _0670_ sky130_fd_sc_hd__mux2_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3185_ tms1x00.RAM\[122\]\[2\] _1331_ _1441_ vssd1 vssd1 vccd1 vccd1 _1444_ sky130_fd_sc_hd__mux2_1
XFILLER_27_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4646__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3820__A1 _1779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2623__A2 _1014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3287__B _1303_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2969_ tms1x00.RAM\[103\]\[1\] _1243_ _1311_ vssd1 vssd1 vccd1 vccd1 _1313_ sky130_fd_sc_hd__mux2_1
X_4708_ clknet_leaf_3_wb_clk_i _0322_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[48\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4639_ clknet_leaf_0_wb_clk_i _0260_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[37\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3887__A1 _1779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2311__A1 tms1x00.wb_step vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2473__S1 _0800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3925__B _1286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3878__A1 _1779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4669__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4990_ clknet_leaf_0_wb_clk_i _0600_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[22\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3388__A _1273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3941_ tms1x00.RAM\[90\]\[3\] _1333_ _1875_ vssd1 vssd1 vccd1 vccd1 _1879_ sky130_fd_sc_hd__mux2_1
XFILLER_32_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3872_ tms1x00.RAM\[8\]\[0\] _1772_ _1840_ vssd1 vssd1 vccd1 vccd1 _1841_ sky130_fd_sc_hd__mux2_1
X_2823_ tms1x00.RAM\[48\]\[3\] tms1x00.RAM\[49\]\[3\] tms1x00.RAM\[50\]\[3\] tms1x00.RAM\[51\]\[3\]
+ _0816_ _0977_ vssd1 vssd1 vccd1 vccd1 _1213_ sky130_fd_sc_hd__mux4_2
X_2754_ tms1x00.RAM\[68\]\[3\] tms1x00.RAM\[69\]\[3\] _0826_ vssd1 vssd1 vccd1 vccd1
+ _1144_ sky130_fd_sc_hd__mux2_1
X_2685_ tms1x00.RAM\[12\]\[2\] tms1x00.RAM\[13\]\[2\] _0823_ vssd1 vssd1 vccd1 vccd1
+ _1076_ sky130_fd_sc_hd__mux2_1
X_4424_ clknet_leaf_26_wb_clk_i _0023_ vssd1 vssd1 vccd1 vccd1 wbs_o_buff\[28\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__3869__A1 _1779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4355_ _1247_ tms1x00.RAM\[13\]\[3\] _2156_ vssd1 vssd1 vccd1 vccd1 _2160_ sky130_fd_sc_hd__mux2_1
XFILLER_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3306_ tms1x00.RAM\[27\]\[0\] _1456_ _1514_ vssd1 vssd1 vccd1 vccd1 _1515_ sky130_fd_sc_hd__mux2_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4286_ tms1x00.RAM\[21\]\[0\] _1323_ _2121_ vssd1 vssd1 vccd1 vccd1 _2122_ sky130_fd_sc_hd__mux2_1
XFILLER_55_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3237_ _1474_ vssd1 vssd1 vccd1 vccd1 _0206_ sky130_fd_sc_hd__clkbuf_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3168_ _1434_ vssd1 vssd1 vccd1 vccd1 _0177_ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_0_wb_clk_i_A clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_82_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3099_ _1366_ tms1x00.RAM\[111\]\[2\] _1391_ vssd1 vssd1 vccd1 vccd1 _1394_ sky130_fd_sc_hd__mux2_1
XFILLER_55_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4811__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input10_A oram_value[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3796__A0 _1703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2824__B _1213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2470_ _0822_ _0862_ vssd1 vssd1 vccd1 vccd1 _0863_ sky130_fd_sc_hd__and2_1
XFILLER_79_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4140_ _0743_ tms1x00.K_latch\[1\] _1956_ _2012_ tms1x00.Y\[1\] vssd1 vssd1 vccd1
+ vccd1 _2016_ sky130_fd_sc_hd__a32o_1
XFILLER_69_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4071_ _1958_ _1964_ _1965_ _1966_ vssd1 vssd1 vccd1 vccd1 _0548_ sky130_fd_sc_hd__o211a_1
XFILLER_49_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3022_ _1130_ tms1x00.RAM\[0\]\[2\] _1346_ vssd1 vssd1 vccd1 vccd1 _1349_ sky130_fd_sc_hd__mux2_1
XANTENNA__2287__B1 _0704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4973_ clknet_leaf_9_wb_clk_i _0583_ vssd1 vssd1 vccd1 vccd1 tms1x00.X\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_24_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3924_ _1869_ vssd1 vssd1 vccd1 vccd1 _0498_ sky130_fd_sc_hd__clkbuf_1
XFILLER_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3855_ _1831_ vssd1 vssd1 vccd1 vccd1 _0467_ sky130_fd_sc_hd__clkbuf_1
X_2806_ _1193_ _1194_ _1195_ _0786_ _0794_ vssd1 vssd1 vccd1 vccd1 _1196_ sky130_fd_sc_hd__a221o_1
X_3786_ _1310_ _1344_ vssd1 vssd1 vccd1 vccd1 _1791_ sky130_fd_sc_hd__nor2_2
X_2737_ _0771_ _1126_ _1127_ _0909_ tms1x00.A\[2\] vssd1 vssd1 vccd1 vccd1 _1128_
+ sky130_fd_sc_hd__a32o_1
XANTENNA__2211__A0 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_22_wb_clk_i clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_2668_ _0819_ _1058_ vssd1 vssd1 vccd1 vccd1 _1059_ sky130_fd_sc_hd__or2_1
XANTENNA__2762__B2 _0786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4834__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4407_ clknet_leaf_29_wb_clk_i _0005_ vssd1 vssd1 vccd1 vccd1 wbs_o_buff\[11\] sky130_fd_sc_hd__dfxtp_1
X_2599_ tms1x00.RAM\[24\]\[1\] tms1x00.RAM\[25\]\[1\] tms1x00.RAM\[26\]\[1\] tms1x00.RAM\[27\]\[1\]
+ _0945_ _0791_ vssd1 vssd1 vccd1 vccd1 _0991_ sky130_fd_sc_hd__mux4_2
XFILLER_59_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4338_ _2150_ vssd1 vssd1 vccd1 vccd1 _0631_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_input2_A io_in[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4269_ _2112_ vssd1 vssd1 vccd1 vccd1 _0600_ sky130_fd_sc_hd__clkbuf_1
XFILLER_75_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4984__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2278__B1 _0703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2817__A2 _1204_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3520__S _1634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3778__A0 _1703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3756__A _1237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input58_A wbs_cyc_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2835__A _1224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4707__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2667__S1 _0800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2441__B1 _0821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3640_ _1707_ vssd1 vssd1 vccd1 vccd1 _0376_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__2570__A _0940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4261__S _2106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3571_ _1666_ vssd1 vssd1 vccd1 vccd1 _0348_ sky130_fd_sc_hd__clkbuf_1
X_2522_ _0905_ _0771_ vssd1 vssd1 vccd1 vccd1 _0915_ sky130_fd_sc_hd__and2_1
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3941__A0 tms1x00.RAM\[90\]\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2453_ _0797_ _0845_ vssd1 vssd1 vccd1 vccd1 _0846_ sky130_fd_sc_hd__or2_1
X_2384_ _0035_ vssd1 vssd1 vccd1 vccd1 _0777_ sky130_fd_sc_hd__buf_6
XFILLER_68_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4123_ _0738_ _2001_ vssd1 vssd1 vccd1 vccd1 _2002_ sky130_fd_sc_hd__or2_1
Xinput2 io_in[6] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_1
XFILLER_68_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4054_ net91 _1952_ _1953_ _1931_ vssd1 vssd1 vccd1 vccd1 _0544_ sky130_fd_sc_hd__o211a_1
XFILLER_56_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3005_ _0914_ _1337_ vssd1 vssd1 vccd1 vccd1 _1338_ sky130_fd_sc_hd__nor2_2
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4956_ clknet_leaf_6_wb_clk_i _0566_ vssd1 vssd1 vccd1 vccd1 tms1x00.PA\[3\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__2658__S1 _0800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3907_ _0917_ _1257_ vssd1 vssd1 vccd1 vccd1 _1860_ sky130_fd_sc_hd__or2_2
XANTENNA__3576__A _0911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4887_ clknet_leaf_22_wb_clk_i _0501_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[91\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2480__A _0815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3838_ _1129_ vssd1 vssd1 vccd1 vccd1 _1821_ sky130_fd_sc_hd__clkbuf_4
XFILLER_20_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3769_ tms1x00.RAM\[73\]\[0\] _1772_ _1781_ vssd1 vssd1 vccd1 vccd1 _1782_ sky130_fd_sc_hd__mux2_1
XANTENNA__5012__CLK clknet_leaf_20_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2639__B _0748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2374__B net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3486__A _1273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3923__A0 _1823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4810_ clknet_leaf_24_wb_clk_i _0424_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[75\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4741_ clknet_leaf_26_wb_clk_i _0355_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[57\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_15_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4672_ clknet_leaf_2_wb_clk_i _0044_ vssd1 vssd1 vccd1 vccd1 _0037_ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2504__S _0826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3623_ _1592_ tms1x00.RAM\[63\]\[3\] _1693_ vssd1 vssd1 vccd1 vccd1 _1697_ sky130_fd_sc_hd__mux2_1
XANTENNA__4004__B _0730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3914__A0 _1823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2717__B2 _0818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2812__S1 _0927_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3554_ tms1x00.RAM\[52\]\[2\] _1576_ _1654_ vssd1 vssd1 vccd1 vccd1 _1657_ sky130_fd_sc_hd__mux2_1
X_2505_ _0895_ _0896_ _0897_ _0785_ _0828_ vssd1 vssd1 vccd1 vccd1 _0898_ sky130_fd_sc_hd__a221o_1
X_3485_ _1618_ vssd1 vssd1 vccd1 vccd1 _0310_ sky130_fd_sc_hd__clkbuf_1
X_2436_ _0786_ _0827_ _0828_ vssd1 vssd1 vccd1 vccd1 _0829_ sky130_fd_sc_hd__a21o_1
XFILLER_69_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2367_ tms1x00.ins_in\[4\] vssd1 vssd1 vccd1 vccd1 _0762_ sky130_fd_sc_hd__clkinv_2
X_4106_ net103 _1989_ vssd1 vssd1 vccd1 vccd1 _1990_ sky130_fd_sc_hd__or2_1
XFILLER_38_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2298_ wbs_o_buff\[28\] _0704_ vssd1 vssd1 vccd1 vccd1 _0709_ sky130_fd_sc_hd__and2_1
X_4037_ _0753_ _1940_ _1941_ _1931_ vssd1 vssd1 vccd1 vccd1 _0539_ sky130_fd_sc_hd__o211a_1
XFILLER_56_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4939_ clknet_leaf_7_wb_clk_i _0549_ vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__dfxtp_2
XANTENNA__2500__S0 _0777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2956__A1 _1235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3905__A0 _1823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2708__A1 _0830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4552__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2385__A _0777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2644__A0 _1035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2832__B _0748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output89_A net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3270_ _1485_ tms1x00.RAM\[125\]\[0\] _1494_ vssd1 vssd1 vccd1 vccd1 _1495_ sky130_fd_sc_hd__mux2_1
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2221_ net24 wbs_o_buff\[19\] _0668_ vssd1 vssd1 vccd1 vccd1 _0678_ sky130_fd_sc_hd__mux2_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_34_wb_clk_i_A clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_46_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2730__S0 _0823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3060__A0 _1364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2938__A1 tms1x00.RAM\[49\]\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4724_ clknet_leaf_28_wb_clk_i _0338_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[53\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2985_ _1322_ vssd1 vssd1 vccd1 vccd1 _0106_ sky130_fd_sc_hd__clkbuf_1
X_4655_ clknet_leaf_10_wb_clk_i _0276_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[33\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4425__CLK clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4586_ clknet_leaf_1_wb_clk_i _0207_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[116\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput60 wbs_dat_i[10] vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__clkbuf_1
X_3606_ _1687_ vssd1 vssd1 vccd1 vccd1 _0362_ sky130_fd_sc_hd__clkbuf_1
X_3537_ _1647_ vssd1 vssd1 vccd1 vccd1 _0333_ sky130_fd_sc_hd__clkbuf_1
XFILLER_1_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4575__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3468_ _1286_ _1525_ vssd1 vssd1 vccd1 vccd1 _1609_ sky130_fd_sc_hd__nor2_2
XFILLER_76_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3399_ _1567_ vssd1 vssd1 vccd1 vccd1 _0275_ sky130_fd_sc_hd__clkbuf_1
X_2419_ _0036_ vssd1 vssd1 vccd1 vccd1 _0812_ sky130_fd_sc_hd__buf_6
XANTENNA__2874__A0 _1035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2721__S0 _0823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2652__B _1042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4379__A0 tms1x00.PC\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2929__A1 _1243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4918__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input40_A ram_val[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4067__C1 _1931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4448__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3042__A0 _1225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2770_ tms1x00.RAM\[96\]\[3\] tms1x00.RAM\[97\]\[3\] tms1x00.RAM\[98\]\[3\] tms1x00.RAM\[99\]\[3\]
+ _0931_ _0932_ vssd1 vssd1 vccd1 vccd1 _1160_ sky130_fd_sc_hd__mux4_2
XFILLER_8_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3674__A _1236_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4440_ clknet_leaf_22_wb_clk_i _0061_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[69\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_4371_ tms1x00.RAM\[9\]\[2\] _1330_ _2166_ vssd1 vssd1 vccd1 vccd1 _2169_ sky130_fd_sc_hd__mux2_1
X_3322_ _1523_ vssd1 vssd1 vccd1 vccd1 _0242_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3253_ _1483_ vssd1 vssd1 vccd1 vccd1 _0213_ sky130_fd_sc_hd__clkbuf_1
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2204_ _0669_ vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__clkbuf_1
X_3184_ _1443_ vssd1 vssd1 vccd1 vccd1 _0184_ sky130_fd_sc_hd__clkbuf_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2608__B1 _0776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2753__A _0822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3033__A0 _1225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2968_ _1312_ vssd1 vssd1 vccd1 vccd1 _0099_ sky130_fd_sc_hd__clkbuf_1
X_4707_ clknet_leaf_3_wb_clk_i _0321_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[48\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3584__A1 _1674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2899_ _1270_ vssd1 vssd1 vccd1 vccd1 _0072_ sky130_fd_sc_hd__clkbuf_1
X_4638_ clknet_leaf_1_wb_clk_i _0259_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[37\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4569_ clknet_leaf_33_wb_clk_i _0190_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[121\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_77_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3523__S _1639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3272__A0 _1488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3759__A _1034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3024__A0 _1225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4740__CLK clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4191__C_N _0747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapped_tms1x00_190 vssd1 vssd1 vccd1 vccd1 io_oeb[0] wrapped_tms1x00_190/LO sky130_fd_sc_hd__conb_1
XFILLER_5_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2602__S _0924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2783__C1 _0806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3940_ _1878_ vssd1 vssd1 vccd1 vccd1 _0505_ sky130_fd_sc_hd__clkbuf_1
XFILLER_17_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2292__B _0704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3871_ _1303_ _1344_ vssd1 vssd1 vccd1 vccd1 _1840_ sky130_fd_sc_hd__nor2_2
XFILLER_31_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2822_ _1209_ _1210_ _1211_ _0787_ _0996_ vssd1 vssd1 vccd1 vccd1 _1212_ sky130_fd_sc_hd__a221o_1
X_2753_ _0822_ _1142_ vssd1 vssd1 vccd1 vccd1 _1143_ sky130_fd_sc_hd__and2_1
XFILLER_8_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2684_ _0788_ tms1x00.RAM\[14\]\[2\] _0812_ vssd1 vssd1 vccd1 vccd1 _1075_ sky130_fd_sc_hd__o21a_1
XANTENNA__4012__B _0763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4423_ clknet_leaf_26_wb_clk_i _0022_ vssd1 vssd1 vccd1 vccd1 wbs_o_buff\[27\] sky130_fd_sc_hd__dfxtp_1
X_4354_ _2159_ vssd1 vssd1 vccd1 vccd1 _0638_ sky130_fd_sc_hd__clkbuf_1
X_3305_ _1250_ _1286_ vssd1 vssd1 vccd1 vccd1 _1514_ sky130_fd_sc_hd__nor2_2
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4285_ _1240_ _1250_ vssd1 vssd1 vccd1 vccd1 _2121_ sky130_fd_sc_hd__nor2_2
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3236_ tms1x00.RAM\[117\]\[3\] _1463_ _1470_ vssd1 vssd1 vccd1 vccd1 _1474_ sky130_fd_sc_hd__mux2_1
XANTENNA__2829__B1 _0920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3167_ _1366_ tms1x00.RAM\[124\]\[2\] _1431_ vssd1 vssd1 vccd1 vccd1 _1434_ sky130_fd_sc_hd__mux2_1
XFILLER_27_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3098_ _1393_ vssd1 vssd1 vccd1 vccd1 _0148_ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3254__A0 _1368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4763__CLK clknet_leaf_20_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2765__C1 _0773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3518__S _1634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2377__B _0768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3493__A0 _1592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2508__C1 _0804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output71_A net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_916 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4636__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3720__A1 _1669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4259__S _2106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4070_ _0718_ vssd1 vssd1 vccd1 vccd1 _1966_ sky130_fd_sc_hd__clkbuf_4
XFILLER_49_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3021_ _1348_ vssd1 vssd1 vccd1 vccd1 _0116_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__2287__A1 net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4972_ clknet_leaf_9_wb_clk_i _0582_ vssd1 vssd1 vccd1 vccd1 tms1x00.X\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_52_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3923_ _1823_ tms1x00.RAM\[92\]\[3\] _1865_ vssd1 vssd1 vccd1 vccd1 _1869_ sky130_fd_sc_hd__mux2_1
XFILLER_32_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3787__A1 _1772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3854_ _1816_ tms1x00.RAM\[81\]\[0\] _1830_ vssd1 vssd1 vccd1 vccd1 _1831_ sky130_fd_sc_hd__mux2_1
X_2805_ tms1x00.RAM\[12\]\[3\] tms1x00.RAM\[13\]\[3\] _0778_ vssd1 vssd1 vccd1 vccd1
+ _1195_ sky130_fd_sc_hd__mux2_1
XFILLER_20_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3785_ _1790_ vssd1 vssd1 vccd1 vccd1 _0438_ sky130_fd_sc_hd__clkbuf_1
X_2736_ _0748_ _0747_ vssd1 vssd1 vccd1 vccd1 _1127_ sky130_fd_sc_hd__or2b_1
X_2667_ tms1x00.RAM\[20\]\[2\] tms1x00.RAM\[21\]\[2\] tms1x00.RAM\[22\]\[2\] tms1x00.RAM\[23\]\[2\]
+ _0799_ _0800_ vssd1 vssd1 vccd1 vccd1 _1058_ sky130_fd_sc_hd__mux4_2
XANTENNA__3862__A _1258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4406_ clknet_leaf_28_wb_clk_i _0004_ vssd1 vssd1 vccd1 vccd1 wbs_o_buff\[10\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__2514__A2 _0858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2598_ _0932_ _0989_ _0819_ vssd1 vssd1 vccd1 vccd1 _0990_ sky130_fd_sc_hd__a21o_1
XANTENNA__3711__A1 _1669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4337_ _1247_ tms1x00.RAM\[15\]\[3\] _2146_ vssd1 vssd1 vccd1 vccd1 _2150_ sky130_fd_sc_hd__mux2_1
XFILLER_59_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4268_ tms1x00.RAM\[22\]\[0\] _1323_ _2111_ vssd1 vssd1 vccd1 vccd1 _2112_ sky130_fd_sc_hd__mux2_1
XFILLER_55_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2278__A1 net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3219_ _1464_ vssd1 vssd1 vccd1 vccd1 _0198_ sky130_fd_sc_hd__clkbuf_1
X_4199_ _2065_ vssd1 vssd1 vccd1 vccd1 _0577_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2803__B_N _0840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_668 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4509__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3756__B _1403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3950__A1 _1333_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4659__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3702__A1 _1669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3466__A0 _1592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2269__A1 net75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3769__A1 _1772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2441__A1 _0806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3570_ tms1x00.RAM\[5\]\[1\] _1574_ _1664_ vssd1 vssd1 vccd1 vccd1 _1666_ sky130_fd_sc_hd__mux2_1
X_2521_ _0913_ vssd1 vssd1 vccd1 vccd1 _0914_ sky130_fd_sc_hd__clkbuf_8
XFILLER_6_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3941__A1 _1333_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2452_ tms1x00.RAM\[120\]\[0\] tms1x00.RAM\[121\]\[0\] tms1x00.RAM\[122\]\[0\] tms1x00.RAM\[123\]\[0\]
+ _0815_ _0812_ vssd1 vssd1 vccd1 vccd1 _0845_ sky130_fd_sc_hd__mux4_1
X_2383_ _0775_ vssd1 vssd1 vccd1 vccd1 _0776_ sky130_fd_sc_hd__clkbuf_4
XFILLER_68_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4122_ tms1x00.PB\[2\] tms1x00.PA\[2\] _1996_ vssd1 vssd1 vccd1 vccd1 _2001_ sky130_fd_sc_hd__mux2_1
X_4053_ _0755_ _0752_ _1932_ vssd1 vssd1 vccd1 vccd1 _1953_ sky130_fd_sc_hd__or3_1
XFILLER_56_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3457__A0 _1592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput3 io_in[7] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_1
X_3004_ _1336_ vssd1 vssd1 vccd1 vccd1 _1337_ sky130_fd_sc_hd__clkbuf_8
XFILLER_64_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4955_ clknet_leaf_6_wb_clk_i _0565_ vssd1 vssd1 vccd1 vccd1 tms1x00.PA\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_40_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3906_ _1859_ vssd1 vssd1 vccd1 vccd1 _0490_ sky130_fd_sc_hd__clkbuf_1
XFILLER_60_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4886_ clknet_leaf_21_wb_clk_i _0500_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[91\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_3837_ _1820_ vssd1 vssd1 vccd1 vccd1 _0460_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4801__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2196__A0 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3768_ _1237_ _1261_ vssd1 vssd1 vccd1 vccd1 _1781_ sky130_fd_sc_hd__nor2_2
X_2719_ _0921_ _1109_ vssd1 vssd1 vccd1 vccd1 _1110_ sky130_fd_sc_hd__or2_1
XANTENNA__3932__A1 _1779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2700__S _0788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3699_ tms1x00.RAM\[72\]\[3\] _1676_ _1737_ vssd1 vssd1 vccd1 vccd1 _1741_ sky130_fd_sc_hd__mux2_1
XANTENNA__4951__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2374__C tms1x00.ins_in\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2671__A _0932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3486__B _1283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2610__S _0975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3439__A0 _1592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_24_wb_clk_i_A clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_19_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4272__S _2111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4740_ clknet_leaf_26_wb_clk_i _0354_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[58\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_4671_ clknet_leaf_11_wb_clk_i _0043_ vssd1 vssd1 vccd1 vccd1 _0036_ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3622_ _1696_ vssd1 vssd1 vccd1 vccd1 _0369_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4004__C _0752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4974__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3553_ _1656_ vssd1 vssd1 vccd1 vccd1 _0340_ sky130_fd_sc_hd__clkbuf_1
X_3484_ tms1x00.RAM\[42\]\[3\] _1578_ _1614_ vssd1 vssd1 vccd1 vccd1 _1618_ sky130_fd_sc_hd__mux2_1
X_2504_ tms1x00.RAM\[52\]\[0\] tms1x00.RAM\[53\]\[0\] _0826_ vssd1 vssd1 vccd1 vccd1
+ _0897_ sky130_fd_sc_hd__mux2_1
X_2435_ _0793_ vssd1 vssd1 vccd1 vccd1 _0828_ sky130_fd_sc_hd__clkbuf_4
X_2366_ _0760_ _0745_ vssd1 vssd1 vccd1 vccd1 _0761_ sky130_fd_sc_hd__nor2_1
X_4105_ tms1x00.PA\[1\] _1973_ _1987_ tms1x00.PB\[1\] vssd1 vssd1 vccd1 vccd1 _1989_
+ sky130_fd_sc_hd__a22o_1
XFILLER_29_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2297_ _0708_ vssd1 vssd1 vccd1 vccd1 _0022_ sky130_fd_sc_hd__clkbuf_1
X_4036_ _0733_ _0739_ _0764_ _1915_ net86 vssd1 vssd1 vccd1 vccd1 _1941_ sky130_fd_sc_hd__a41o_1
XFILLER_71_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2653__A1 _0948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4061__A_N _0742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4938_ clknet_leaf_7_wb_clk_i _0548_ vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__dfxtp_2
XFILLER_40_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4869_ clknet_leaf_23_wb_clk_i _0483_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[87\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2500__S1 _0779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2892__A1 _1247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4847__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4997__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2220_ _0677_ vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__clkbuf_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_527 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2730__S1 _0850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5002__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2984_ tms1x00.RAM\[102\]\[3\] _1247_ _1318_ vssd1 vssd1 vccd1 vccd1 _1322_ sky130_fd_sc_hd__mux2_1
X_4723_ clknet_leaf_29_wb_clk_i _0337_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[53\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2494__S0 _0799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4654_ clknet_leaf_6_wb_clk_i _0275_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[33\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3899__A0 _1816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4585_ clknet_leaf_3_wb_clk_i _0206_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[117\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput50 wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__clkbuf_1
Xinput61 wbs_dat_i[11] vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__clkbuf_1
X_3605_ tms1x00.RAM\[56\]\[3\] _1676_ _1683_ vssd1 vssd1 vccd1 vccd1 _1687_ sky130_fd_sc_hd__mux2_1
XANTENNA__2250__S net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4031__A _0718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3536_ tms1x00.RAM\[54\]\[2\] _1576_ _1644_ vssd1 vssd1 vccd1 vccd1 _1647_ sky130_fd_sc_hd__mux2_1
X_3467_ _1608_ vssd1 vssd1 vccd1 vccd1 _0302_ sky130_fd_sc_hd__clkbuf_1
X_3398_ _1485_ tms1x00.RAM\[33\]\[0\] _1566_ vssd1 vssd1 vccd1 vccd1 _1567_ sky130_fd_sc_hd__mux2_1
XANTENNA__2323__A0 tms1x00.Y\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2418_ tms1x00.RAM\[79\]\[0\] _0789_ vssd1 vssd1 vccd1 vccd1 _0811_ sky130_fd_sc_hd__or2b_1
X_2349_ _0743_ tms1x00.ins_in\[2\] vssd1 vssd1 vccd1 vccd1 _0744_ sky130_fd_sc_hd__nand2_1
XFILLER_45_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4019_ tms1x00.Y\[2\] _1915_ vssd1 vssd1 vccd1 vccd1 _1928_ sky130_fd_sc_hd__nand2_1
XFILLER_26_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2721__S1 _0850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4206__A _0766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4379__A1 net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2562__B1 _0953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2396__A _0788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input33_A ram_val[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5025__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3290__A1 _1459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2335__S _0726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2476__S0 _0808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3674__B _1251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4370_ _2168_ vssd1 vssd1 vccd1 vccd1 _0645_ sky130_fd_sc_hd__clkbuf_1
X_3321_ tms1x00.RAM\[26\]\[3\] _1463_ _1519_ vssd1 vssd1 vccd1 vccd1 _1523_ sky130_fd_sc_hd__mux2_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3252_ _1366_ tms1x00.RAM\[115\]\[2\] _1480_ vssd1 vssd1 vccd1 vccd1 _1483_ sky130_fd_sc_hd__mux2_1
XFILLER_39_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2203_ net15 wbs_o_buff\[10\] _0668_ vssd1 vssd1 vccd1 vccd1 _0669_ sky130_fd_sc_hd__mux2_1
X_3183_ tms1x00.RAM\[122\]\[1\] _1328_ _1441_ vssd1 vssd1 vccd1 vccd1 _1443_ sky130_fd_sc_hd__mux2_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3805__A0 _1703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2608__A1 _0948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_16_wb_clk_i clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__3281__A1 _1459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4026__A _0732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2967_ tms1x00.RAM\[103\]\[0\] _1235_ _1311_ vssd1 vssd1 vccd1 vccd1 _1312_ sky130_fd_sc_hd__mux2_1
XANTENNA__2467__S0 _0830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2898_ _1035_ tms1x00.RAM\[79\]\[1\] _1268_ vssd1 vssd1 vccd1 vccd1 _1270_ sky130_fd_sc_hd__mux2_1
X_4706_ clknet_leaf_3_wb_clk_i _0320_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[48\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4542__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4637_ clknet_leaf_3_wb_clk_i _0258_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[2\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4568_ clknet_leaf_32_wb_clk_i _0189_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[121\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_4499_ clknet_leaf_15_wb_clk_i _0120_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[98\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_3519_ _1637_ vssd1 vssd1 vccd1 vccd1 _0325_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4692__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4297__A0 _1819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2944__A _1229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwrapped_tms1x00_180 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_180/HI io_out[3] sky130_fd_sc_hd__conb_1
Xwrapped_tms1x00_191 vssd1 vssd1 vccd1 vccd1 io_oeb[1] wrapped_tms1x00_191/LO sky130_fd_sc_hd__conb_1
XANTENNA__3980__C1 _1901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3015__A _1343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3870_ _1839_ vssd1 vssd1 vccd1 vccd1 _0474_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__2449__S0 _0815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2821_ tms1x00.RAM\[52\]\[3\] tms1x00.RAM\[53\]\[3\] _0975_ vssd1 vssd1 vccd1 vccd1
+ _1211_ sky130_fd_sc_hd__mux2_1
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2752_ tms1x00.RAM\[70\]\[3\] tms1x00.RAM\[71\]\[3\] _0823_ vssd1 vssd1 vccd1 vccd1
+ _1142_ sky130_fd_sc_hd__mux2_1
X_2683_ tms1x00.RAM\[15\]\[2\] _0788_ vssd1 vssd1 vccd1 vccd1 _1074_ sky130_fd_sc_hd__or2b_1
X_4422_ clknet_leaf_27_wb_clk_i _0021_ vssd1 vssd1 vccd1 vccd1 wbs_o_buff\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_8_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2526__A0 _0912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4353_ _1245_ tms1x00.RAM\[13\]\[2\] _2156_ vssd1 vssd1 vccd1 vccd1 _2159_ sky130_fd_sc_hd__mux2_1
XANTENNA__4279__A0 _1819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3304_ _1513_ vssd1 vssd1 vccd1 vccd1 _0234_ sky130_fd_sc_hd__clkbuf_1
X_4284_ _2120_ vssd1 vssd1 vccd1 vccd1 _0607_ sky130_fd_sc_hd__clkbuf_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3235_ _1473_ vssd1 vssd1 vccd1 vccd1 _0205_ sky130_fd_sc_hd__clkbuf_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2829__A1 _0944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3166_ _1433_ vssd1 vssd1 vccd1 vccd1 _0176_ sky130_fd_sc_hd__clkbuf_1
XFILLER_54_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3097_ _1364_ tms1x00.RAM\[111\]\[1\] _1391_ vssd1 vssd1 vccd1 vccd1 _1393_ sky130_fd_sc_hd__mux2_1
XFILLER_54_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2764__A _0821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4908__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3999_ _1909_ _1912_ _1913_ _1901_ vssd1 vssd1 vccd1 vccd1 _0529_ sky130_fd_sc_hd__o211a_1
XFILLER_50_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3006__A1 _1324_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4438__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4588__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3245__A1 _1463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_928 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3020_ _1035_ tms1x00.RAM\[0\]\[1\] _1346_ vssd1 vssd1 vccd1 vccd1 _1348_ sky130_fd_sc_hd__mux2_1
XANTENNA__2287__A2 _0697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3484__A1 _1578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4971_ clknet_leaf_9_wb_clk_i _0581_ vssd1 vssd1 vccd1 vccd1 tms1x00.X\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3236__A1 _1463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4007__C _0763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3922_ _1868_ vssd1 vssd1 vccd1 vccd1 _0497_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3853_ _1251_ _1257_ vssd1 vssd1 vccd1 vccd1 _1830_ sky130_fd_sc_hd__or2_2
XFILLER_32_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2804_ _0840_ tms1x00.RAM\[14\]\[3\] _0780_ vssd1 vssd1 vccd1 vccd1 _1194_ sky130_fd_sc_hd__o21a_1
X_3784_ _1710_ tms1x00.RAM\[80\]\[3\] _1786_ vssd1 vssd1 vccd1 vccd1 _1790_ sky130_fd_sc_hd__mux2_1
XFILLER_9_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2735_ _0041_ _1056_ _1080_ _1104_ _1125_ vssd1 vssd1 vccd1 vccd1 _1126_ sky130_fd_sc_hd__o32a_1
X_2666_ tms1x00.RAM\[16\]\[2\] tms1x00.RAM\[17\]\[2\] tms1x00.RAM\[18\]\[2\] tms1x00.RAM\[19\]\[2\]
+ _0955_ _0956_ vssd1 vssd1 vccd1 vccd1 _1057_ sky130_fd_sc_hd__mux4_2
X_4405_ clknet_leaf_35_wb_clk_i _0034_ vssd1 vssd1 vccd1 vccd1 wbs_o_buff\[9\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__3862__B _1317_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2514__A3 _0903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2597_ tms1x00.RAM\[30\]\[1\] tms1x00.RAM\[31\]\[1\] _0816_ vssd1 vssd1 vccd1 vccd1
+ _0989_ sky130_fd_sc_hd__mux2_1
X_4336_ _2149_ vssd1 vssd1 vccd1 vccd1 _0630_ sky130_fd_sc_hd__clkbuf_1
XFILLER_75_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4267_ _1250_ _1317_ vssd1 vssd1 vccd1 vccd1 _2111_ sky130_fd_sc_hd__nor2_2
XFILLER_74_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4198_ _0766_ _2064_ vssd1 vssd1 vccd1 vccd1 _2065_ sky130_fd_sc_hd__and2_1
XANTENNA__4730__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3475__A1 _1578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_31_wb_clk_i clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_3218_ tms1x00.RAM\[11\]\[3\] _1463_ _1457_ vssd1 vssd1 vccd1 vccd1 _1464_ sky130_fd_sc_hd__mux2_1
XFILLER_55_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3149_ _1423_ vssd1 vssd1 vccd1 vccd1 _0169_ sky130_fd_sc_hd__clkbuf_1
XFILLER_82_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4880__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3227__A1 _1463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4214__A _0766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3529__S _1639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3163__A0 _1361_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2910__A0 _1130_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_14_wb_clk_i_A clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_65_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3218__A1 _1463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4603__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2520_ tms1x00.ram_addr_buff\[4\] tms1x00.ram_addr_buff\[5\] tms1x00.ram_addr_buff\[6\]
+ vssd1 vssd1 vccd1 vccd1 _0913_ sky130_fd_sc_hd__nand3b_4
XFILLER_6_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2451_ _0798_ _0841_ _0843_ _0775_ vssd1 vssd1 vccd1 vccd1 _0844_ sky130_fd_sc_hd__o211a_1
XFILLER_69_703 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4753__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2382_ _0774_ vssd1 vssd1 vccd1 vccd1 _0775_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__2298__B _0704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4121_ _2000_ vssd1 vssd1 vccd1 vccd1 _0564_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4052_ _0733_ _0730_ _0763_ _1918_ vssd1 vssd1 vccd1 vccd1 _1952_ sky130_fd_sc_hd__and4_1
XFILLER_49_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput4 io_in[8] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_1
X_3003_ tms1x00.ram_addr_buff\[0\] tms1x00.ram_addr_buff\[1\] _1238_ vssd1 vssd1 vccd1
+ vccd1 _1336_ sky130_fd_sc_hd__or3_1
XFILLER_37_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3209__A1 _1456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4954_ clknet_leaf_5_wb_clk_i _0564_ vssd1 vssd1 vccd1 vccd1 tms1x00.PA\[1\] sky130_fd_sc_hd__dfxtp_1
X_3905_ _1823_ tms1x00.RAM\[94\]\[3\] _1855_ vssd1 vssd1 vccd1 vccd1 _1859_ sky130_fd_sc_hd__mux2_1
XFILLER_33_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4885_ clknet_leaf_21_wb_clk_i _0499_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[91\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3836_ _1819_ tms1x00.RAM\[83\]\[1\] _1817_ vssd1 vssd1 vccd1 vccd1 _1820_ sky130_fd_sc_hd__mux2_1
XANTENNA__2815__S0 _0826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3767_ _1780_ vssd1 vssd1 vccd1 vccd1 _0430_ sky130_fd_sc_hd__clkbuf_1
X_2718_ tms1x00.RAM\[112\]\[2\] tms1x00.RAM\[113\]\[2\] tms1x00.RAM\[114\]\[2\] tms1x00.RAM\[115\]\[2\]
+ _0873_ _0822_ vssd1 vssd1 vccd1 vccd1 _1109_ sky130_fd_sc_hd__mux4_1
XANTENNA__3393__A0 _1490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2196__A1 wbs_o_buff\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3698_ _1740_ vssd1 vssd1 vccd1 vccd1 _0401_ sky130_fd_sc_hd__clkbuf_1
X_2649_ _0940_ _1037_ _1039_ _0942_ vssd1 vssd1 vccd1 vccd1 _1040_ sky130_fd_sc_hd__o211a_1
XFILLER_59_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4319_ _1823_ tms1x00.RAM\[12\]\[3\] _2136_ vssd1 vssd1 vccd1 vccd1 _2140_ sky130_fd_sc_hd__mux2_1
XFILLER_0_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3448__A1 _1578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4626__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3384__A0 _1490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input63_A wbs_dat_i[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2862__A _1129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4670_ clknet_leaf_3_wb_clk_i _0042_ vssd1 vssd1 vccd1 vccd1 _0035_ sky130_fd_sc_hd__dfxtp_2
XFILLER_30_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3621_ _1590_ tms1x00.RAM\[63\]\[2\] _1693_ vssd1 vssd1 vccd1 vccd1 _1696_ sky130_fd_sc_hd__mux2_1
X_3552_ tms1x00.RAM\[52\]\[1\] _1574_ _1654_ vssd1 vssd1 vccd1 vccd1 _1656_ sky130_fd_sc_hd__mux2_1
X_2503_ _0778_ tms1x00.RAM\[54\]\[0\] _0812_ vssd1 vssd1 vccd1 vccd1 _0896_ sky130_fd_sc_hd__o21a_1
X_3483_ _1617_ vssd1 vssd1 vccd1 vccd1 _0309_ sky130_fd_sc_hd__clkbuf_1
X_2434_ tms1x00.RAM\[68\]\[0\] tms1x00.RAM\[69\]\[0\] _0826_ vssd1 vssd1 vccd1 vccd1
+ _0827_ sky130_fd_sc_hd__mux2_1
X_2365_ _0759_ vssd1 vssd1 vccd1 vccd1 _0760_ sky130_fd_sc_hd__buf_2
XFILLER_57_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4104_ tms1x00.PA\[0\] _1978_ _1988_ vssd1 vssd1 vccd1 vccd1 _0559_ sky130_fd_sc_hd__o21a_1
XFILLER_69_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2296_ wbs_o_buff\[27\] _0704_ vssd1 vssd1 vccd1 vccd1 _0708_ sky130_fd_sc_hd__and2_1
XANTENNA__2248__S net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4035_ _0755_ _0730_ _1915_ vssd1 vssd1 vccd1 vccd1 _1940_ sky130_fd_sc_hd__or3b_1
XFILLER_49_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4649__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2653__A2 _1041_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2772__A _0996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4937_ clknet_leaf_7_wb_clk_i _0547_ vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__dfxtp_2
XANTENNA__4799__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4868_ clknet_leaf_22_wb_clk_i _0482_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[88\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_3819_ _1809_ vssd1 vssd1 vccd1 vccd1 _0453_ sky130_fd_sc_hd__clkbuf_1
XFILLER_21_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4799_ clknet_leaf_22_wb_clk_i _0413_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[6\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2801__C1 _0775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3357__A0 _1490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3109__A0 _1366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4941__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2983_ _1321_ vssd1 vssd1 vccd1 vccd1 _0105_ sky130_fd_sc_hd__clkbuf_1
X_4722_ clknet_leaf_28_wb_clk_i _0336_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[53\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2494__S1 _0800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3348__A0 _1490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4653_ clknet_leaf_5_wb_clk_i _0274_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[34\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput40 ram_val[4] vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__clkbuf_2
XANTENNA__4312__A _1344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4584_ clknet_leaf_1_wb_clk_i _0205_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[117\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput51 wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__clkbuf_1
Xinput62 wbs_dat_i[1] vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__clkbuf_1
X_3604_ _1686_ vssd1 vssd1 vccd1 vccd1 _0361_ sky130_fd_sc_hd__clkbuf_1
X_3535_ _1646_ vssd1 vssd1 vccd1 vccd1 _0332_ sky130_fd_sc_hd__clkbuf_1
X_3466_ _1592_ tms1x00.RAM\[44\]\[3\] _1604_ vssd1 vssd1 vccd1 vccd1 _1608_ sky130_fd_sc_hd__mux2_1
X_2417_ _0807_ _0809_ vssd1 vssd1 vccd1 vccd1 _0810_ sky130_fd_sc_hd__or2_1
X_3397_ _1251_ _1524_ vssd1 vssd1 vccd1 vccd1 _1566_ sky130_fd_sc_hd__or2_2
XANTENNA__3520__A0 _1592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2348_ tms1x00.ins_in\[3\] vssd1 vssd1 vccd1 vccd1 _0743_ sky130_fd_sc_hd__buf_2
XANTENNA__4471__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2279_ net83 _0702_ _0703_ wbs_o_buff\[14\] vssd1 vssd1 vccd1 vccd1 _0008_ sky130_fd_sc_hd__a22o_1
X_4018_ _0753_ _1926_ _1927_ _1901_ vssd1 vssd1 vccd1 vccd1 _0534_ sky130_fd_sc_hd__o211a_1
XFILLER_26_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3598__A _1284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3823__A1 _1772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3339__A0 _1490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4000__A1 net76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2562__A1 _0928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3511__A0 _1592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2677__A _0813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4814__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input26_A ram_val[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3814__A1 _1772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2476__S1 _0780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output94_A net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3320_ _1522_ vssd1 vssd1 vccd1 vccd1 _0241_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4494__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3251_ _1482_ vssd1 vssd1 vccd1 vccd1 _0212_ sky130_fd_sc_hd__clkbuf_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2202_ net49 vssd1 vssd1 vccd1 vccd1 _0668_ sky130_fd_sc_hd__clkbuf_4
X_3182_ _1442_ vssd1 vssd1 vccd1 vccd1 _0183_ sky130_fd_sc_hd__clkbuf_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3211__A _1327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2966_ _0914_ _1310_ vssd1 vssd1 vccd1 vccd1 _1311_ sky130_fd_sc_hd__nor2_2
XANTENNA__2467__S1 _0831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2897_ _1269_ vssd1 vssd1 vccd1 vccd1 _0071_ sky130_fd_sc_hd__clkbuf_1
X_4705_ clknet_leaf_3_wb_clk_i _0319_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[48\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_4636_ clknet_leaf_10_wb_clk_i _0257_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[2\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_4567_ clknet_leaf_35_wb_clk_i _0188_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[121\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_4498_ clknet_leaf_16_wb_clk_i _0119_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[98\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_3518_ _1590_ tms1x00.RAM\[47\]\[2\] _1634_ vssd1 vssd1 vccd1 vccd1 _1637_ sky130_fd_sc_hd__mux2_1
XFILLER_77_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3449_ _1598_ vssd1 vssd1 vccd1 vccd1 _0294_ sky130_fd_sc_hd__clkbuf_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3820__S _1806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2944__B _1249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2232__A0 net30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapped_tms1x00_170 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_170/HI io_oeb[31] sky130_fd_sc_hd__conb_1
Xwrapped_tms1x00_181 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_181/HI io_out[4] sky130_fd_sc_hd__conb_1
XANTENNA__3980__B1 _1900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2783__A1 _0940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapped_tms1x00_192 vssd1 vssd1 vccd1 vccd1 io_oeb[2] wrapped_tms1x00_192/LO sky130_fd_sc_hd__conb_1
XFILLER_4_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4288__A1 _1327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3966__A tms1x00.wb_step vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2449__S1 _0779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2820_ _0931_ tms1x00.RAM\[54\]\[3\] _0791_ vssd1 vssd1 vccd1 vccd1 _1210_ sky130_fd_sc_hd__o21a_1
X_2751_ _1137_ _1139_ _1140_ _0922_ _0942_ vssd1 vssd1 vccd1 vccd1 _1141_ sky130_fd_sc_hd__o221a_1
XANTENNA__3971__A0 _0742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2682_ tms1x00.RAM\[8\]\[2\] tms1x00.RAM\[9\]\[2\] tms1x00.RAM\[10\]\[2\] tms1x00.RAM\[11\]\[2\]
+ _0830_ _0800_ vssd1 vssd1 vccd1 vccd1 _1073_ sky130_fd_sc_hd__mux4_1
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4421_ clknet_leaf_27_wb_clk_i _0020_ vssd1 vssd1 vccd1 vccd1 wbs_o_buff\[25\] sky130_fd_sc_hd__dfxtp_1
X_4352_ _2158_ vssd1 vssd1 vccd1 vccd1 _0637_ sky130_fd_sc_hd__clkbuf_1
X_4283_ _1823_ tms1x00.RAM\[29\]\[3\] _2116_ vssd1 vssd1 vccd1 vccd1 _2120_ sky130_fd_sc_hd__mux2_1
X_3303_ _1492_ tms1x00.RAM\[28\]\[3\] _1509_ vssd1 vssd1 vccd1 vccd1 _1513_ sky130_fd_sc_hd__mux2_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3234_ tms1x00.RAM\[117\]\[2\] _1461_ _1470_ vssd1 vssd1 vccd1 vccd1 _1473_ sky130_fd_sc_hd__mux2_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3165_ _1364_ tms1x00.RAM\[124\]\[1\] _1431_ vssd1 vssd1 vccd1 vccd1 _1433_ sky130_fd_sc_hd__mux2_1
XFILLER_82_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3096_ _1392_ vssd1 vssd1 vccd1 vccd1 _0147_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3998_ _0701_ _1908_ net75 vssd1 vssd1 vccd1 vccd1 _1913_ sky130_fd_sc_hd__a21o_1
XFILLER_50_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2949_ _1130_ tms1x00.RAM\[19\]\[2\] _1297_ vssd1 vssd1 vccd1 vccd1 _1300_ sky130_fd_sc_hd__mux2_1
XANTENNA__2765__A1 _0920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4619_ clknet_leaf_0_wb_clk_i _0240_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[26\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3190__A1 _1324_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2955__A _0914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3786__A _1310_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4381__S _2006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2205__A0 net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_1_wb_clk_i clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_79_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3181__A1 _1324_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3026__A _0913_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2865__A _1224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4970_ clknet_leaf_9_wb_clk_i _0580_ vssd1 vssd1 vccd1 vccd1 tms1x00.Y\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3921_ _1821_ tms1x00.RAM\[92\]\[2\] _1865_ vssd1 vssd1 vccd1 vccd1 _1868_ sky130_fd_sc_hd__mux2_1
XANTENNA__4682__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3852_ _1829_ vssd1 vssd1 vccd1 vccd1 _0466_ sky130_fd_sc_hd__clkbuf_1
XFILLER_32_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4197__A0 tms1x00.Y\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2803_ tms1x00.RAM\[15\]\[3\] _0840_ vssd1 vssd1 vccd1 vccd1 _1193_ sky130_fd_sc_hd__or2b_1
X_3783_ _1789_ vssd1 vssd1 vccd1 vccd1 _0437_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5038__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2734_ _0040_ _1115_ _1124_ _0835_ vssd1 vssd1 vccd1 vccd1 _1125_ sky130_fd_sc_hd__a31o_1
X_2665_ _0821_ _1040_ _1044_ _0040_ _1055_ vssd1 vssd1 vccd1 vccd1 _1056_ sky130_fd_sc_hd__o311a_1
X_2596_ _0818_ _0987_ vssd1 vssd1 vccd1 vccd1 _0988_ sky130_fd_sc_hd__and2_1
X_4404_ clknet_leaf_35_wb_clk_i _0033_ vssd1 vssd1 vccd1 vccd1 wbs_o_buff\[8\] sky130_fd_sc_hd__dfxtp_1
X_4335_ _1245_ tms1x00.RAM\[15\]\[2\] _2146_ vssd1 vssd1 vccd1 vccd1 _2149_ sky130_fd_sc_hd__mux2_1
XANTENNA__3172__A1 _1324_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4266_ _2110_ vssd1 vssd1 vccd1 vccd1 _0599_ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4197_ tms1x00.Y\[0\] _2062_ _2063_ vssd1 vssd1 vccd1 vccd1 _2064_ sky130_fd_sc_hd__mux2_1
X_3217_ _1333_ vssd1 vssd1 vccd1 vccd1 _1463_ sky130_fd_sc_hd__buf_2
XFILLER_67_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3148_ tms1x00.RAM\[106\]\[2\] _1331_ _1420_ vssd1 vssd1 vccd1 vccd1 _1423_ sky130_fd_sc_hd__mux2_1
XFILLER_54_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3079_ _1364_ tms1x00.RAM\[113\]\[1\] _1381_ vssd1 vssd1 vccd1 vccd1 _1383_ sky130_fd_sc_hd__mux2_1
XFILLER_54_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4188__B1 _0760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3935__A0 tms1x00.RAM\[90\]\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4360__A0 _1243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3455__S _1599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2450_ _0828_ _0842_ vssd1 vssd1 vccd1 vccd1 _0843_ sky130_fd_sc_hd__or2_1
XFILLER_6_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4351__A0 _1243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2381_ _0038_ vssd1 vssd1 vccd1 vccd1 _0774_ sky130_fd_sc_hd__inv_2
XFILLER_68_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4120_ net103 _1999_ vssd1 vssd1 vccd1 vccd1 _2000_ sky130_fd_sc_hd__or2_1
XFILLER_68_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4051_ net90 _1950_ _1951_ _1931_ vssd1 vssd1 vccd1 vccd1 _0543_ sky130_fd_sc_hd__o211a_1
Xinput5 io_in[9] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_1
XFILLER_65_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3002_ _1335_ vssd1 vssd1 vccd1 vccd1 _0110_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__2665__B1 _0040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4953_ clknet_leaf_6_wb_clk_i _0563_ vssd1 vssd1 vccd1 vccd1 tms1x00.PA\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_17_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3090__A0 _1366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3904_ _1858_ vssd1 vssd1 vccd1 vccd1 _0489_ sky130_fd_sc_hd__clkbuf_1
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4884_ clknet_leaf_17_wb_clk_i _0498_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[92\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3917__A0 _1816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3835_ _1034_ vssd1 vssd1 vccd1 vccd1 _1819_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__4428__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3766_ tms1x00.RAM\[74\]\[3\] _1779_ _1773_ vssd1 vssd1 vccd1 vccd1 _1780_ sky130_fd_sc_hd__mux2_1
X_2717_ _1105_ _1106_ _1107_ _0818_ _0953_ vssd1 vssd1 vccd1 vccd1 _1108_ sky130_fd_sc_hd__a221o_1
XANTENNA__2815__S1 _0780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4578__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3697_ tms1x00.RAM\[72\]\[2\] _1674_ _1737_ vssd1 vssd1 vccd1 vccd1 _1740_ sky130_fd_sc_hd__mux2_1
XANTENNA__4342__A0 _1243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2648_ _0807_ _1038_ vssd1 vssd1 vccd1 vccd1 _1039_ sky130_fd_sc_hd__or2_1
XANTENNA__2579__S0 _0808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2579_ tms1x00.RAM\[120\]\[1\] tms1x00.RAM\[121\]\[1\] tms1x00.RAM\[122\]\[1\] tms1x00.RAM\[123\]\[1\]
+ _0808_ _0831_ vssd1 vssd1 vccd1 vccd1 _0971_ sky130_fd_sc_hd__mux4_2
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4318_ _2139_ vssd1 vssd1 vccd1 vccd1 _0622_ sky130_fd_sc_hd__clkbuf_1
XFILLER_75_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2709__S _0788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4249_ _1310_ _1430_ vssd1 vssd1 vccd1 vccd1 _2101_ sky130_fd_sc_hd__nor2_2
XFILLER_68_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3081__A0 _1366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3908__A0 _1816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4333__A0 _1243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input56_A wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2742__S0 _0931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3072__A0 _1366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3620_ _1695_ vssd1 vssd1 vccd1 vccd1 _0368_ sky130_fd_sc_hd__clkbuf_1
X_3551_ _1655_ vssd1 vssd1 vccd1 vccd1 _0339_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__3375__A1 _1461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2502_ tms1x00.RAM\[55\]\[0\] _0778_ vssd1 vssd1 vccd1 vccd1 _0895_ sky130_fd_sc_hd__or2b_1
XANTENNA__4324__A0 _1819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3482_ tms1x00.RAM\[42\]\[2\] _1576_ _1614_ vssd1 vssd1 vccd1 vccd1 _1617_ sky130_fd_sc_hd__mux2_1
X_2433_ _0035_ vssd1 vssd1 vccd1 vccd1 _0826_ sky130_fd_sc_hd__buf_6
X_2364_ net148 _0721_ vssd1 vssd1 vccd1 vccd1 _0759_ sky130_fd_sc_hd__and2_1
X_4103_ tms1x00.PB\[0\] _0738_ _1987_ vssd1 vssd1 vccd1 vccd1 _1988_ sky130_fd_sc_hd__or3b_1
XFILLER_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3214__A _1330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2295_ _0707_ vssd1 vssd1 vccd1 vccd1 _0021_ sky130_fd_sc_hd__clkbuf_1
XFILLER_65_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4034_ _0755_ _0741_ _0753_ _1939_ _0766_ vssd1 vssd1 vccd1 vccd1 _0538_ sky130_fd_sc_hd__o311a_1
XFILLER_2_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4936_ clknet_leaf_8_wb_clk_i _0546_ vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__dfxtp_2
XFILLER_33_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4867_ clknet_leaf_22_wb_clk_i _0481_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[88\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_3818_ tms1x00.RAM\[85\]\[2\] _1777_ _1806_ vssd1 vssd1 vccd1 vccd1 _1809_ sky130_fd_sc_hd__mux2_1
XANTENNA__3366__A1 _1461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4798_ clknet_leaf_22_wb_clk_i _0412_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[6\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3749_ tms1x00.RAM\[75\]\[1\] _1672_ _1767_ vssd1 vssd1 vccd1 vccd1 _1769_ sky130_fd_sc_hd__mux2_1
XANTENNA__4315__A0 _1819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3118__A1 _1328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3823__S _1811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4743__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2801__B1 _1190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4893__CLK clknet_leaf_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2982_ tms1x00.RAM\[102\]\[2\] _1245_ _1318_ vssd1 vssd1 vccd1 vccd1 _1321_ sky130_fd_sc_hd__mux2_1
XFILLER_21_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3596__A1 _1676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4721_ clknet_leaf_28_wb_clk_i _0335_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[53\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_4652_ clknet_leaf_6_wb_clk_i _0273_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[34\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput30 ram_val[24] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__dlymetal6s2s_1
X_3603_ tms1x00.RAM\[56\]\[2\] _1674_ _1683_ vssd1 vssd1 vccd1 vccd1 _1686_ sky130_fd_sc_hd__mux2_1
XANTENNA__4312__B _1409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4583_ clknet_leaf_0_wb_clk_i _0204_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[117\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput52 wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__clkbuf_1
Xinput63 wbs_dat_i[2] vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__clkbuf_1
Xinput41 ram_val[5] vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__clkbuf_2
X_3534_ tms1x00.RAM\[54\]\[1\] _1574_ _1644_ vssd1 vssd1 vccd1 vccd1 _1646_ sky130_fd_sc_hd__mux2_1
X_3465_ _1607_ vssd1 vssd1 vccd1 vccd1 _0301_ sky130_fd_sc_hd__clkbuf_1
X_2416_ tms1x00.RAM\[72\]\[0\] tms1x00.RAM\[73\]\[0\] tms1x00.RAM\[74\]\[0\] tms1x00.RAM\[75\]\[0\]
+ _0808_ _0780_ vssd1 vssd1 vccd1 vccd1 _0809_ sky130_fd_sc_hd__mux4_1
X_3396_ _1565_ vssd1 vssd1 vccd1 vccd1 _0274_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4616__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2347_ tms1x00.ins_in\[0\] vssd1 vssd1 vccd1 vccd1 _0742_ sky130_fd_sc_hd__buf_2
XFILLER_29_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2278_ net82 _0702_ _0703_ wbs_o_buff\[13\] vssd1 vssd1 vccd1 vccd1 _0007_ sky130_fd_sc_hd__a22o_1
X_4017_ _0755_ _0730_ _0740_ _0764_ net81 vssd1 vssd1 vccd1 vccd1 _1927_ sky130_fd_sc_hd__a41o_1
XFILLER_38_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2706__S0 _0873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3598__B _1303_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4766__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3036__A0 _0912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4919_ clknet_leaf_8_wb_clk_i tms1x00.K_in\[2\] vssd1 vssd1 vccd1 vccd1 tms1x00.K_latch\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_52_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3587__A1 _1676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2795__C1 _0942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3818__S _1806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input19_A ram_val[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3027__A0 _0912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3578__A1 _1669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2250__A1 K_override\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4132__B _0768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output87_A net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4639__CLK clknet_leaf_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3250_ _1364_ tms1x00.RAM\[115\]\[1\] _1480_ vssd1 vssd1 vccd1 vccd1 _1482_ sky130_fd_sc_hd__mux2_1
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2201_ _0667_ vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__clkbuf_1
XANTENNA__3502__A1 _1578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3181_ tms1x00.RAM\[122\]\[0\] _1324_ _1441_ vssd1 vssd1 vccd1 vccd1 _1442_ sky130_fd_sc_hd__mux2_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4789__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2710__C1 _0794_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3018__A0 _0912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2965_ _1309_ vssd1 vssd1 vccd1 vccd1 _1310_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__2777__C1 _0996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4704_ clknet_leaf_28_wb_clk_i _0318_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[4\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_2896_ _0912_ tms1x00.RAM\[79\]\[0\] _1268_ vssd1 vssd1 vccd1 vccd1 _1269_ sky130_fd_sc_hd__mux2_1
XANTENNA__4042__B _0752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4635_ clknet_leaf_10_wb_clk_i _0256_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[2\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_25_wb_clk_i clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_4566_ clknet_leaf_1_wb_clk_i _0187_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[121\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_3517_ _1636_ vssd1 vssd1 vccd1 vccd1 _0324_ sky130_fd_sc_hd__clkbuf_1
X_4497_ clknet_leaf_11_wb_clk_i _0118_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[0\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3448_ tms1x00.RAM\[38\]\[3\] _1578_ _1594_ vssd1 vssd1 vccd1 vccd1 _1598_ sky130_fd_sc_hd__mux2_1
XFILLER_76_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3379_ _1229_ _1525_ vssd1 vssd1 vccd1 vccd1 _1556_ sky130_fd_sc_hd__or2_2
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_3__f_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_2_3__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_43_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapped_tms1x00_171 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_171/HI io_oeb[32] sky130_fd_sc_hd__conb_1
Xwrapped_tms1x00_160 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_160/HI io_oeb[21] sky130_fd_sc_hd__conb_1
Xwrapped_tms1x00_182 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_182/HI io_out[5] sky130_fd_sc_hd__conb_1
Xwrapped_tms1x00_193 vssd1 vssd1 vccd1 vccd1 io_oeb[3] wrapped_tms1x00_193/LO sky130_fd_sc_hd__conb_1
XANTENNA__4379__S _2006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_33_wb_clk_i_A clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_4_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2688__A _0039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4931__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3248__A0 _1361_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3966__B _0766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2750_ tms1x00.RAM\[88\]\[3\] tms1x00.RAM\[89\]\[3\] tms1x00.RAM\[90\]\[3\] tms1x00.RAM\[91\]\[3\]
+ _0931_ _0932_ vssd1 vssd1 vccd1 vccd1 _1140_ sky130_fd_sc_hd__mux4_1
XFILLER_31_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3971__A1 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2681_ _1068_ _1070_ _1071_ _0807_ _0774_ vssd1 vssd1 vccd1 vccd1 _1072_ sky130_fd_sc_hd__o221a_1
X_4420_ clknet_leaf_32_wb_clk_i _0019_ vssd1 vssd1 vccd1 vccd1 wbs_o_buff\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_8_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4351_ _1243_ tms1x00.RAM\[13\]\[1\] _2156_ vssd1 vssd1 vccd1 vccd1 _2158_ sky130_fd_sc_hd__mux2_1
X_3302_ _1512_ vssd1 vssd1 vccd1 vccd1 _0233_ sky130_fd_sc_hd__clkbuf_1
X_4282_ _2119_ vssd1 vssd1 vccd1 vccd1 _0606_ sky130_fd_sc_hd__clkbuf_1
XFILLER_4_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3487__A0 _1585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3233_ _1472_ vssd1 vssd1 vccd1 vccd1 _0204_ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4963__D _0573_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3164_ _1432_ vssd1 vssd1 vccd1 vccd1 _0175_ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3095_ _1361_ tms1x00.RAM\[111\]\[0\] _1391_ vssd1 vssd1 vccd1 vccd1 _1392_ sky130_fd_sc_hd__mux2_1
XFILLER_39_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2537__S _0924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3997_ net76 net75 vssd1 vssd1 vccd1 vccd1 _1912_ sky130_fd_sc_hd__nor2_1
XFILLER_50_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4804__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2948_ _1299_ vssd1 vssd1 vccd1 vccd1 _0092_ sky130_fd_sc_hd__clkbuf_1
XFILLER_10_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2879_ _1256_ vssd1 vssd1 vccd1 vccd1 _0066_ sky130_fd_sc_hd__clkbuf_1
X_4618_ clknet_leaf_0_wb_clk_i _0239_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[26\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4954__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4549_ clknet_leaf_31_wb_clk_i _0170_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[106\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_77_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2955__B _1303_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3650__A0 _1706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3786__B _1344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3402__A0 _1490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3026__B _1273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2881__A _1257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3977__A _0701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3920_ _1867_ vssd1 vssd1 vccd1 vccd1 _0496_ sky130_fd_sc_hd__clkbuf_1
XFILLER_45_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4827__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3851_ _1823_ tms1x00.RAM\[82\]\[3\] _1825_ vssd1 vssd1 vccd1 vccd1 _1829_ sky130_fd_sc_hd__mux2_1
XFILLER_32_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3782_ _1708_ tms1x00.RAM\[80\]\[2\] _1786_ vssd1 vssd1 vccd1 vccd1 _1789_ sky130_fd_sc_hd__mux2_1
X_2802_ tms1x00.RAM\[8\]\[3\] tms1x00.RAM\[9\]\[3\] tms1x00.RAM\[10\]\[3\] tms1x00.RAM\[11\]\[3\]
+ _0816_ _0927_ vssd1 vssd1 vccd1 vccd1 _1192_ sky130_fd_sc_hd__mux4_1
XANTENNA__4977__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2733_ _0776_ _1117_ _1119_ _0821_ _1123_ vssd1 vssd1 vccd1 vccd1 _1124_ sky130_fd_sc_hd__a311o_1
XFILLER_13_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3944__A1 _1323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2664_ _0776_ _1048_ _1050_ _0804_ _1054_ vssd1 vssd1 vccd1 vccd1 _1055_ sky130_fd_sc_hd__a311o_1
X_2595_ tms1x00.RAM\[28\]\[1\] tms1x00.RAM\[29\]\[1\] _0873_ vssd1 vssd1 vccd1 vccd1
+ _0987_ sky130_fd_sc_hd__mux2_1
X_4403_ clknet_leaf_35_wb_clk_i _0032_ vssd1 vssd1 vccd1 vccd1 wbs_o_buff\[7\] sky130_fd_sc_hd__dfxtp_1
X_4334_ _2148_ vssd1 vssd1 vccd1 vccd1 _0629_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__3217__A _1333_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4265_ tms1x00.RAM\[39\]\[3\] _1333_ _2106_ vssd1 vssd1 vccd1 vccd1 _2110_ sky130_fd_sc_hd__mux2_1
X_4196_ tms1x00.ins_in\[4\] _0746_ _1127_ tms1x00.ins_in\[5\] vssd1 vssd1 vccd1 vccd1
+ _2063_ sky130_fd_sc_hd__nor4b_4
XFILLER_55_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3216_ _1462_ vssd1 vssd1 vccd1 vccd1 _0197_ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3147_ _1422_ vssd1 vssd1 vccd1 vccd1 _0168_ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3078_ _1382_ vssd1 vssd1 vccd1 vccd1 _0139_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3632__A0 _1592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2791__A _0928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4188__A1 tms1x00.PC\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3935__A1 _1323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2966__A _0914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3623__A0 _1592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2206__A _0670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3926__A1 _1772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2380_ _0040_ vssd1 vssd1 vccd1 vccd1 _0773_ sky130_fd_sc_hd__clkinv_2
X_4050_ _0755_ _0752_ _1928_ vssd1 vssd1 vccd1 vccd1 _1951_ sky130_fd_sc_hd__or3_1
XFILLER_49_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2665__A1 _0821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput6 oram_value[0] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__dlymetal6s2s_1
X_3001_ tms1x00.RAM\[101\]\[3\] _1334_ _1325_ vssd1 vssd1 vccd1 vccd1 _1335_ sky130_fd_sc_hd__mux2_1
XFILLER_65_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5005__CLK clknet_leaf_20_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4952_ clknet_leaf_5_wb_clk_i _0562_ vssd1 vssd1 vccd1 vccd1 tms1x00.PB\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_45_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3903_ _1821_ tms1x00.RAM\[94\]\[2\] _1855_ vssd1 vssd1 vccd1 vccd1 _1858_ sky130_fd_sc_hd__mux2_1
X_4883_ clknet_leaf_15_wb_clk_i _0497_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[92\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_3834_ _1818_ vssd1 vssd1 vccd1 vccd1 _0459_ sky130_fd_sc_hd__clkbuf_1
XFILLER_20_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3765_ _1224_ vssd1 vssd1 vccd1 vccd1 _1779_ sky130_fd_sc_hd__clkbuf_4
X_2716_ tms1x00.RAM\[116\]\[2\] tms1x00.RAM\[117\]\[2\] _0789_ vssd1 vssd1 vccd1 vccd1
+ _1107_ sky130_fd_sc_hd__mux2_1
XFILLER_9_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3696_ _1739_ vssd1 vssd1 vccd1 vccd1 _0400_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4050__B _0752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2647_ tms1x00.RAM\[40\]\[2\] tms1x00.RAM\[41\]\[2\] tms1x00.RAM\[42\]\[2\] tms1x00.RAM\[43\]\[2\]
+ _0830_ _0831_ vssd1 vssd1 vccd1 vccd1 _1038_ sky130_fd_sc_hd__mux4_1
X_2578_ tms1x00.RAM\[124\]\[1\] tms1x00.RAM\[125\]\[1\] tms1x00.RAM\[126\]\[1\] tms1x00.RAM\[127\]\[1\]
+ _0945_ _0956_ vssd1 vssd1 vccd1 vccd1 _0970_ sky130_fd_sc_hd__mux4_1
XFILLER_0_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2579__S1 _0831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4317_ _1821_ tms1x00.RAM\[12\]\[2\] _2136_ vssd1 vssd1 vccd1 vccd1 _2139_ sky130_fd_sc_hd__mux2_1
X_4248_ _2100_ vssd1 vssd1 vccd1 vccd1 _0591_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4179_ tms1x00.PC\[3\] _2043_ vssd1 vssd1 vccd1 vccd1 _2048_ sky130_fd_sc_hd__and2_1
XFILLER_35_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3410__A _1034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4387__S _2006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input49_A wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4672__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2742__S1 _0932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3550_ tms1x00.RAM\[52\]\[0\] _1571_ _1654_ vssd1 vssd1 vccd1 vccd1 _1655_ sky130_fd_sc_hd__mux2_1
X_2501_ _0828_ _0893_ _0038_ vssd1 vssd1 vccd1 vccd1 _0894_ sky130_fd_sc_hd__o21a_1
X_3481_ _1616_ vssd1 vssd1 vccd1 vccd1 _0308_ sky130_fd_sc_hd__clkbuf_1
XFILLER_69_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2432_ _0822_ _0824_ vssd1 vssd1 vccd1 vccd1 _0825_ sky130_fd_sc_hd__and2_1
X_2363_ _0749_ vssd1 vssd1 vccd1 vccd1 _0758_ sky130_fd_sc_hd__inv_2
XANTENNA__2886__A1 _1235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4102_ _0722_ _0758_ _1986_ _1973_ vssd1 vssd1 vccd1 vccd1 _1987_ sky130_fd_sc_hd__a31oi_4
X_4033_ _0733_ _0756_ _0764_ net85 vssd1 vssd1 vccd1 vccd1 _1939_ sky130_fd_sc_hd__a31o_1
X_2294_ wbs_o_buff\[26\] _0704_ vssd1 vssd1 vccd1 vccd1 _0707_ sky130_fd_sc_hd__and2_1
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2638__A1 _0960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4045__B tms1x00.Y\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4935_ clknet_leaf_13_wb_clk_i _0545_ vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__dfxtp_4
X_4866_ clknet_leaf_21_wb_clk_i _0480_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[88\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4545__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3817_ _1808_ vssd1 vssd1 vccd1 vccd1 _0452_ sky130_fd_sc_hd__clkbuf_1
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4797_ clknet_leaf_22_wb_clk_i _0411_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[6\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3748_ _1768_ vssd1 vssd1 vccd1 vccd1 _0423_ sky130_fd_sc_hd__clkbuf_1
XFILLER_4_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4695__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3679_ _1708_ tms1x00.RAM\[65\]\[2\] _1727_ vssd1 vssd1 vccd1 vccd1 _1730_ sky130_fd_sc_hd__mux2_1
XANTENNA__2326__A0 tms1x00.Y\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput140 net140 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[31] sky130_fd_sc_hd__buf_2
XFILLER_0_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2801__B2 _0921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2660__S0 _0840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4306__A1 _1327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4418__CLK clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4568__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2981_ _1320_ vssd1 vssd1 vccd1 vccd1 _0104_ sky130_fd_sc_hd__clkbuf_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4720_ clknet_leaf_29_wb_clk_i _0334_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[54\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_4651_ clknet_leaf_6_wb_clk_i _0272_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[34\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput31 ram_val[25] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput20 ram_val[15] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__dlymetal6s2s_1
X_3602_ _1685_ vssd1 vssd1 vccd1 vccd1 _0360_ sky130_fd_sc_hd__clkbuf_1
X_4582_ clknet_leaf_1_wb_clk_i _0203_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[117\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput42 ram_val[6] vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__clkbuf_2
Xinput53 wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__clkbuf_1
Xinput64 wbs_dat_i[3] vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__clkbuf_1
XANTENNA__2651__S0 _0799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3533_ _1645_ vssd1 vssd1 vccd1 vccd1 _0331_ sky130_fd_sc_hd__clkbuf_1
X_3464_ _1590_ tms1x00.RAM\[44\]\[2\] _1604_ vssd1 vssd1 vccd1 vccd1 _1607_ sky130_fd_sc_hd__mux2_1
X_2415_ _0777_ vssd1 vssd1 vccd1 vccd1 _0808_ sky130_fd_sc_hd__buf_8
X_3395_ _1492_ tms1x00.RAM\[34\]\[3\] _1561_ vssd1 vssd1 vccd1 vccd1 _1565_ sky130_fd_sc_hd__mux2_1
X_2346_ _0739_ _0740_ vssd1 vssd1 vccd1 vccd1 _0741_ sky130_fd_sc_hd__nand2_1
XFILLER_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2277_ net81 _0702_ _0703_ wbs_o_buff\[12\] vssd1 vssd1 vccd1 vccd1 _0006_ sky130_fd_sc_hd__a22o_1
X_4016_ _0732_ _0739_ _0740_ vssd1 vssd1 vccd1 vccd1 _1926_ sky130_fd_sc_hd__or3b_1
XANTENNA__2706__S1 _0822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_2_2__f_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_2_2__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_52_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4918_ clknet_leaf_8_wb_clk_i tms1x00.K_in\[1\] vssd1 vssd1 vccd1 vccd1 tms1x00.K_latch\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2795__B1 _1184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4849_ clknet_leaf_17_wb_clk_i _0463_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[82\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4222__C tms1x00.ins_in\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_23_wb_clk_i_A clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_4_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4710__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2633__S0 _0788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3045__A _0913_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2200_ net45 wbs_o_buff\[9\] _0657_ vssd1 vssd1 vccd1 vccd1 _0667_ sky130_fd_sc_hd__mux2_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3180_ _1430_ _1403_ vssd1 vssd1 vccd1 vccd1 _1441_ sky130_fd_sc_hd__nor2_2
XFILLER_78_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2474__C1 _0802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2964_ _1227_ _1238_ vssd1 vssd1 vccd1 vccd1 _1309_ sky130_fd_sc_hd__or2_1
XFILLER_34_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4703_ clknet_leaf_28_wb_clk_i _0317_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[4\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_2895_ _1237_ _1267_ vssd1 vssd1 vccd1 vccd1 _1268_ sky130_fd_sc_hd__or2_2
X_4634_ clknet_leaf_10_wb_clk_i _0255_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[2\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_4565_ clknet_leaf_33_wb_clk_i _0186_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[122\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_3516_ _1588_ tms1x00.RAM\[47\]\[1\] _1634_ vssd1 vssd1 vccd1 vccd1 _1636_ sky130_fd_sc_hd__mux2_1
X_4496_ clknet_leaf_11_wb_clk_i _0117_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[0\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_3447_ _1597_ vssd1 vssd1 vccd1 vccd1 _0293_ sky130_fd_sc_hd__clkbuf_1
XFILLER_58_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3378_ _1555_ vssd1 vssd1 vccd1 vccd1 _0266_ sky130_fd_sc_hd__clkbuf_1
XFILLER_69_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2329_ _0730_ tms1x00.ram_addr_buff\[2\] _0726_ vssd1 vssd1 vccd1 vccd1 _0731_ sky130_fd_sc_hd__mux2_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3829__S _1811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwrapped_tms1x00_172 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_172/HI io_oeb[33] sky130_fd_sc_hd__conb_1
Xwrapped_tms1x00_161 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_161/HI io_oeb[22] sky130_fd_sc_hd__conb_1
Xwrapped_tms1x00_150 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_150/HI io_oeb[11] sky130_fd_sc_hd__conb_1
XANTENNA__3980__A2 _0724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapped_tms1x00_183 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_183/HI io_out[6] sky130_fd_sc_hd__conb_1
Xwrapped_tms1x00_194 vssd1 vssd1 vccd1 vccd1 io_oeb[4] wrapped_tms1x00_194/LO sky130_fd_sc_hd__conb_1
XFILLER_4_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2940__A0 _1130_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3496__A1 _1571_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input31_A ram_val[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4143__B _1126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4606__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3420__A1 _1571_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2680_ tms1x00.RAM\[0\]\[2\] tms1x00.RAM\[1\]\[2\] tms1x00.RAM\[2\]\[2\] tms1x00.RAM\[3\]\[2\]
+ _0808_ _0831_ vssd1 vssd1 vccd1 vccd1 _1071_ sky130_fd_sc_hd__mux4_1
XFILLER_8_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4350_ _2157_ vssd1 vssd1 vccd1 vccd1 _0636_ sky130_fd_sc_hd__clkbuf_1
X_3301_ _1490_ tms1x00.RAM\[28\]\[2\] _1509_ vssd1 vssd1 vccd1 vccd1 _1512_ sky130_fd_sc_hd__mux2_1
X_4281_ _1821_ tms1x00.RAM\[29\]\[2\] _2116_ vssd1 vssd1 vccd1 vccd1 _2119_ sky130_fd_sc_hd__mux2_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3232_ tms1x00.RAM\[117\]\[1\] _1459_ _1470_ vssd1 vssd1 vccd1 vccd1 _1472_ sky130_fd_sc_hd__mux2_1
XFILLER_67_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3163_ _1361_ tms1x00.RAM\[124\]\[0\] _1431_ vssd1 vssd1 vccd1 vccd1 _1432_ sky130_fd_sc_hd__mux2_1
XFILLER_39_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3094_ _0913_ _1267_ vssd1 vssd1 vccd1 vccd1 _1391_ sky130_fd_sc_hd__or2_2
XFILLER_39_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3239__A1 _1456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2462__A2 _0854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3996_ _1911_ vssd1 vssd1 vccd1 vccd1 _0528_ sky130_fd_sc_hd__clkbuf_1
XFILLER_23_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4053__B _0752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2947_ _1035_ tms1x00.RAM\[19\]\[1\] _1297_ vssd1 vssd1 vccd1 vccd1 _1299_ sky130_fd_sc_hd__mux2_1
XANTENNA__3411__A1 _1574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2878_ _1225_ tms1x00.RAM\[17\]\[3\] _1252_ vssd1 vssd1 vccd1 vccd1 _1256_ sky130_fd_sc_hd__mux2_1
X_4617_ clknet_leaf_4_wb_clk_i _0238_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[27\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_4548_ clknet_leaf_31_wb_clk_i _0169_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[106\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_4479_ clknet_leaf_29_wb_clk_i _0100_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[103\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_58_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3478__A1 _1571_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3413__A _1129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4629__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3469__A1 _1571_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3977__B _0760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3850_ _1828_ vssd1 vssd1 vccd1 vccd1 _0465_ sky130_fd_sc_hd__clkbuf_1
X_3781_ _1788_ vssd1 vssd1 vccd1 vccd1 _0436_ sky130_fd_sc_hd__clkbuf_1
X_2801_ _1187_ _1189_ _1190_ _0921_ _0775_ vssd1 vssd1 vccd1 vccd1 _1191_ sky130_fd_sc_hd__o221a_1
XFILLER_13_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3993__A _0701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2601__C1 _0920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2732_ _0996_ _1120_ _1122_ _0806_ vssd1 vssd1 vccd1 vccd1 _1123_ sky130_fd_sc_hd__o211a_1
XFILLER_9_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2663_ _0953_ _1051_ _1053_ _0802_ vssd1 vssd1 vccd1 vccd1 _1054_ sky130_fd_sc_hd__o211a_1
X_2594_ _0984_ _0985_ _0921_ vssd1 vssd1 vccd1 vccd1 _0986_ sky130_fd_sc_hd__mux2_1
X_4402_ clknet_leaf_35_wb_clk_i _0031_ vssd1 vssd1 vccd1 vccd1 wbs_o_buff\[6\] sky130_fd_sc_hd__dfxtp_1
X_4333_ _1243_ tms1x00.RAM\[15\]\[1\] _2146_ vssd1 vssd1 vccd1 vccd1 _2148_ sky130_fd_sc_hd__mux2_1
XFILLER_59_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4264_ _2109_ vssd1 vssd1 vccd1 vccd1 _0598_ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3215_ tms1x00.RAM\[11\]\[2\] _1461_ _1457_ vssd1 vssd1 vccd1 vccd1 _1462_ sky130_fd_sc_hd__mux2_1
XFILLER_67_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4195_ tms1x00.P\[0\] _2061_ vssd1 vssd1 vccd1 vccd1 _2062_ sky130_fd_sc_hd__xor2_1
XFILLER_67_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3146_ tms1x00.RAM\[106\]\[1\] _1328_ _1420_ vssd1 vssd1 vccd1 vccd1 _1422_ sky130_fd_sc_hd__mux2_1
XFILLER_82_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3077_ _1361_ tms1x00.RAM\[113\]\[0\] _1381_ vssd1 vssd1 vccd1 vccd1 _1382_ sky130_fd_sc_hd__mux2_1
XFILLER_55_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3632__A1 tms1x00.RAM\[62\]\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4921__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3979_ _0718_ vssd1 vssd1 vccd1 vccd1 _1901_ sky130_fd_sc_hd__buf_4
XANTENNA__3699__A1 _1676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2966__B _1310_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3143__A _0914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4451__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2819__B_N _0931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2222__A _0678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput7 oram_value[1] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__dlymetal6s2s_1
X_3000_ _1333_ vssd1 vssd1 vccd1 vccd1 _1334_ sky130_fd_sc_hd__clkbuf_4
XFILLER_36_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4951_ clknet_leaf_6_wb_clk_i _0561_ vssd1 vssd1 vccd1 vccd1 tms1x00.PB\[2\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__3614__A1 _1676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3902_ _1857_ vssd1 vssd1 vccd1 vccd1 _0488_ sky130_fd_sc_hd__clkbuf_1
X_4882_ clknet_leaf_17_wb_clk_i _0496_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[92\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2822__C1 _0996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3833_ _1816_ tms1x00.RAM\[83\]\[0\] _1817_ vssd1 vssd1 vccd1 vccd1 _1818_ sky130_fd_sc_hd__mux2_1
XFILLER_33_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3764_ _1778_ vssd1 vssd1 vccd1 vccd1 _0429_ sky130_fd_sc_hd__clkbuf_1
X_2715_ _0945_ tms1x00.RAM\[118\]\[2\] _0927_ vssd1 vssd1 vccd1 vccd1 _1106_ sky130_fd_sc_hd__o21a_1
X_3695_ tms1x00.RAM\[72\]\[1\] _1672_ _1737_ vssd1 vssd1 vccd1 vccd1 _1739_ sky130_fd_sc_hd__mux2_1
X_2646_ tms1x00.RAM\[44\]\[2\] tms1x00.RAM\[45\]\[2\] tms1x00.RAM\[46\]\[2\] tms1x00.RAM\[47\]\[2\]
+ _0955_ _0956_ vssd1 vssd1 vccd1 vccd1 _1037_ sky130_fd_sc_hd__mux4_2
X_2577_ _0944_ _0962_ _0964_ _0821_ _0968_ vssd1 vssd1 vccd1 vccd1 _0969_ sky130_fd_sc_hd__a311o_1
XFILLER_59_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4316_ _2138_ vssd1 vssd1 vccd1 vccd1 _0621_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4474__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4247_ tms1x00.A\[3\] _2082_ _2096_ vssd1 vssd1 vccd1 vccd1 _2100_ sky130_fd_sc_hd__mux2_1
X_4178_ _0760_ _2046_ _2047_ _1966_ vssd1 vssd1 vccd1 vccd1 _0574_ sky130_fd_sc_hd__o211a_1
XFILLER_28_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3898__A _1257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3129_ _1412_ vssd1 vssd1 vccd1 vccd1 _0160_ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2408__A2 tms1x00.RAM\[90\]\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3605__A1 _1676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2307__A net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4817__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2977__A _0914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4097__A1 tms1x00.PC\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4967__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2916__S _0715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2280__B1 _0703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3048__A _1034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3780__A0 _1706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2500_ tms1x00.RAM\[60\]\[0\] tms1x00.RAM\[61\]\[0\] tms1x00.RAM\[62\]\[0\] tms1x00.RAM\[63\]\[0\]
+ _0777_ _0779_ vssd1 vssd1 vccd1 vccd1 _0893_ sky130_fd_sc_hd__mux4_1
XFILLER_6_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3480_ tms1x00.RAM\[42\]\[1\] _1574_ _1614_ vssd1 vssd1 vccd1 vccd1 _1616_ sky130_fd_sc_hd__mux2_1
XFILLER_6_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2431_ tms1x00.RAM\[70\]\[0\] tms1x00.RAM\[71\]\[0\] _0823_ vssd1 vssd1 vccd1 vccd1
+ _0824_ sky130_fd_sc_hd__mux2_1
X_2362_ _0744_ tms1x00.ins_in\[1\] _0742_ vssd1 vssd1 vccd1 vccd1 _0757_ sky130_fd_sc_hd__or3b_1
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4101_ _0762_ _0745_ vssd1 vssd1 vccd1 vccd1 _1986_ sky130_fd_sc_hd__nor2_1
X_2293_ _0706_ vssd1 vssd1 vccd1 vccd1 _0020_ sky130_fd_sc_hd__clkbuf_1
X_4032_ _1938_ vssd1 vssd1 vccd1 vccd1 _0537_ sky130_fd_sc_hd__clkbuf_1
XFILLER_38_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_1__f_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_2_1__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_37_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4934_ clknet_leaf_14_wb_clk_i _0544_ vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__dfxtp_2
XFILLER_24_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_19_wb_clk_i clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_32_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4865_ clknet_leaf_21_wb_clk_i _0479_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[88\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_3816_ tms1x00.RAM\[85\]\[1\] _1775_ _1806_ vssd1 vssd1 vccd1 vccd1 _1808_ sky130_fd_sc_hd__mux2_1
X_4796_ clknet_leaf_25_wb_clk_i _0410_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[70\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_13_wb_clk_i_A clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_20_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3747_ tms1x00.RAM\[75\]\[0\] _1669_ _1767_ vssd1 vssd1 vccd1 vccd1 _1768_ sky130_fd_sc_hd__mux2_1
XFILLER_21_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3678_ _1729_ vssd1 vssd1 vccd1 vccd1 _0392_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__3523__A0 _1585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput141 net141 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[3] sky130_fd_sc_hd__buf_2
Xoutput130 net130 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[22] sky130_fd_sc_hd__buf_2
XFILLER_0_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2797__A _0927_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2629_ tms1x00.RAM\[55\]\[1\] _0873_ vssd1 vssd1 vccd1 vccd1 _1021_ sky130_fd_sc_hd__or2b_1
XFILLER_75_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4236__B _2007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2471__S _0826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2660__S1 _0822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input61_A wbs_dat_i[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3514__A0 _1585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2980_ tms1x00.RAM\[102\]\[1\] _1243_ _1318_ vssd1 vssd1 vccd1 vccd1 _1320_ sky130_fd_sc_hd__mux2_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4650_ clknet_leaf_5_wb_clk_i _0271_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[34\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput21 ram_val[16] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_1
X_3601_ tms1x00.RAM\[56\]\[1\] _1672_ _1683_ vssd1 vssd1 vccd1 vccd1 _1685_ sky130_fd_sc_hd__mux2_1
Xinput10 oram_value[4] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_1
X_4581_ clknet_leaf_2_wb_clk_i _0202_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[118\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput54 wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__clkbuf_1
Xinput32 ram_val[26] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__clkbuf_1
Xinput43 ram_val[7] vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__clkbuf_2
Xinput65 wbs_dat_i[8] vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2651__S1 _0800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3532_ tms1x00.RAM\[54\]\[0\] _1571_ _1644_ vssd1 vssd1 vccd1 vccd1 _1645_ sky130_fd_sc_hd__mux2_1
X_3463_ _1606_ vssd1 vssd1 vccd1 vccd1 _0300_ sky130_fd_sc_hd__clkbuf_1
XFILLER_69_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3505__A0 _1585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2414_ _0797_ vssd1 vssd1 vccd1 vccd1 _0807_ sky130_fd_sc_hd__clkbuf_4
X_3394_ _1564_ vssd1 vssd1 vccd1 vccd1 _0273_ sky130_fd_sc_hd__clkbuf_1
XFILLER_69_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2345_ tms1x00.Y\[1\] tms1x00.Y\[0\] vssd1 vssd1 vccd1 vccd1 _0740_ sky130_fd_sc_hd__nor2_1
X_2276_ net80 _0702_ _0703_ wbs_o_buff\[11\] vssd1 vssd1 vccd1 vccd1 _0005_ sky130_fd_sc_hd__a22o_1
X_4015_ net80 _1924_ _1925_ _1901_ vssd1 vssd1 vccd1 vccd1 _0533_ sky130_fd_sc_hd__o211a_1
XANTENNA__4512__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4917_ clknet_leaf_8_wb_clk_i tms1x00.K_in\[0\] vssd1 vssd1 vccd1 vccd1 tms1x00.K_latch\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2244__A0 net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4662__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4848_ clknet_leaf_16_wb_clk_i _0462_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[83\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2795__B2 _0922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4222__D _0742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3744__A0 _1710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4779_ clknet_leaf_18_wb_clk_i _0393_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[65\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2304__B _0699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5018__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3416__A _1224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2633__S1 _0780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3045__B _1345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3760__S _1773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2710__B2 _0786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4685__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2474__B1 _0866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2226__A0 net27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2963_ _1308_ vssd1 vssd1 vccd1 vccd1 _0098_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__3974__A0 tms1x00.ins_in\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4702_ clknet_leaf_29_wb_clk_i _0316_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[4\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2777__B2 _0787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2894_ _0717_ _0728_ _0916_ vssd1 vssd1 vccd1 vccd1 _1267_ sky130_fd_sc_hd__nand3_4
X_4633_ clknet_leaf_10_wb_clk_i _0254_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[30\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4564_ clknet_leaf_33_wb_clk_i _0185_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[122\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_3515_ _1635_ vssd1 vssd1 vccd1 vccd1 _0323_ sky130_fd_sc_hd__clkbuf_1
X_4495_ clknet_leaf_11_wb_clk_i _0116_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[0\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2388__S0 _0778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3446_ tms1x00.RAM\[38\]\[2\] _1576_ _1594_ vssd1 vssd1 vccd1 vccd1 _1597_ sky130_fd_sc_hd__mux2_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3377_ tms1x00.RAM\[36\]\[3\] _1463_ _1551_ vssd1 vssd1 vccd1 vccd1 _1555_ sky130_fd_sc_hd__mux2_1
XFILLER_69_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2328_ tms1x00.Y\[2\] vssd1 vssd1 vccd1 vccd1 _0730_ sky130_fd_sc_hd__buf_2
XFILLER_57_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_34_wb_clk_i clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_34_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_2259_ _0697_ vssd1 vssd1 vccd1 vccd1 _0698_ sky130_fd_sc_hd__buf_2
XFILLER_26_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2315__A net76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapped_tms1x00_173 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_173/HI io_oeb[34] sky130_fd_sc_hd__conb_1
Xwrapped_tms1x00_162 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_162/HI io_oeb[23] sky130_fd_sc_hd__conb_1
Xwrapped_tms1x00_151 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_151/HI io_oeb[12] sky130_fd_sc_hd__conb_1
XANTENNA__4408__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapped_tms1x00_184 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_184/HI io_out[7] sky130_fd_sc_hd__conb_1
Xwrapped_tms1x00_195 vssd1 vssd1 vccd1 vccd1 io_oeb[5] wrapped_tms1x00_195/LO sky130_fd_sc_hd__conb_1
XFILLER_5_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4558__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input24_A ram_val[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3956__A0 _0730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output92_A net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4381__A0 tms1x00.PC\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3300_ _1511_ vssd1 vssd1 vccd1 vccd1 _0232_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__2931__A1 _1245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4280_ _2118_ vssd1 vssd1 vccd1 vccd1 _0605_ sky130_fd_sc_hd__clkbuf_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2895__A _1237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3231_ _1471_ vssd1 vssd1 vccd1 vccd1 _0203_ sky130_fd_sc_hd__clkbuf_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3162_ _1430_ _1409_ vssd1 vssd1 vccd1 vccd1 _1431_ sky130_fd_sc_hd__or2_2
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3093_ _1390_ vssd1 vssd1 vccd1 vccd1 _0146_ sky130_fd_sc_hd__clkbuf_1
XFILLER_81_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3995_ _0718_ _1909_ _1910_ vssd1 vssd1 vccd1 vccd1 _1911_ sky130_fd_sc_hd__and3_1
XFILLER_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2946_ _1298_ vssd1 vssd1 vccd1 vccd1 _0091_ sky130_fd_sc_hd__clkbuf_1
X_2877_ _1255_ vssd1 vssd1 vccd1 vccd1 _0065_ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4616_ clknet_leaf_4_wb_clk_i _0237_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[27\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4700__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4547_ clknet_leaf_31_wb_clk_i _0168_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[106\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_4478_ clknet_leaf_30_wb_clk_i _0099_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[103\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4850__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3429_ _1229_ _1343_ vssd1 vssd1 vccd1 vccd1 _1586_ sky130_fd_sc_hd__or2_2
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2781__S0 _0823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2989__A1 _1324_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4051__C1 _1931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3780_ _1706_ tms1x00.RAM\[80\]\[1\] _1786_ vssd1 vssd1 vccd1 vccd1 _1788_ sky130_fd_sc_hd__mux2_1
X_2800_ tms1x00.RAM\[0\]\[3\] tms1x00.RAM\[1\]\[3\] tms1x00.RAM\[2\]\[3\] tms1x00.RAM\[3\]\[3\]
+ _0816_ _0977_ vssd1 vssd1 vccd1 vccd1 _1190_ sky130_fd_sc_hd__mux4_2
XFILLER_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2731_ _0783_ _1121_ vssd1 vssd1 vccd1 vccd1 _1122_ sky130_fd_sc_hd__or2_1
XFILLER_9_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2662_ _0797_ _1052_ vssd1 vssd1 vccd1 vccd1 _1053_ sky130_fd_sc_hd__or2_1
XANTENNA__3157__A1 _1331_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4401_ clknet_leaf_35_wb_clk_i _0030_ vssd1 vssd1 vccd1 vccd1 wbs_o_buff\[5\] sky130_fd_sc_hd__dfxtp_1
X_2593_ tms1x00.RAM\[20\]\[1\] tms1x00.RAM\[21\]\[1\] tms1x00.RAM\[22\]\[1\] tms1x00.RAM\[23\]\[1\]
+ _0975_ _0791_ vssd1 vssd1 vccd1 vccd1 _0985_ sky130_fd_sc_hd__mux4_2
X_4332_ _2147_ vssd1 vssd1 vccd1 vccd1 _0628_ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4263_ tms1x00.RAM\[39\]\[2\] _1330_ _2106_ vssd1 vssd1 vccd1 vccd1 _2109_ sky130_fd_sc_hd__mux2_1
X_3214_ _1330_ vssd1 vssd1 vccd1 vccd1 _1461_ sky130_fd_sc_hd__clkbuf_4
X_4194_ _2059_ _2060_ vssd1 vssd1 vccd1 vccd1 _2061_ sky130_fd_sc_hd__and2_1
XFILLER_39_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3145_ _1421_ vssd1 vssd1 vccd1 vccd1 _0167_ sky130_fd_sc_hd__clkbuf_1
XFILLER_54_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3076_ _1251_ _1375_ vssd1 vssd1 vccd1 vccd1 _1381_ sky130_fd_sc_hd__or2_2
XFILLER_36_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3978_ net8 _1899_ vssd1 vssd1 vccd1 vccd1 _1900_ sky130_fd_sc_hd__or2_1
XFILLER_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2929_ tms1x00.RAM\[59\]\[1\] _1243_ _1287_ vssd1 vssd1 vccd1 vccd1 _1289_ sky130_fd_sc_hd__mux2_1
XANTENNA__3148__A1 _1331_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3143__B _1403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2506__S0 _0815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4896__CLK clknet_leaf_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3139__A1 _1331_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2898__A0 _1035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3334__A _1249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput8 oram_value[2] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_1
Xclkbuf_2_0__f_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_2_0__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_36_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4950_ clknet_leaf_5_wb_clk_i _0560_ vssd1 vssd1 vccd1 vccd1 tms1x00.PB\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_33_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3901_ _1819_ tms1x00.RAM\[94\]\[1\] _1855_ vssd1 vssd1 vccd1 vccd1 _1857_ sky130_fd_sc_hd__mux2_1
X_4881_ clknet_leaf_17_wb_clk_i _0495_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[92\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_3832_ _1229_ _1257_ vssd1 vssd1 vccd1 vccd1 _1817_ sky130_fd_sc_hd__or2_2
XFILLER_20_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3763_ tms1x00.RAM\[74\]\[2\] _1777_ _1773_ vssd1 vssd1 vccd1 vccd1 _1778_ sky130_fd_sc_hd__mux2_1
X_2714_ tms1x00.RAM\[119\]\[2\] _0945_ vssd1 vssd1 vccd1 vccd1 _1105_ sky130_fd_sc_hd__or2b_1
X_3694_ _1738_ vssd1 vssd1 vccd1 vccd1 _0399_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__2413__A _0038_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2645_ _1036_ vssd1 vssd1 vccd1 vccd1 _0052_ sky130_fd_sc_hd__clkbuf_1
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4315_ _1819_ tms1x00.RAM\[12\]\[1\] _2136_ vssd1 vssd1 vccd1 vccd1 _2138_ sky130_fd_sc_hd__mux2_1
X_2576_ _0940_ _0965_ _0967_ _0942_ vssd1 vssd1 vccd1 vccd1 _0968_ sky130_fd_sc_hd__o211a_1
XFILLER_0_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3550__A1 _1571_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4619__CLK clknet_leaf_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4059__B _0768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4246_ _2099_ vssd1 vssd1 vccd1 vccd1 _0590_ sky130_fd_sc_hd__clkbuf_1
XFILLER_74_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4177_ tms1x00.PC\[3\] _1908_ vssd1 vssd1 vccd1 vccd1 _2047_ sky130_fd_sc_hd__or2_1
XFILLER_28_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3898__B _1396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3128_ _1364_ tms1x00.RAM\[108\]\[1\] _1410_ vssd1 vssd1 vccd1 vccd1 _1412_ sky130_fd_sc_hd__mux2_1
XFILLER_56_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3059_ _1371_ vssd1 vssd1 vccd1 vccd1 _0131_ sky130_fd_sc_hd__clkbuf_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4015__C1 _1901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3419__A _1303_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2977__B _1317_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3541__A1 _1571_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2469__S _0823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2727__S0 _0873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2804__B1 _0780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2280__A1 net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2430_ _0035_ vssd1 vssd1 vccd1 vccd1 _0823_ sky130_fd_sc_hd__buf_6
XANTENNA__3763__S _1773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3532__A1 _1571_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2361_ _0739_ _0740_ vssd1 vssd1 vccd1 vccd1 _0756_ sky130_fd_sc_hd__and2_1
XFILLER_69_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4100_ _1985_ vssd1 vssd1 vccd1 vccd1 _0558_ sky130_fd_sc_hd__clkbuf_1
X_2292_ wbs_o_buff\[25\] _0704_ vssd1 vssd1 vccd1 vccd1 _0706_ sky130_fd_sc_hd__and2_1
XANTENNA__2718__S0 _0873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4031_ _0718_ _1936_ _1937_ vssd1 vssd1 vccd1 vccd1 _1938_ sky130_fd_sc_hd__and3_1
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4933_ clknet_leaf_14_wb_clk_i _0543_ vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__dfxtp_2
XFILLER_52_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3599__A1 _1669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4864_ clknet_leaf_29_wb_clk_i _0478_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[8\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2271__A1 net77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2271__B2 wbs_o_buff\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3815_ _1807_ vssd1 vssd1 vccd1 vccd1 _0451_ sky130_fd_sc_hd__clkbuf_1
X_4795_ clknet_leaf_24_wb_clk_i _0409_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[70\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_3746_ _1237_ _1286_ vssd1 vssd1 vccd1 vccd1 _1767_ sky130_fd_sc_hd__nor2_2
XANTENNA__4441__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3771__A1 _1775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3677_ _1706_ tms1x00.RAM\[65\]\[1\] _1727_ vssd1 vssd1 vccd1 vccd1 _1729_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_9_wb_clk_i_A clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_2628_ _0794_ _1019_ _0038_ vssd1 vssd1 vccd1 vccd1 _1020_ sky130_fd_sc_hd__o21a_1
Xoutput142 net142 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[4] sky130_fd_sc_hd__buf_2
Xoutput120 net120 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[13] sky130_fd_sc_hd__buf_2
Xoutput131 net131 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[23] sky130_fd_sc_hd__buf_2
X_2559_ _0818_ _0950_ vssd1 vssd1 vccd1 vccd1 _0951_ sky130_fd_sc_hd__and2_1
X_4229_ tms1x00.X\[1\] _2088_ _2090_ _0766_ vssd1 vssd1 vccd1 vccd1 _0582_ sky130_fd_sc_hd__o211a_1
XFILLER_75_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2318__A net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2752__S _0823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2262__A1 net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2565__A2 tms1x00.RAM\[90\]\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2988__A _0914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input54_A wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4227__C1 _1966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2789__C1 _0944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4464__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4580_ clknet_leaf_1_wb_clk_i _0201_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[118\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput22 ram_val[17] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__clkbuf_1
X_3600_ _1684_ vssd1 vssd1 vccd1 vccd1 _0359_ sky130_fd_sc_hd__clkbuf_1
Xinput11 oram_value[5] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_1
Xinput55 wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__clkbuf_1
Xinput33 ram_val[27] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_1
Xinput44 ram_val[8] vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__clkbuf_2
XANTENNA__3753__A1 _1676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3531_ _1284_ _1317_ vssd1 vssd1 vccd1 vccd1 _1644_ sky130_fd_sc_hd__nor2_2
Xinput66 wbs_dat_i[9] vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__clkbuf_1
X_3462_ _1588_ tms1x00.RAM\[44\]\[1\] _1604_ vssd1 vssd1 vccd1 vccd1 _1606_ sky130_fd_sc_hd__mux2_1
XFILLER_6_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3393_ _1490_ tms1x00.RAM\[34\]\[2\] _1561_ vssd1 vssd1 vccd1 vccd1 _1564_ sky130_fd_sc_hd__mux2_1
X_2413_ _0038_ vssd1 vssd1 vccd1 vccd1 _0806_ sky130_fd_sc_hd__clkbuf_4
XFILLER_69_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2344_ tms1x00.Y\[2\] vssd1 vssd1 vccd1 vccd1 _0739_ sky130_fd_sc_hd__clkinv_2
XANTENNA__2713__C1 _0773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3522__A _1396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2275_ net79 _0702_ _0703_ wbs_o_buff\[10\] vssd1 vssd1 vccd1 vccd1 _0004_ sky130_fd_sc_hd__a22o_1
X_4014_ _0732_ _0753_ _1922_ vssd1 vssd1 vccd1 vccd1 _1925_ sky130_fd_sc_hd__or3b_1
XFILLER_38_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4916_ clknet_leaf_7_wb_clk_i _0530_ vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__dfxtp_4
XFILLER_21_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4847_ clknet_leaf_16_wb_clk_i _0461_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[83\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4957__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4778_ clknet_leaf_18_wb_clk_i _0392_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[65\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3729_ tms1x00.RAM\[68\]\[0\] _1669_ _1757_ vssd1 vssd1 vccd1 vccd1 _1758_ sky130_fd_sc_hd__mux2_1
XFILLER_76_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3432__A _1034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3735__A1 _1676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3607__A _1284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2511__A _0747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_4_wb_clk_i clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_4_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2474__B2 _0798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4173__A tms1x00.PC\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2962_ tms1x00.RAM\[104\]\[3\] _1247_ _1304_ vssd1 vssd1 vccd1 vccd1 _1308_ sky130_fd_sc_hd__mux2_1
XFILLER_22_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3974__A1 net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4701_ clknet_leaf_27_wb_clk_i _0315_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[4\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_4632_ clknet_leaf_10_wb_clk_i _0253_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[30\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_2893_ _1266_ vssd1 vssd1 vccd1 vccd1 _0070_ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2654__B_N _0975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3726__A1 _1676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4563_ clknet_leaf_33_wb_clk_i _0184_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[122\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_4494_ clknet_leaf_10_wb_clk_i _0115_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[0\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_3514_ _1585_ tms1x00.RAM\[47\]\[0\] _1634_ vssd1 vssd1 vccd1 vccd1 _1635_ sky130_fd_sc_hd__mux2_1
X_3445_ _1596_ vssd1 vssd1 vccd1 vccd1 _0292_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__2388__S1 _0780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3376_ _1554_ vssd1 vssd1 vccd1 vccd1 _0265_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4348__A _0917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2327_ _0729_ vssd1 vssd1 vccd1 vccd1 _0043_ sky130_fd_sc_hd__clkbuf_1
XFILLER_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2258_ _0696_ vssd1 vssd1 vccd1 vccd1 _0697_ sky130_fd_sc_hd__buf_4
XFILLER_27_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2189_ _0661_ vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__clkbuf_1
XANTENNA__2465__A1 _0773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapped_tms1x00_163 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_163/HI io_oeb[24] sky130_fd_sc_hd__conb_1
Xwrapped_tms1x00_152 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_152/HI io_oeb[13] sky130_fd_sc_hd__conb_1
Xwrapped_tms1x00_174 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_174/HI io_oeb[35] sky130_fd_sc_hd__conb_1
Xwrapped_tms1x00_185 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_185/HI io_out[8] sky130_fd_sc_hd__conb_1
Xwrapped_tms1x00_196 vssd1 vssd1 vccd1 vccd1 io_oeb[6] wrapped_tms1x00_196/LO sky130_fd_sc_hd__conb_1
XFILLER_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3717__A1 _1676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4258__A _1310_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3162__A _1430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input17_A ram_val[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3956__A1 tms1x00.ram_addr_buff\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3708__A1 _1676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4502__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4381__A1 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output85_A net85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2895__B _1267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3230_ tms1x00.RAM\[117\]\[0\] _1456_ _1470_ vssd1 vssd1 vccd1 vccd1 _1471_ sky130_fd_sc_hd__mux2_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3161_ _1375_ vssd1 vssd1 vccd1 vccd1 _1430_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__4652__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3092_ _1368_ tms1x00.RAM\[112\]\[3\] _1386_ vssd1 vssd1 vccd1 vccd1 _1390_ sky130_fd_sc_hd__mux2_1
XFILLER_48_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5008__CLK clknet_leaf_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3994_ _0701_ _1908_ vssd1 vssd1 vccd1 vccd1 _1910_ sky130_fd_sc_hd__or2_1
XFILLER_50_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2945_ _0912_ tms1x00.RAM\[19\]\[0\] _1297_ vssd1 vssd1 vccd1 vccd1 _1298_ sky130_fd_sc_hd__mux2_1
XANTENNA__3946__S _1880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2876_ _1130_ tms1x00.RAM\[17\]\[2\] _1252_ vssd1 vssd1 vccd1 vccd1 _1255_ sky130_fd_sc_hd__mux2_1
XFILLER_31_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4615_ clknet_leaf_4_wb_clk_i _0236_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[27\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3247__A _1229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4546_ clknet_leaf_31_wb_clk_i _0167_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[106\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_4477_ clknet_leaf_31_wb_clk_i _0098_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[104\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_3428_ _0911_ vssd1 vssd1 vccd1 vccd1 _1585_ sky130_fd_sc_hd__buf_2
XFILLER_58_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4078__A net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3359_ _1492_ tms1x00.RAM\[2\]\[3\] _1541_ vssd1 vssd1 vccd1 vccd1 _1545_ sky130_fd_sc_hd__mux2_1
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input9_A oram_value[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2781__S1 _0850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5029_ clknet_leaf_22_wb_clk_i _0639_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[13\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3710__A _1237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4525__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2996__A _1330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3626__A0 _1585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3766__S _1773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2670__S _0923_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2601__A1 _0944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2730_ tms1x00.RAM\[104\]\[2\] tms1x00.RAM\[105\]\[2\] tms1x00.RAM\[106\]\[2\] tms1x00.RAM\[107\]\[2\]
+ _0823_ _0850_ vssd1 vssd1 vccd1 vccd1 _1121_ sky130_fd_sc_hd__mux4_1
XFILLER_9_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2661_ tms1x00.RAM\[56\]\[2\] tms1x00.RAM\[57\]\[2\] tms1x00.RAM\[58\]\[2\] tms1x00.RAM\[59\]\[2\]
+ _0815_ _0812_ vssd1 vssd1 vccd1 vccd1 _1052_ sky130_fd_sc_hd__mux4_1
XANTENNA__3067__A _1273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4400_ clknet_leaf_35_wb_clk_i _0029_ vssd1 vssd1 vccd1 vccd1 wbs_o_buff\[4\] sky130_fd_sc_hd__dfxtp_1
X_2592_ tms1x00.RAM\[16\]\[1\] tms1x00.RAM\[17\]\[1\] tms1x00.RAM\[18\]\[1\] tms1x00.RAM\[19\]\[1\]
+ _0975_ _0791_ vssd1 vssd1 vccd1 vccd1 _0984_ sky130_fd_sc_hd__mux4_1
X_4331_ _1235_ tms1x00.RAM\[15\]\[0\] _2146_ vssd1 vssd1 vccd1 vccd1 _2147_ sky130_fd_sc_hd__mux2_1
X_4262_ _2108_ vssd1 vssd1 vccd1 vccd1 _0597_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3213_ _1460_ vssd1 vssd1 vccd1 vccd1 _0196_ sky130_fd_sc_hd__clkbuf_1
XFILLER_79_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4193_ tms1x00.ins_in\[4\] _2058_ tms1x00.N\[0\] vssd1 vssd1 vccd1 vccd1 _2060_ sky130_fd_sc_hd__o21ai_1
XFILLER_28_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3144_ tms1x00.RAM\[106\]\[0\] _1324_ _1420_ vssd1 vssd1 vccd1 vccd1 _1421_ sky130_fd_sc_hd__mux2_1
XFILLER_82_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3075_ _1380_ vssd1 vssd1 vccd1 vccd1 _0138_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3617__A0 _1585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_32_wb_clk_i_A clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_63_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4548__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3977_ _0701_ _0760_ _0720_ vssd1 vssd1 vccd1 vccd1 _1899_ sky130_fd_sc_hd__or3b_1
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2928_ _1288_ vssd1 vssd1 vccd1 vccd1 _0083_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4698__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4080__B _0747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2859_ _1034_ vssd1 vssd1 vccd1 vccd1 _1243_ sky130_fd_sc_hd__buf_4
X_4529_ clknet_leaf_14_wb_clk_i _0150_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[111\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3856__A0 _1819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2506__S1 _0812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4281__A0 _1821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4033__B1 net85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2690__S0 _0931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3334__B _1267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3847__A0 _1819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput9 oram_value[3] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_1
XFILLER_80_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3900_ _1856_ vssd1 vssd1 vccd1 vccd1 _0487_ sky130_fd_sc_hd__clkbuf_1
X_4880_ clknet_leaf_17_wb_clk_i _0494_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[93\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2822__B2 _0787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3831_ _0911_ vssd1 vssd1 vccd1 vccd1 _1816_ sky130_fd_sc_hd__clkbuf_4
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3762_ _1129_ vssd1 vssd1 vccd1 vccd1 _1777_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__2586__B1 _0977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2713_ _0920_ _1084_ _1090_ _1103_ _0773_ vssd1 vssd1 vccd1 vccd1 _1104_ sky130_fd_sc_hd__o311a_1
X_3693_ tms1x00.RAM\[72\]\[0\] _1669_ _1737_ vssd1 vssd1 vccd1 vccd1 _1738_ sky130_fd_sc_hd__mux2_1
X_2644_ _1035_ tms1x00.RAM\[109\]\[1\] _0918_ vssd1 vssd1 vccd1 vccd1 _1036_ sky130_fd_sc_hd__mux2_1
XANTENNA__4990__CLK clknet_leaf_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2575_ _0798_ _0966_ vssd1 vssd1 vccd1 vccd1 _0967_ sky130_fd_sc_hd__or2_1
X_4314_ _2137_ vssd1 vssd1 vccd1 vccd1 _0620_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4059__C tms1x00.ins_in\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4245_ tms1x00.A\[2\] _2077_ _2096_ vssd1 vssd1 vccd1 vccd1 _2099_ sky130_fd_sc_hd__mux2_1
XFILLER_59_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4176_ _2043_ _2045_ vssd1 vssd1 vccd1 vccd1 _2046_ sky130_fd_sc_hd__xor2_1
XFILLER_56_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3127_ _1411_ vssd1 vssd1 vccd1 vccd1 _0159_ sky130_fd_sc_hd__clkbuf_1
XFILLER_56_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3260__A _1034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3058_ _1361_ tms1x00.RAM\[95\]\[0\] _1370_ vssd1 vssd1 vccd1 vccd1 _1371_ sky130_fd_sc_hd__mux2_1
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2307__C valid vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2604__A _0794_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2577__B1 _0821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3419__B _1525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2329__A0 _0730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3435__A _1129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2727__S1 _0822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4713__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2485__S _0826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2501__B1 _0038_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2804__A1 _0840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5097__A net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2568__B1 _0040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2740__A0 _1130_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2360_ _0754_ vssd1 vssd1 vccd1 vccd1 _0755_ sky130_fd_sc_hd__clkbuf_2
XFILLER_2_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2291_ _0705_ vssd1 vssd1 vccd1 vccd1 _0019_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__2718__S1 _0822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4030_ tms1x00.Y\[3\] _0752_ _1935_ vssd1 vssd1 vccd1 vccd1 _1937_ sky130_fd_sc_hd__or3b_1
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4932_ clknet_leaf_13_wb_clk_i _0542_ vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__dfxtp_2
XFILLER_61_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4863_ clknet_leaf_29_wb_clk_i _0477_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[8\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_3814_ tms1x00.RAM\[85\]\[0\] _1772_ _1806_ vssd1 vssd1 vccd1 vccd1 _1807_ sky130_fd_sc_hd__mux2_1
X_4794_ clknet_leaf_24_wb_clk_i _0408_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[70\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3954__S _0726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3745_ _1766_ vssd1 vssd1 vccd1 vccd1 _0422_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3676_ _1728_ vssd1 vssd1 vccd1 vccd1 _0391_ sky130_fd_sc_hd__clkbuf_1
Xoutput110 net110 vssd1 vssd1 vccd1 vccd1 ram_adrb[6] sky130_fd_sc_hd__buf_2
X_2627_ tms1x00.RAM\[60\]\[1\] tms1x00.RAM\[61\]\[1\] tms1x00.RAM\[62\]\[1\] tms1x00.RAM\[63\]\[1\]
+ _0826_ _0850_ vssd1 vssd1 vccd1 vccd1 _1019_ sky130_fd_sc_hd__mux4_1
Xoutput143 net143 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[5] sky130_fd_sc_hd__buf_2
Xoutput121 net121 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[14] sky130_fd_sc_hd__buf_2
Xoutput132 net132 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[24] sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_28_wb_clk_i clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_2558_ tms1x00.RAM\[92\]\[1\] tms1x00.RAM\[93\]\[1\] _0816_ vssd1 vssd1 vccd1 vccd1
+ _0950_ sky130_fd_sc_hd__mux2_1
XFILLER_0_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4736__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2489_ _0806_ _0870_ _0875_ _0039_ _0881_ vssd1 vssd1 vccd1 vccd1 _0882_ sky130_fd_sc_hd__a311o_1
X_4228_ tms1x00.X\[1\] _2087_ vssd1 vssd1 vccd1 vccd1 _2090_ sky130_fd_sc_hd__nand2_1
XANTENNA__4886__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4159_ _0719_ net75 _2029_ _2030_ _2031_ vssd1 vssd1 vccd1 vccd1 _2032_ sky130_fd_sc_hd__o32a_1
XFILLER_56_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2988__B _1240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4172__C1 _1966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input47_A wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5041__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4609__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput12 oram_value[6] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_1
X_3530_ _1643_ vssd1 vssd1 vccd1 vccd1 _0330_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4759__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput45 ram_val[9] vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__clkbuf_2
Xinput34 ram_val[28] vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__clkbuf_1
Xinput23 ram_val[18] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput67 wbs_stb_i vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__clkbuf_1
Xinput56 wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3461_ _1605_ vssd1 vssd1 vccd1 vccd1 _0299_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3392_ _1563_ vssd1 vssd1 vccd1 vccd1 _0272_ sky130_fd_sc_hd__clkbuf_1
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2412_ _0776_ _0784_ _0796_ _0803_ _0804_ vssd1 vssd1 vccd1 vccd1 _0805_ sky130_fd_sc_hd__a221o_1
X_2343_ net48 valid vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__nand2_1
XFILLER_69_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4013_ _1923_ vssd1 vssd1 vccd1 vccd1 _1924_ sky130_fd_sc_hd__inv_2
X_2274_ _0699_ vssd1 vssd1 vccd1 vccd1 _0703_ sky130_fd_sc_hd__clkbuf_4
XFILLER_38_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4915_ clknet_leaf_8_wb_clk_i _0529_ vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__dfxtp_4
XFILLER_21_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4846_ clknet_leaf_16_wb_clk_i _0460_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[83\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4777_ clknet_leaf_19_wb_clk_i _0391_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[65\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2627__S0 _0826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3728_ _1237_ _1337_ vssd1 vssd1 vccd1 vccd1 _1757_ sky130_fd_sc_hd__nor2_2
X_3659_ _1706_ tms1x00.RAM\[67\]\[1\] _1717_ vssd1 vssd1 vccd1 vccd1 _1719_ sky130_fd_sc_hd__mux2_1
XFILLER_57_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4901__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2618__S0 _0808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2456__B_N _0808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_3__f_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3607__B _1310_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2961_ _1307_ vssd1 vssd1 vccd1 vccd1 _0097_ sky130_fd_sc_hd__clkbuf_1
XFILLER_15_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4700_ clknet_leaf_3_wb_clk_i _0314_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[50\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4581__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4631_ clknet_leaf_10_wb_clk_i _0252_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[30\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_2892_ tms1x00.RAM\[89\]\[3\] _1247_ _1262_ vssd1 vssd1 vccd1 vccd1 _1266_ sky130_fd_sc_hd__mux2_1
XFILLER_30_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4562_ clknet_leaf_33_wb_clk_i _0183_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[122\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_3513_ _1267_ _1524_ vssd1 vssd1 vccd1 vccd1 _1634_ sky130_fd_sc_hd__or2_2
X_4493_ clknet_leaf_30_wb_clk_i _0114_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[100\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_3444_ tms1x00.RAM\[38\]\[1\] _1574_ _1594_ vssd1 vssd1 vccd1 vccd1 _1596_ sky130_fd_sc_hd__mux2_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3375_ tms1x00.RAM\[36\]\[2\] _1461_ _1551_ vssd1 vssd1 vccd1 vccd1 _1554_ sky130_fd_sc_hd__mux2_1
XANTENNA__4348__B _1343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2326_ tms1x00.Y\[1\] _0728_ _0726_ vssd1 vssd1 vccd1 vccd1 _0729_ sky130_fd_sc_hd__mux2_1
XFILLER_73_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5045_ clknet_leaf_4_wb_clk_i _0655_ vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__dfxtp_1
X_2257_ net49 net114 valid vssd1 vssd1 vccd1 vccd1 _0696_ sky130_fd_sc_hd__and3_1
XANTENNA__3111__A0 _1368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2188_ net39 wbs_o_buff\[3\] _0657_ vssd1 vssd1 vccd1 vccd1 _0661_ sky130_fd_sc_hd__mux2_1
XFILLER_25_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3414__A1 _1576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapped_tms1x00_164 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_164/HI io_oeb[25] sky130_fd_sc_hd__conb_1
Xwrapped_tms1x00_153 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_153/HI io_oeb[14] sky130_fd_sc_hd__conb_1
X_4829_ clknet_leaf_20_wb_clk_i _0443_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[78\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xwrapped_tms1x00_175 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_175/HI io_oeb[36] sky130_fd_sc_hd__conb_1
Xwrapped_tms1x00_186 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_186/HI io_out[9] sky130_fd_sc_hd__conb_1
Xwrapped_tms1x00_197 vssd1 vssd1 vccd1 vccd1 io_oeb[7] wrapped_tms1x00_197/LO sky130_fd_sc_hd__conb_1
XFILLER_4_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4142__A2 _2007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3350__A0 _1492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2689__C1 _0773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4258__B _1525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3162__B _1409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4454__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3169__A0 _1368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2916__A0 K_override\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output78_A net78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3341__A0 _1492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3160_ _1429_ vssd1 vssd1 vccd1 vccd1 _0174_ sky130_fd_sc_hd__clkbuf_1
XFILLER_66_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3091_ _1389_ vssd1 vssd1 vccd1 vccd1 _0145_ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1 feedback_delay vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3892__A1 _1775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_22_wb_clk_i_A clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_81_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3993_ _0701_ _1908_ vssd1 vssd1 vccd1 vccd1 _1909_ sky130_fd_sc_hd__nand2_1
XFILLER_16_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2944_ _1229_ _1249_ vssd1 vssd1 vccd1 vccd1 _1297_ sky130_fd_sc_hd__or2_2
XFILLER_31_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2875_ _1254_ vssd1 vssd1 vccd1 vccd1 _0064_ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4614_ clknet_leaf_0_wb_clk_i _0235_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[27\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2432__A _0822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3247__B _1375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4545_ clknet_leaf_31_wb_clk_i _0166_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[107\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_4476_ clknet_leaf_31_wb_clk_i _0097_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[104\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4477__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3263__A _1129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3332__A0 _1492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3427_ _1584_ vssd1 vssd1 vccd1 vccd1 _0286_ sky130_fd_sc_hd__clkbuf_1
X_3358_ _1544_ vssd1 vssd1 vccd1 vccd1 _0257_ sky130_fd_sc_hd__clkbuf_1
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2309_ net59 _0715_ vssd1 vssd1 vccd1 vccd1 _0716_ sky130_fd_sc_hd__and2_1
XANTENNA__3883__A1 _1775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3289_ _1505_ vssd1 vssd1 vccd1 vccd1 _0227_ sky130_fd_sc_hd__clkbuf_1
X_5028_ clknet_leaf_19_wb_clk_i _0638_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[13\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_54_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3710__B _1317_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3438__A _1224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2342__A _0738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3874__A1 _1775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4051__A1 net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2660_ tms1x00.RAM\[60\]\[2\] tms1x00.RAM\[61\]\[2\] tms1x00.RAM\[62\]\[2\] tms1x00.RAM\[63\]\[2\]
+ _0840_ _0822_ vssd1 vssd1 vccd1 vccd1 _1051_ sky130_fd_sc_hd__mux4_1
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3067__B _1375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2591_ _0969_ _0982_ _0835_ vssd1 vssd1 vccd1 vccd1 _0983_ sky130_fd_sc_hd__a21oi_1
X_4330_ _1267_ _1343_ vssd1 vssd1 vccd1 vccd1 _2146_ sky130_fd_sc_hd__or2_2
XANTENNA__4179__A tms1x00.PC\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4261_ tms1x00.RAM\[39\]\[1\] _1327_ _2106_ vssd1 vssd1 vccd1 vccd1 _2108_ sky130_fd_sc_hd__mux2_1
XFILLER_68_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3212_ tms1x00.RAM\[11\]\[1\] _1459_ _1457_ vssd1 vssd1 vccd1 vccd1 _1460_ sky130_fd_sc_hd__mux2_1
XFILLER_79_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4192_ tms1x00.ins_in\[4\] tms1x00.N\[0\] _2058_ vssd1 vssd1 vccd1 vccd1 _2059_ sky130_fd_sc_hd__or3_1
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3865__A1 _1775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3143_ _0914_ _1403_ vssd1 vssd1 vccd1 vccd1 _1420_ sky130_fd_sc_hd__nor2_2
XFILLER_67_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3074_ _1368_ tms1x00.RAM\[114\]\[3\] _1376_ vssd1 vssd1 vccd1 vccd1 _1380_ sky130_fd_sc_hd__mux2_1
XFILLER_36_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3617__A1 tms1x00.RAM\[63\]\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4290__A1 _1330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3976_ _1898_ vssd1 vssd1 vccd1 vccd1 _0521_ sky130_fd_sc_hd__clkbuf_1
XFILLER_50_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2927_ tms1x00.RAM\[59\]\[0\] _1235_ _1287_ vssd1 vssd1 vccd1 vccd1 _1288_ sky130_fd_sc_hd__mux2_1
XFILLER_31_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4080__C _0748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2858_ _1242_ vssd1 vssd1 vccd1 vccd1 _0059_ sky130_fd_sc_hd__clkbuf_1
X_2789_ _0922_ _1176_ _1178_ _0944_ vssd1 vssd1 vccd1 vccd1 _1179_ sky130_fd_sc_hd__o211a_1
X_4528_ clknet_leaf_14_wb_clk_i _0149_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[111\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_49_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4459_ clknet_leaf_33_wb_clk_i _0080_ vssd1 vssd1 vccd1 vccd1 K_override\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_58_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3608__A1 _1669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2831__A2 _1155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4642__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2690__S1 _0932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4272__A1 _1330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2807__C1 _0806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2283__B1 _0703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3830_ _1815_ vssd1 vssd1 vccd1 vccd1 _0458_ sky130_fd_sc_hd__clkbuf_1
XFILLER_60_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3761_ _1776_ vssd1 vssd1 vccd1 vccd1 _0428_ sky130_fd_sc_hd__clkbuf_1
X_2712_ _0821_ _1096_ _1102_ vssd1 vssd1 vccd1 vccd1 _1103_ sky130_fd_sc_hd__or3_1
XANTENNA__2586__A1 _0975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3692_ _1237_ _1303_ vssd1 vssd1 vccd1 vccd1 _1737_ sky130_fd_sc_hd__nor2_2
X_2643_ _1034_ vssd1 vssd1 vccd1 vccd1 _1035_ sky130_fd_sc_hd__clkbuf_4
X_2574_ tms1x00.RAM\[104\]\[1\] tms1x00.RAM\[105\]\[1\] tms1x00.RAM\[106\]\[1\] tms1x00.RAM\[107\]\[1\]
+ _0799_ _0813_ vssd1 vssd1 vccd1 vccd1 _0966_ sky130_fd_sc_hd__mux4_1
X_4313_ _1816_ tms1x00.RAM\[12\]\[0\] _2136_ vssd1 vssd1 vccd1 vccd1 _2137_ sky130_fd_sc_hd__mux2_1
X_4244_ _2098_ vssd1 vssd1 vccd1 vccd1 _0589_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4175_ tms1x00.PC\[3\] _2030_ _2044_ _1971_ vssd1 vssd1 vccd1 vccd1 _2045_ sky130_fd_sc_hd__o22a_1
XFILLER_68_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3126_ _1361_ tms1x00.RAM\[108\]\[0\] _1410_ vssd1 vssd1 vccd1 vccd1 _1411_ sky130_fd_sc_hd__mux2_1
XANTENNA__2510__A1 _0773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3057_ _1258_ _1267_ vssd1 vssd1 vccd1 vccd1 _1370_ sky130_fd_sc_hd__or2_2
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4263__A1 _1330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4015__A1 net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3959_ _1888_ vssd1 vssd1 vccd1 vccd1 _0514_ sky130_fd_sc_hd__clkbuf_1
XFILLER_51_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2577__A1 _0944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2329__A1 tms1x00.ram_addr_buff\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3829__A1 _1779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2501__A1 _0828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4254__A1 _1330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2568__A1 _0920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2530__A _0921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2290_ wbs_o_buff\[24\] _0704_ vssd1 vssd1 vccd1 vccd1 _0705_ sky130_fd_sc_hd__and2_1
XFILLER_49_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2676__S _0815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3361__A _1240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4688__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4931_ clknet_leaf_9_wb_clk_i _0541_ vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__dfxtp_2
XFILLER_45_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4192__A tms1x00.ins_in\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4862_ clknet_leaf_21_wb_clk_i _0476_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[8\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3813_ _1240_ _1258_ vssd1 vssd1 vccd1 vccd1 _1806_ sky130_fd_sc_hd__nor2_2
X_4793_ clknet_leaf_24_wb_clk_i _0407_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[70\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_3744_ _1710_ tms1x00.RAM\[76\]\[3\] _1762_ vssd1 vssd1 vccd1 vccd1 _1766_ sky130_fd_sc_hd__mux2_1
X_3675_ _1703_ tms1x00.RAM\[65\]\[0\] _1727_ vssd1 vssd1 vccd1 vccd1 _1728_ sky130_fd_sc_hd__mux2_1
X_2626_ _0783_ _1017_ vssd1 vssd1 vccd1 vccd1 _1018_ sky130_fd_sc_hd__or2_1
Xoutput100 net100 vssd1 vssd1 vccd1 vccd1 oram_addr[5] sky130_fd_sc_hd__buf_2
Xoutput111 net111 vssd1 vssd1 vccd1 vccd1 ram_adrb[7] sky130_fd_sc_hd__buf_2
Xoutput122 net122 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[15] sky130_fd_sc_hd__buf_2
Xoutput133 net133 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[25] sky130_fd_sc_hd__buf_2
X_2557_ _0946_ _0947_ _0948_ vssd1 vssd1 vccd1 vccd1 _0949_ sky130_fd_sc_hd__mux2_1
Xoutput144 net144 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[6] sky130_fd_sc_hd__buf_2
X_2488_ _0877_ _0879_ _0880_ _0807_ _0775_ vssd1 vssd1 vccd1 vccd1 _0881_ sky130_fd_sc_hd__o221a_1
XFILLER_68_550 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4227_ tms1x00.X\[0\] _2088_ _2089_ _1966_ vssd1 vssd1 vccd1 vccd1 _0581_ sky130_fd_sc_hd__o211a_1
XFILLER_56_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4158_ tms1x00.PC\[0\] vssd1 vssd1 vccd1 vccd1 _2031_ sky130_fd_sc_hd__inv_2
X_4089_ tms1x00.SR\[0\] tms1x00.PC\[0\] _1979_ vssd1 vssd1 vccd1 vccd1 _1980_ sky130_fd_sc_hd__mux2_1
X_3109_ _1366_ tms1x00.RAM\[110\]\[2\] _1397_ vssd1 vssd1 vccd1 vccd1 _1400_ sky130_fd_sc_hd__mux2_1
XFILLER_44_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4830__CLK clknet_leaf_20_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2486__B1 _0828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4980__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2238__A0 net33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2525__A _0914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2789__A1 _0922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3738__A0 _1703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput13 oram_value[7] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_1
Xinput35 ram_val[29] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__clkbuf_1
Xinput24 ram_val[19] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__clkbuf_1
Xinput46 wb_rst_i vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__clkbuf_4
XFILLER_7_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2410__B1 _0802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput57 wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__clkbuf_1
Xinput68 wbs_we_i vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3460_ _1585_ tms1x00.RAM\[44\]\[0\] _1604_ vssd1 vssd1 vccd1 vccd1 _1605_ sky130_fd_sc_hd__mux2_1
X_3391_ _1488_ tms1x00.RAM\[34\]\[1\] _1561_ vssd1 vssd1 vccd1 vccd1 _1563_ sky130_fd_sc_hd__mux2_1
X_2411_ _0039_ vssd1 vssd1 vccd1 vccd1 _0804_ sky130_fd_sc_hd__inv_2
XANTENNA__3910__A0 _1819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2342_ _0738_ vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__clkbuf_4
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2713__A1 _0920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4012_ _0754_ _0763_ _1922_ vssd1 vssd1 vccd1 vccd1 _1923_ sky130_fd_sc_hd__nand3_1
XFILLER_38_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2273_ _0697_ vssd1 vssd1 vccd1 vccd1 _0702_ sky130_fd_sc_hd__clkbuf_4
XFILLER_77_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4914_ clknet_leaf_8_wb_clk_i _0528_ vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__dfxtp_2
XFILLER_40_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4845_ clknet_leaf_18_wb_clk_i _0459_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[83\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4776_ clknet_leaf_19_wb_clk_i _0390_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[66\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4703__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2627__S1 _0850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3727_ _1756_ vssd1 vssd1 vccd1 vccd1 _0414_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__3266__A _1224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3658_ _1718_ vssd1 vssd1 vccd1 vccd1 _0383_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4853__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2609_ tms1x00.RAM\[14\]\[1\] tms1x00.RAM\[15\]\[1\] _0924_ vssd1 vssd1 vccd1 vccd1
+ _1001_ sky130_fd_sc_hd__mux2_1
X_3589_ _1261_ _1284_ vssd1 vssd1 vccd1 vccd1 _1678_ sky130_fd_sc_hd__nor2_2
XANTENNA__3901__A0 _1819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2468__A0 _0859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2345__A tms1x00.Y\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2618__S1 _0780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3196__A1 _1334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2511__C _0748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_12_wb_clk_i_A clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2554__S0 _0945_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3120__A1 _1331_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4726__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2960_ tms1x00.RAM\[104\]\[2\] _1245_ _1304_ vssd1 vssd1 vccd1 vccd1 _1307_ sky130_fd_sc_hd__mux2_1
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2891_ _1265_ vssd1 vssd1 vccd1 vccd1 _0069_ sky130_fd_sc_hd__clkbuf_1
X_4630_ clknet_leaf_10_wb_clk_i _0251_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[30\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3187__A1 _1334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4876__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4561_ clknet_leaf_33_wb_clk_i _0182_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[123\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_3512_ _1633_ vssd1 vssd1 vccd1 vccd1 _0322_ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4492_ clknet_leaf_29_wb_clk_i _0113_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[100\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_3443_ _1595_ vssd1 vssd1 vccd1 vccd1 _0291_ sky130_fd_sc_hd__clkbuf_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3374_ _1553_ vssd1 vssd1 vccd1 vccd1 _0264_ sky130_fd_sc_hd__clkbuf_1
XFILLER_57_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2325_ tms1x00.ram_addr_buff\[1\] vssd1 vssd1 vccd1 vccd1 _0728_ sky130_fd_sc_hd__clkbuf_4
X_5044_ clknet_leaf_6_wb_clk_i _0654_ vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__dfxtp_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2256_ net68 vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__clkinv_2
XFILLER_72_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2187_ _0660_ vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__clkbuf_1
XFILLER_81_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4828_ clknet_leaf_22_wb_clk_i _0442_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[7\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
Xwrapped_tms1x00_154 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_154/HI io_oeb[15] sky130_fd_sc_hd__conb_1
XANTENNA__4375__A0 tms1x00.PC\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3178__A1 _1334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapped_tms1x00_176 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_176/HI io_oeb[37] sky130_fd_sc_hd__conb_1
Xwrapped_tms1x00_187 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_187/HI io_out[34] sky130_fd_sc_hd__conb_1
Xwrapped_tms1x00_165 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_165/HI io_oeb[26] sky130_fd_sc_hd__conb_1
Xwrapped_tms1x00_198 vssd1 vssd1 vccd1 vccd1 io_oeb[8] wrapped_tms1x00_198/LO sky130_fd_sc_hd__conb_1
X_4759_ clknet_leaf_10_wb_clk_i _0373_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[62\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_12_wb_clk_i clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__5031__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4749__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4899__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3634__A _0911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3090_ _1366_ tms1x00.RAM\[112\]\[2\] _1386_ vssd1 vssd1 vccd1 vccd1 _1389_ sky130_fd_sc_hd__mux2_1
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4054__C1 _1931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3992_ _0722_ vssd1 vssd1 vccd1 vccd1 _1908_ sky130_fd_sc_hd__buf_2
XFILLER_23_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2943_ _1296_ vssd1 vssd1 vccd1 vccd1 _0090_ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2874_ _1035_ tms1x00.RAM\[17\]\[1\] _1252_ vssd1 vssd1 vccd1 vccd1 _1254_ sky130_fd_sc_hd__mux2_1
X_4613_ clknet_leaf_11_wb_clk_i _0234_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[28\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_4544_ clknet_leaf_31_wb_clk_i _0165_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[107\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_4475_ clknet_leaf_30_wb_clk_i _0096_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[104\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_3426_ tms1x00.RAM\[40\]\[3\] _1578_ _1580_ vssd1 vssd1 vccd1 vccd1 _1584_ sky130_fd_sc_hd__mux2_1
XANTENNA__2766__S0 _0931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3357_ _1490_ tms1x00.RAM\[2\]\[2\] _1541_ vssd1 vssd1 vccd1 vccd1 _1544_ sky130_fd_sc_hd__mux2_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2308_ net49 net68 valid vssd1 vssd1 vccd1 vccd1 _0715_ sky130_fd_sc_hd__and3_2
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5027_ clknet_leaf_20_wb_clk_i _0637_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[13\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2594__S _0921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3288_ tms1x00.RAM\[24\]\[0\] _1456_ _1504_ vssd1 vssd1 vccd1 vccd1 _1505_ sky130_fd_sc_hd__mux2_1
XFILLER_73_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2239_ _0687_ vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__clkbuf_1
XFILLER_72_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3719__A _1317_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3020__A0 _1035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input22_A ram_val[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4285__A _1240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output109_A net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output90_A net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2590_ _0920_ _0973_ _0981_ _0040_ vssd1 vssd1 vccd1 vccd1 _0982_ sky130_fd_sc_hd__o31a_1
XFILLER_4_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4914__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4260_ _2107_ vssd1 vssd1 vccd1 vccd1 _0596_ sky130_fd_sc_hd__clkbuf_1
X_4191_ _0748_ tms1x00.ins_in\[5\] _0747_ vssd1 vssd1 vccd1 vccd1 _2058_ sky130_fd_sc_hd__or3b_2
X_3211_ _1327_ vssd1 vssd1 vccd1 vccd1 _1459_ sky130_fd_sc_hd__buf_2
XFILLER_79_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3142_ _1419_ vssd1 vssd1 vccd1 vccd1 _0166_ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3073_ _1379_ vssd1 vssd1 vccd1 vccd1 _0137_ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4027__C1 _1931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3975_ net103 _1897_ vssd1 vssd1 vccd1 vccd1 _1898_ sky130_fd_sc_hd__or2_1
XANTENNA__2589__C1 _0776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3250__A0 _1364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2926_ _1284_ _1286_ vssd1 vssd1 vccd1 vccd1 _1287_ sky130_fd_sc_hd__nor2_2
XANTENNA__4444__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2857_ tms1x00.RAM\[69\]\[0\] _1235_ _1241_ vssd1 vssd1 vccd1 vccd1 _1242_ sky130_fd_sc_hd__mux2_1
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2788_ _0996_ _1177_ vssd1 vssd1 vccd1 vccd1 _1178_ sky130_fd_sc_hd__or2_1
XFILLER_3_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4151__A_N _0701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4527_ clknet_leaf_13_wb_clk_i _0148_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[111\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_49_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4458_ clknet_leaf_33_wb_clk_i _0079_ vssd1 vssd1 vccd1 vccd1 K_override\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_59_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3409_ _1573_ vssd1 vssd1 vccd1 vccd1 _0279_ sky130_fd_sc_hd__clkbuf_1
X_4389_ tms1x00.PA\[3\] net102 _2006_ vssd1 vssd1 vccd1 vccd1 _2178_ sky130_fd_sc_hd__mux2_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4018__C1 _1901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2528__A _0804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4009__C1 _1901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2283__A1 net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4467__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3760_ tms1x00.RAM\[74\]\[1\] _1775_ _1773_ vssd1 vssd1 vccd1 vccd1 _1776_ sky130_fd_sc_hd__mux2_1
X_2711_ _0921_ _1097_ _1101_ _0802_ vssd1 vssd1 vccd1 vccd1 _1102_ sky130_fd_sc_hd__o211a_1
XFILLER_13_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3691_ _1736_ vssd1 vssd1 vccd1 vccd1 _0398_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2642_ _1033_ vssd1 vssd1 vccd1 vccd1 _1034_ sky130_fd_sc_hd__buf_4
XANTENNA__3094__A _0913_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2573_ tms1x00.RAM\[108\]\[1\] tms1x00.RAM\[109\]\[1\] tms1x00.RAM\[110\]\[1\] tms1x00.RAM\[111\]\[1\]
+ _0955_ _0956_ vssd1 vssd1 vccd1 vccd1 _0965_ sky130_fd_sc_hd__mux4_1
X_4312_ _1344_ _1409_ vssd1 vssd1 vccd1 vccd1 _2136_ sky130_fd_sc_hd__or2_2
X_4243_ tms1x00.A\[1\] _2070_ _2096_ vssd1 vssd1 vccd1 vccd1 _2098_ sky130_fd_sc_hd__mux2_1
XANTENNA__3299__A0 _1488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3822__A _1258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4174_ tms1x00.ins_in\[5\] _1995_ _2027_ tms1x00.SR\[3\] vssd1 vssd1 vccd1 vccd1
+ _2044_ sky130_fd_sc_hd__o22a_1
XFILLER_56_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3125_ _0913_ _1409_ vssd1 vssd1 vccd1 vccd1 _1410_ sky130_fd_sc_hd__or2_2
XFILLER_55_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2438__A _0779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3056_ _1369_ vssd1 vssd1 vccd1 vccd1 _0130_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3968__S net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3269__A _0917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3958_ _0733_ tms1x00.ram_addr_buff\[3\] _0725_ vssd1 vssd1 vccd1 vccd1 _1888_ sky130_fd_sc_hd__mux2_1
X_2909_ _1276_ vssd1 vssd1 vccd1 vccd1 _0076_ sky130_fd_sc_hd__clkbuf_1
X_3889_ _1258_ _1310_ vssd1 vssd1 vccd1 vccd1 _1850_ sky130_fd_sc_hd__nor2_2
XFILLER_4_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3462__A0 _1588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2265__A1 net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2639__A_N _0747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3907__A _0917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2811__A _0996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3361__B _1525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4930_ clknet_leaf_9_wb_clk_i _0540_ vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__dfxtp_2
XANTENNA__3453__A0 _1588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4861_ clknet_leaf_29_wb_clk_i _0475_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[8\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_60_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3812_ _1805_ vssd1 vssd1 vccd1 vccd1 _0450_ sky130_fd_sc_hd__clkbuf_1
XFILLER_21_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4792_ clknet_leaf_25_wb_clk_i _0406_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[71\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3743_ _1765_ vssd1 vssd1 vccd1 vccd1 _0421_ sky130_fd_sc_hd__clkbuf_1
X_3674_ _1236_ _1251_ vssd1 vssd1 vccd1 vccd1 _1727_ sky130_fd_sc_hd__or2_2
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2625_ tms1x00.RAM\[56\]\[1\] tms1x00.RAM\[57\]\[1\] tms1x00.RAM\[58\]\[1\] tms1x00.RAM\[59\]\[1\]
+ _0823_ _0850_ vssd1 vssd1 vccd1 vccd1 _1017_ sky130_fd_sc_hd__mux4_1
Xoutput101 net101 vssd1 vssd1 vccd1 vccd1 oram_addr[6] sky130_fd_sc_hd__buf_2
XANTENNA__4181__A1 tms1x00.PC\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput112 net112 vssd1 vssd1 vccd1 vccd1 ram_adrb[8] sky130_fd_sc_hd__buf_2
Xoutput123 net123 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[16] sky130_fd_sc_hd__buf_2
Xoutput134 net134 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[26] sky130_fd_sc_hd__buf_2
X_2556_ _0783_ vssd1 vssd1 vccd1 vccd1 _0948_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__2192__A0 net41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput145 net145 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[7] sky130_fd_sc_hd__buf_2
X_2487_ tms1x00.RAM\[0\]\[0\] tms1x00.RAM\[1\]\[0\] tms1x00.RAM\[2\]\[0\] tms1x00.RAM\[3\]\[0\]
+ _0830_ _0831_ vssd1 vssd1 vccd1 vccd1 _0880_ sky130_fd_sc_hd__mux4_1
X_4226_ tms1x00.X\[0\] _2087_ vssd1 vssd1 vccd1 vccd1 _2089_ sky130_fd_sc_hd__nand2_1
XFILLER_29_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4157_ _1995_ _2027_ _1971_ vssd1 vssd1 vccd1 vccd1 _2030_ sky130_fd_sc_hd__a21oi_4
XFILLER_56_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4632__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3108_ _1399_ vssd1 vssd1 vccd1 vccd1 _0152_ sky130_fd_sc_hd__clkbuf_1
XFILLER_56_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4088_ tms1x00.CL _1978_ vssd1 vssd1 vccd1 vccd1 _1979_ sky130_fd_sc_hd__nor2_4
XFILLER_44_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3039_ _1358_ vssd1 vssd1 vccd1 vccd1 _0124_ sky130_fd_sc_hd__clkbuf_1
XFILLER_52_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3747__A1 _1669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2350__B net75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4172__A1 tms1x00.PC\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2486__A1 _0786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2525__B _0917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4505__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput25 ram_val[1] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_2
Xinput14 ram_val[0] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_2
Xinput36 ram_val[2] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2410__A1 _0798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput58 wbs_cyc_i vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__clkbuf_1
Xinput47 wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2410_ _0798_ _0801_ _0802_ vssd1 vssd1 vccd1 vccd1 _0803_ sky130_fd_sc_hd__o21a_1
XANTENNA__2260__B _0697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3390_ _1562_ vssd1 vssd1 vccd1 vccd1 _0271_ sky130_fd_sc_hd__clkbuf_1
XFILLER_69_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2341_ _0718_ vssd1 vssd1 vccd1 vccd1 _0738_ sky130_fd_sc_hd__clkinv_4
XANTENNA__4655__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2272_ net78 _0698_ _0700_ wbs_o_buff\[9\] vssd1 vssd1 vccd1 vccd1 _0034_ sky130_fd_sc_hd__a22o_1
X_4011_ tms1x00.Y\[2\] _1921_ vssd1 vssd1 vccd1 vccd1 _1922_ sky130_fd_sc_hd__nor2_1
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4913_ clknet_leaf_6_wb_clk_i _0527_ vssd1 vssd1 vccd1 vccd1 tms1x00.ins_in\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_34_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4844_ clknet_leaf_23_wb_clk_i _0458_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[84\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_4775_ clknet_leaf_18_wb_clk_i _0389_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[66\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3729__A1 _1669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3726_ tms1x00.RAM\[6\]\[3\] _1676_ _1752_ vssd1 vssd1 vccd1 vccd1 _1756_ sky130_fd_sc_hd__mux2_1
X_3657_ _1703_ tms1x00.RAM\[67\]\[0\] _1717_ vssd1 vssd1 vccd1 vccd1 _1718_ sky130_fd_sc_hd__mux2_1
X_2608_ _0948_ _0999_ _0776_ vssd1 vssd1 vccd1 vccd1 _1000_ sky130_fd_sc_hd__o21ai_1
X_3588_ _1677_ vssd1 vssd1 vccd1 vccd1 _0354_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__2597__S _0816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2539_ _0840_ vssd1 vssd1 vccd1 vccd1 _0931_ sky130_fd_sc_hd__buf_6
XFILLER_0_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4209_ tms1x00.P\[2\] tms1x00.N\[2\] vssd1 vssd1 vccd1 vccd1 _2074_ sky130_fd_sc_hd__nor2_1
XANTENNA__2468__A1 _0860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2626__A _0783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3968__A1 chip_sel_override vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2345__B tms1x00.Y\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4678__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4145__A1 _0730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input52_A wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2554__S1 _0791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2536__A _0927_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_8_wb_clk_i_A clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_35_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2890_ tms1x00.RAM\[89\]\[2\] _1245_ _1262_ vssd1 vssd1 vccd1 vccd1 _1265_ sky130_fd_sc_hd__mux2_1
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4560_ clknet_leaf_33_wb_clk_i _0181_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[123\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_3511_ _1592_ tms1x00.RAM\[48\]\[3\] _1629_ vssd1 vssd1 vccd1 vccd1 _1633_ sky130_fd_sc_hd__mux2_1
XANTENNA__2490__S0 _0808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4491_ clknet_leaf_30_wb_clk_i _0112_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[100\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4136__B2 tms1x00.Y\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3442_ tms1x00.RAM\[38\]\[0\] _1571_ _1594_ vssd1 vssd1 vccd1 vccd1 _1595_ sky130_fd_sc_hd__mux2_1
XANTENNA__4198__A _0766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3373_ tms1x00.RAM\[36\]\[1\] _1459_ _1551_ vssd1 vssd1 vccd1 vccd1 _1553_ sky130_fd_sc_hd__mux2_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2324_ _0727_ vssd1 vssd1 vccd1 vccd1 _0042_ sky130_fd_sc_hd__clkbuf_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3306__S _1514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2255_ _0695_ vssd1 vssd1 vccd1 vccd1 tms1x00.K_in\[3\] sky130_fd_sc_hd__clkbuf_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5043_ clknet_leaf_4_wb_clk_i _0653_ vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__dfxtp_1
XFILLER_66_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2186_ net36 wbs_o_buff\[2\] _0657_ vssd1 vssd1 vccd1 vccd1 _0660_ sky130_fd_sc_hd__mux2_1
XFILLER_81_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4827_ clknet_leaf_21_wb_clk_i _0441_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[7\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xwrapped_tms1x00_155 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_155/HI io_oeb[16] sky130_fd_sc_hd__conb_1
XANTENNA__4375__A1 net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2181__A net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4820__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwrapped_tms1x00_188 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_188/HI io_out[35] sky130_fd_sc_hd__conb_1
Xwrapped_tms1x00_166 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_166/HI io_oeb[27] sky130_fd_sc_hd__conb_1
Xwrapped_tms1x00_177 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_177/HI io_out[0] sky130_fd_sc_hd__conb_1
X_4758_ clknet_leaf_2_wb_clk_i _0372_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[62\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xwrapped_tms1x00_199 vssd1 vssd1 vccd1 vccd1 io_oeb[9] wrapped_tms1x00_199/LO sky130_fd_sc_hd__conb_1
X_4689_ clknet_leaf_32_wb_clk_i _0303_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[43\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3709_ _1746_ vssd1 vssd1 vccd1 vccd1 _0406_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4970__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2689__A1 _0920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2790__S _0945_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3991_ _0747_ _0724_ _1907_ _1901_ vssd1 vssd1 vccd1 vccd1 _0527_ sky130_fd_sc_hd__o211a_1
X_2942_ _1225_ tms1x00.RAM\[49\]\[3\] _1292_ vssd1 vssd1 vccd1 vccd1 _1296_ sky130_fd_sc_hd__mux2_1
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2873_ _1253_ vssd1 vssd1 vccd1 vccd1 _0063_ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4612_ clknet_leaf_11_wb_clk_i _0233_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[28\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2205__S _0668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4993__CLK clknet_leaf_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4543_ clknet_leaf_31_wb_clk_i _0164_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[107\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_4474_ clknet_leaf_31_wb_clk_i _0095_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[104\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_3425_ _1583_ vssd1 vssd1 vccd1 vccd1 _0285_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__2766__S1 _0932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3356_ _1543_ vssd1 vssd1 vccd1 vccd1 _0256_ sky130_fd_sc_hd__clkbuf_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3287_ _1250_ _1303_ vssd1 vssd1 vccd1 vccd1 _1504_ sky130_fd_sc_hd__nor2_2
X_2307_ net49 net68 valid vssd1 vssd1 vccd1 vccd1 _0714_ sky130_fd_sc_hd__nand3_2
XFILLER_39_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5026_ clknet_leaf_20_wb_clk_i _0636_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[13\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_2238_ net33 wbs_o_buff\[27\] _0679_ vssd1 vssd1 vccd1 vccd1 _0687_ sky130_fd_sc_hd__mux2_1
XFILLER_54_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3719__B _1344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2454__S0 _0815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4716__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4866__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input15_A ram_val[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4285__B _1250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4036__B1 net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2598__B1 _0819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output83_A net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4190_ _2055_ _2056_ _2057_ vssd1 vssd1 vccd1 vccd1 _0576_ sky130_fd_sc_hd__o21a_1
X_3210_ _1458_ vssd1 vssd1 vccd1 vccd1 _0195_ sky130_fd_sc_hd__clkbuf_1
XFILLER_79_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3141_ tms1x00.RAM\[107\]\[3\] _1334_ _1415_ vssd1 vssd1 vccd1 vccd1 _1419_ sky130_fd_sc_hd__mux2_1
XFILLER_67_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3072_ _1366_ tms1x00.RAM\[114\]\[2\] _1376_ vssd1 vssd1 vccd1 vccd1 _1379_ sky130_fd_sc_hd__mux2_1
XFILLER_54_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3974_ tms1x00.ins_in\[1\] net7 _0724_ vssd1 vssd1 vccd1 vccd1 _1897_ sky130_fd_sc_hd__mux2_1
XANTENNA__5100__A net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5021__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2925_ _1285_ vssd1 vssd1 vccd1 vccd1 _1286_ sky130_fd_sc_hd__buf_6
X_2856_ _1237_ _1240_ vssd1 vssd1 vccd1 vccd1 _1241_ sky130_fd_sc_hd__nor2_2
X_2787_ tms1x00.RAM\[20\]\[3\] tms1x00.RAM\[21\]\[3\] tms1x00.RAM\[22\]\[3\] tms1x00.RAM\[23\]\[3\]
+ _0923_ _0927_ vssd1 vssd1 vccd1 vccd1 _1177_ sky130_fd_sc_hd__mux4_2
X_4526_ clknet_leaf_13_wb_clk_i _0147_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[111\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4739__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4457_ clknet_leaf_12_wb_clk_i _0078_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[18\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_49_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3408_ tms1x00.RAM\[41\]\[0\] _1571_ _1572_ vssd1 vssd1 vccd1 vccd1 _1573_ sky130_fd_sc_hd__mux2_1
XFILLER_59_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4388_ _2177_ vssd1 vssd1 vccd1 vccd1 _0654_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_input7_A oram_value[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3339_ _1490_ tms1x00.RAM\[31\]\[2\] _1531_ vssd1 vssd1 vccd1 vccd1 _1534_ sky130_fd_sc_hd__mux2_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5009_ clknet_leaf_0_wb_clk_i _0619_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[20\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_27_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3241__A1 _1459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2807__A1 _0921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5044__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3480__A1 _1574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2666__S0 _0955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3232__A1 _1459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2710_ _1098_ _1099_ _1100_ _0786_ _0794_ vssd1 vssd1 vccd1 vccd1 _1101_ sky130_fd_sc_hd__a221o_1
XANTENNA__2440__C1 _0775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3690_ _1710_ tms1x00.RAM\[64\]\[3\] _1732_ vssd1 vssd1 vccd1 vccd1 _1736_ sky130_fd_sc_hd__mux2_1
X_2641_ _0771_ _1030_ _1032_ _0909_ tms1x00.A\[1\] vssd1 vssd1 vccd1 vccd1 _1033_
+ sky130_fd_sc_hd__a32o_1
XFILLER_9_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2572_ _0948_ _0963_ vssd1 vssd1 vccd1 vccd1 _0964_ sky130_fd_sc_hd__or2_1
XANTENNA__3094__B _1267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4311_ _2135_ vssd1 vssd1 vccd1 vccd1 _0619_ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4242_ _2097_ vssd1 vssd1 vccd1 vccd1 _0588_ sky130_fd_sc_hd__clkbuf_1
XFILLER_4_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3822__B _1337_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2719__A _0921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4173_ tms1x00.PC\[2\] tms1x00.PC\[1\] _2025_ vssd1 vssd1 vccd1 vccd1 _2043_ sky130_fd_sc_hd__and3_1
X_3124_ _0717_ _0728_ _0916_ vssd1 vssd1 vccd1 vccd1 _1409_ sky130_fd_sc_hd__or3b_4
X_3055_ _1368_ tms1x00.RAM\[96\]\[3\] _1362_ vssd1 vssd1 vccd1 vccd1 _1369_ sky130_fd_sc_hd__mux2_1
XFILLER_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3471__A1 _1574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3269__B _1375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3957_ _1887_ vssd1 vssd1 vccd1 vccd1 _0513_ sky130_fd_sc_hd__clkbuf_1
XFILLER_51_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3223__A1 _1459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2908_ _1035_ tms1x00.RAM\[18\]\[1\] _1274_ vssd1 vssd1 vccd1 vccd1 _1276_ sky130_fd_sc_hd__mux2_1
XFILLER_32_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3888_ _1849_ vssd1 vssd1 vccd1 vccd1 _0482_ sky130_fd_sc_hd__clkbuf_1
X_2839_ tms1x00.ram_addr_buff\[2\] tms1x00.ram_addr_buff\[3\] _0915_ vssd1 vssd1 vccd1
+ vccd1 _1228_ sky130_fd_sc_hd__or3_1
XANTENNA__4184__C1 _1966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4509_ clknet_leaf_16_wb_clk_i _0130_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[96\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_3_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2364__A net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3907__B _1257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_31_wb_clk_i_A clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_7_wb_clk_i clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_2_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2539__A _0840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4434__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3989__C1 _1901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4584__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2274__A _0699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4860_ clknet_leaf_23_wb_clk_i _0474_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[86\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_60_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3811_ _1710_ tms1x00.RAM\[77\]\[3\] _1801_ vssd1 vssd1 vccd1 vccd1 _1805_ sky130_fd_sc_hd__mux2_1
XFILLER_33_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3205__A1 _1334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4791_ clknet_leaf_24_wb_clk_i _0405_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[71\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_3742_ _1708_ tms1x00.RAM\[76\]\[2\] _1762_ vssd1 vssd1 vccd1 vccd1 _1765_ sky130_fd_sc_hd__mux2_1
XFILLER_13_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3673_ _1726_ vssd1 vssd1 vccd1 vccd1 _0390_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4166__C1 _1966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2624_ _1009_ _1011_ _1013_ _1015_ _0804_ vssd1 vssd1 vccd1 vccd1 _1016_ sky130_fd_sc_hd__o221a_1
XANTENNA__2213__S _0668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput102 net102 vssd1 vssd1 vccd1 vccd1 oram_addr[7] sky130_fd_sc_hd__buf_2
Xoutput124 net124 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[17] sky130_fd_sc_hd__buf_2
Xoutput113 net113 vssd1 vssd1 vccd1 vccd1 ram_csb sky130_fd_sc_hd__buf_2
X_2555_ tms1x00.RAM\[84\]\[1\] tms1x00.RAM\[85\]\[1\] tms1x00.RAM\[86\]\[1\] tms1x00.RAM\[87\]\[1\]
+ _0945_ _0791_ vssd1 vssd1 vccd1 vccd1 _0947_ sky130_fd_sc_hd__mux4_1
Xoutput146 net146 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[8] sky130_fd_sc_hd__buf_2
Xoutput135 net135 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[27] sky130_fd_sc_hd__buf_2
X_2486_ _0786_ _0878_ _0828_ vssd1 vssd1 vccd1 vccd1 _0879_ sky130_fd_sc_hd__a21o_1
X_4225_ tms1x00.ins_in\[5\] _2087_ vssd1 vssd1 vccd1 vccd1 _2088_ sky130_fd_sc_hd__and2b_1
XFILLER_68_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4156_ _0768_ _1995_ _2027_ _2028_ _0701_ vssd1 vssd1 vccd1 vccd1 _2029_ sky130_fd_sc_hd__o221a_1
XFILLER_29_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3107_ _1364_ tms1x00.RAM\[110\]\[1\] _1397_ vssd1 vssd1 vccd1 vccd1 _1399_ sky130_fd_sc_hd__mux2_1
XFILLER_55_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4927__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4087_ _0718_ _1973_ vssd1 vssd1 vccd1 vccd1 _1978_ sky130_fd_sc_hd__nand2_1
X_3038_ _1035_ tms1x00.RAM\[97\]\[1\] _1356_ vssd1 vssd1 vccd1 vccd1 _1358_ sky130_fd_sc_hd__mux2_1
XANTENNA__3444__A1 _1574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4989_ clknet_leaf_1_wb_clk_i _0599_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[39\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2350__C net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3380__A0 _1485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2802__S0 _0816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4457__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3132__A0 _1368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput37 ram_val[30] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__clkbuf_1
Xinput26 ram_val[20] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_1
Xinput15 ram_val[10] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput48 wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__clkbuf_1
Xinput59 wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2340_ _0737_ vssd1 vssd1 vccd1 vccd1 _0048_ sky130_fd_sc_hd__clkbuf_1
XFILLER_69_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2271_ net77 _0698_ _0700_ wbs_o_buff\[8\] vssd1 vssd1 vccd1 vccd1 _0033_ sky130_fd_sc_hd__a22o_1
XFILLER_78_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4010_ tms1x00.Y\[1\] tms1x00.Y\[0\] vssd1 vssd1 vccd1 vccd1 _1921_ sky130_fd_sc_hd__nand2_1
XFILLER_77_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3426__A1 _1578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4912_ clknet_leaf_6_wb_clk_i _0526_ vssd1 vssd1 vccd1 vccd1 tms1x00.ins_in\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2774__B_N _0955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4843_ clknet_leaf_23_wb_clk_i _0457_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[84\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_4774_ clknet_leaf_17_wb_clk_i _0388_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[66\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3725_ _1755_ vssd1 vssd1 vccd1 vccd1 _0413_ sky130_fd_sc_hd__clkbuf_1
X_3656_ _1229_ _1236_ vssd1 vssd1 vccd1 vccd1 _1717_ sky130_fd_sc_hd__or2_2
X_2607_ tms1x00.RAM\[0\]\[1\] tms1x00.RAM\[1\]\[1\] tms1x00.RAM\[2\]\[1\] tms1x00.RAM\[3\]\[1\]
+ _0955_ _0956_ vssd1 vssd1 vccd1 vccd1 _0999_ sky130_fd_sc_hd__mux4_1
X_3587_ tms1x00.RAM\[58\]\[3\] _1676_ _1670_ vssd1 vssd1 vccd1 vccd1 _1677_ sky130_fd_sc_hd__mux2_1
XFILLER_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2538_ _0928_ _0929_ vssd1 vssd1 vccd1 vccd1 _0930_ sky130_fd_sc_hd__nand2_1
X_4208_ tms1x00.P\[2\] tms1x00.N\[2\] vssd1 vssd1 vccd1 vccd1 _2073_ sky130_fd_sc_hd__and2_1
XFILLER_57_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2469_ tms1x00.RAM\[30\]\[0\] tms1x00.RAM\[31\]\[0\] _0823_ vssd1 vssd1 vccd1 vccd1
+ _0862_ sky130_fd_sc_hd__mux2_1
XFILLER_56_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4139_ _2009_ _1030_ vssd1 vssd1 vccd1 vccd1 _2015_ sky130_fd_sc_hd__and2b_1
XFILLER_56_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3417__A1 _1578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3353__A0 _1485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input45_A ram_val[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3105__A0 _1361_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3408__A1 _1571_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2552__A _0775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4622__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3510_ _1632_ vssd1 vssd1 vccd1 vccd1 _0321_ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2490__S1 _0831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4490_ clknet_leaf_31_wb_clk_i _0111_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[100\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3344__A0 _1485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3441_ _1317_ _1525_ vssd1 vssd1 vccd1 vccd1 _1594_ sky130_fd_sc_hd__nor2_2
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3372_ _1552_ vssd1 vssd1 vccd1 vccd1 _0263_ sky130_fd_sc_hd__clkbuf_1
XFILLER_69_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2323_ tms1x00.Y\[0\] _0717_ _0726_ vssd1 vssd1 vccd1 vccd1 _0727_ sky130_fd_sc_hd__mux2_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2698__A2 tms1x00.RAM\[90\]\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2254_ net5 K_override\[3\] net148 vssd1 vssd1 vccd1 vccd1 _0695_ sky130_fd_sc_hd__mux2_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5042_ clknet_leaf_4_wb_clk_i _0652_ vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__dfxtp_1
XFILLER_66_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2185_ _0659_ vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__clkbuf_1
XFILLER_81_801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3558__A _1229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4826_ clknet_leaf_22_wb_clk_i _0440_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[7\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xwrapped_tms1x00_167 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_167/HI io_oeb[28] sky130_fd_sc_hd__conb_1
Xwrapped_tms1x00_156 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_156/HI io_oeb[17] sky130_fd_sc_hd__conb_1
Xwrapped_tms1x00_178 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_178/HI io_out[1] sky130_fd_sc_hd__conb_1
X_4757_ clknet_leaf_2_wb_clk_i _0371_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[62\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xwrapped_tms1x00_189 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_189/HI oram_addr[8] sky130_fd_sc_hd__conb_1
X_4688_ clknet_leaf_5_wb_clk_i _0302_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[44\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_3708_ tms1x00.RAM\[71\]\[3\] _1676_ _1742_ vssd1 vssd1 vccd1 vccd1 _1746_ sky130_fd_sc_hd__mux2_1
X_3639_ _1706_ tms1x00.RAM\[61\]\[1\] _1704_ vssd1 vssd1 vccd1 vccd1 _1707_ sky130_fd_sc_hd__mux2_1
XANTENNA__3335__A0 _1485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_21_wb_clk_i clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_13_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4645__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3468__A _1286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4795__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3326__A0 _1485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4054__A1 net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3990_ net13 _1899_ vssd1 vssd1 vccd1 vccd1 _1907_ sky130_fd_sc_hd__or2_1
XFILLER_35_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2941_ _1295_ vssd1 vssd1 vccd1 vccd1 _0089_ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4611_ clknet_leaf_11_wb_clk_i _0232_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[28\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_2872_ _0912_ tms1x00.RAM\[17\]\[0\] _1252_ vssd1 vssd1 vccd1 vccd1 _1253_ sky130_fd_sc_hd__mux2_1
XFILLER_30_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3565__A0 _1592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4542_ clknet_leaf_31_wb_clk_i _0163_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[107\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_4473_ clknet_leaf_17_wb_clk_i _0094_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[19\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3317__S _1519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2221__S _0668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3424_ tms1x00.RAM\[40\]\[2\] _1576_ _1580_ vssd1 vssd1 vccd1 vccd1 _1583_ sky130_fd_sc_hd__mux2_1
XANTENNA__3841__A _1224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3355_ _1488_ tms1x00.RAM\[2\]\[1\] _1541_ vssd1 vssd1 vccd1 vccd1 _1543_ sky130_fd_sc_hd__mux2_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3286_ _1503_ vssd1 vssd1 vccd1 vccd1 _0226_ sky130_fd_sc_hd__clkbuf_1
X_2306_ net46 vssd1 vssd1 vccd1 vccd1 _0713_ sky130_fd_sc_hd__inv_2
XFILLER_73_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5025_ clknet_leaf_2_wb_clk_i _0635_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[1\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_2237_ _0686_ vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__clkbuf_1
XANTENNA__2457__A _0779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2828__C1 _0806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4225__A_N tms1x00.ins_in\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4668__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4809_ clknet_leaf_24_wb_clk_i _0423_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[75\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_79_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2454__S1 _0812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2367__A tms1x00.ins_in\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2598__A1 _0932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3198__A _1303_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output76_A net76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3140_ _1418_ vssd1 vssd1 vccd1 vccd1 _0165_ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4810__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3071_ _1378_ vssd1 vssd1 vccd1 vccd1 _0136_ sky130_fd_sc_hd__clkbuf_1
XFILLER_48_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2825__A2 tms1x00.RAM\[62\]\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2286__B1 _0704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4027__A1 net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4960__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3973_ _1896_ vssd1 vssd1 vccd1 vccd1 _0520_ sky130_fd_sc_hd__clkbuf_1
XFILLER_51_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2589__A1 _0948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2853__C_N tms1x00.ram_addr_buff\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2924_ _1227_ _1259_ vssd1 vssd1 vccd1 vccd1 _1285_ sky130_fd_sc_hd__or2_1
XFILLER_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2855_ _1239_ vssd1 vssd1 vccd1 vccd1 _1240_ sky130_fd_sc_hd__buf_4
X_4525_ clknet_leaf_16_wb_clk_i _0146_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[112\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_2786_ tms1x00.RAM\[16\]\[3\] tms1x00.RAM\[17\]\[3\] tms1x00.RAM\[18\]\[3\] tms1x00.RAM\[19\]\[3\]
+ _0924_ _0928_ vssd1 vssd1 vccd1 vccd1 _1176_ sky130_fd_sc_hd__mux4_1
X_4456_ clknet_leaf_12_wb_clk_i _0077_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[18\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_4387_ tms1x00.PA\[2\] net101 _2006_ vssd1 vssd1 vccd1 vccd1 _2177_ sky130_fd_sc_hd__mux2_1
X_3407_ _1261_ _1525_ vssd1 vssd1 vccd1 vccd1 _1572_ sky130_fd_sc_hd__nor2_2
XFILLER_59_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3338_ _1533_ vssd1 vssd1 vccd1 vccd1 _0248_ sky130_fd_sc_hd__clkbuf_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4490__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3269_ _0917_ _1375_ vssd1 vssd1 vccd1 vccd1 _1494_ sky130_fd_sc_hd__or2_1
XFILLER_27_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2277__B1 _0703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5008_ clknet_leaf_0_wb_clk_i _0618_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[20\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_54_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3529__A0 _1592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3746__A _1237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_21_wb_clk_i_A clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_5_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4833__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2796__S _0788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4983__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4009__A1 net79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output114_A net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2666__S1 _0956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3656__A _1229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2640_ _1031_ vssd1 vssd1 vccd1 vccd1 _1032_ sky130_fd_sc_hd__inv_2
X_2571_ tms1x00.RAM\[96\]\[1\] tms1x00.RAM\[97\]\[1\] tms1x00.RAM\[98\]\[1\] tms1x00.RAM\[99\]\[1\]
+ _0945_ _0791_ vssd1 vssd1 vccd1 vccd1 _0963_ sky130_fd_sc_hd__mux4_1
X_4310_ tms1x00.RAM\[20\]\[3\] _1333_ _2131_ vssd1 vssd1 vccd1 vccd1 _2135_ sky130_fd_sc_hd__mux2_1
X_4241_ tms1x00.A\[0\] _2062_ _2096_ vssd1 vssd1 vccd1 vccd1 _2097_ sky130_fd_sc_hd__mux2_1
XFILLER_4_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4172_ tms1x00.PC\[2\] _1908_ _2042_ _1966_ vssd1 vssd1 vccd1 vccd1 _0573_ sky130_fd_sc_hd__o211a_1
XFILLER_67_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3123_ _1408_ vssd1 vssd1 vccd1 vccd1 _0158_ sky130_fd_sc_hd__clkbuf_1
XFILLER_82_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3054_ _1224_ vssd1 vssd1 vccd1 vccd1 _1368_ sky130_fd_sc_hd__clkbuf_4
XFILLER_82_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3956_ _0730_ tms1x00.ram_addr_buff\[2\] _0726_ vssd1 vssd1 vccd1 vccd1 _1887_ sky130_fd_sc_hd__mux2_1
XANTENNA__4706__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2907_ _1275_ vssd1 vssd1 vccd1 vccd1 _0075_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__2470__A _0822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3887_ tms1x00.RAM\[88\]\[3\] _1779_ _1845_ vssd1 vssd1 vccd1 vccd1 _1849_ sky130_fd_sc_hd__mux2_1
XANTENNA__2982__A1 _1245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2838_ tms1x00.ram_addr_buff\[0\] tms1x00.ram_addr_buff\[1\] vssd1 vssd1 vccd1 vccd1
+ _1227_ sky130_fd_sc_hd__nand2_1
XANTENNA__4856__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2769_ _0940_ _1156_ _1158_ _0942_ vssd1 vssd1 vccd1 vccd1 _1159_ sky130_fd_sc_hd__o211a_1
XFILLER_3_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4508_ clknet_leaf_16_wb_clk_i _0129_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[96\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2734__A1 _0040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4439_ clknet_leaf_28_wb_clk_i _0060_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[69\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2593__S0 _0975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3998__B1 net75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2380__A _0040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2973__A1 _1247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5011__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2489__B1 _0039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3150__A1 _1334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4729__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3810_ _1804_ vssd1 vssd1 vccd1 vccd1 _0449_ sky130_fd_sc_hd__clkbuf_1
X_4790_ clknet_leaf_24_wb_clk_i _0404_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[71\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3741_ _1764_ vssd1 vssd1 vccd1 vccd1 _0420_ sky130_fd_sc_hd__clkbuf_1
XFILLER_32_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4879__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3672_ _1710_ tms1x00.RAM\[66\]\[3\] _1722_ vssd1 vssd1 vccd1 vccd1 _1726_ sky130_fd_sc_hd__mux2_1
X_2623_ _0819_ _1014_ _0775_ vssd1 vssd1 vccd1 vccd1 _1015_ sky130_fd_sc_hd__o21ai_1
X_2554_ tms1x00.RAM\[80\]\[1\] tms1x00.RAM\[81\]\[1\] tms1x00.RAM\[82\]\[1\] tms1x00.RAM\[83\]\[1\]
+ _0945_ _0791_ vssd1 vssd1 vccd1 vccd1 _0946_ sky130_fd_sc_hd__mux4_1
Xoutput103 net103 vssd1 vssd1 vccd1 vccd1 oram_csb sky130_fd_sc_hd__buf_2
Xoutput125 net125 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[18] sky130_fd_sc_hd__buf_2
Xoutput114 net114 vssd1 vssd1 vccd1 vccd1 ram_web sky130_fd_sc_hd__buf_2
Xoutput147 net147 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[9] sky130_fd_sc_hd__buf_2
Xoutput136 net136 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[28] sky130_fd_sc_hd__buf_2
X_2485_ tms1x00.RAM\[4\]\[0\] tms1x00.RAM\[5\]\[0\] _0826_ vssd1 vssd1 vccd1 vccd1
+ _0878_ sky130_fd_sc_hd__mux2_1
XFILLER_68_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4010__A tms1x00.Y\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4224_ _0746_ _2086_ vssd1 vssd1 vccd1 vccd1 _2087_ sky130_fd_sc_hd__nor2_1
XFILLER_68_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4155_ tms1x00.SR\[0\] vssd1 vssd1 vccd1 vccd1 _2028_ sky130_fd_sc_hd__inv_2
XANTENNA__3141__A1 _1334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3106_ _1398_ vssd1 vssd1 vccd1 vccd1 _0151_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4086_ _1977_ vssd1 vssd1 vccd1 vccd1 _0552_ sky130_fd_sc_hd__clkbuf_1
XFILLER_71_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3037_ _1357_ vssd1 vssd1 vccd1 vccd1 _0123_ sky130_fd_sc_hd__clkbuf_1
XFILLER_36_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4988_ clknet_leaf_0_wb_clk_i _0598_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[39\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3296__A _1249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3939_ tms1x00.RAM\[90\]\[2\] _1330_ _1875_ vssd1 vssd1 vccd1 vccd1 _1878_ sky130_fd_sc_hd__mux2_1
XFILLER_20_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2802__S1 _0927_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3199__A1 _1324_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput27 ram_val[21] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput16 ram_val[11] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput38 ram_val[31] vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__clkbuf_1
Xinput49 wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__clkbuf_4
XFILLER_6_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3934__A _1258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3371__A1 _1456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2270_ net76 _0698_ _0700_ wbs_o_buff\[7\] vssd1 vssd1 vccd1 vccd1 _0032_ sky130_fd_sc_hd__a22o_1
XFILLER_77_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4551__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4084__C1 _1966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2285__A _0699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4911_ clknet_leaf_7_wb_clk_i _0525_ vssd1 vssd1 vccd1 vccd1 tms1x00.ins_in\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XANTENNA_clkbuf_2_0__f_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4842_ clknet_leaf_19_wb_clk_i _0456_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[84\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4773_ clknet_leaf_19_wb_clk_i _0387_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[66\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3724_ tms1x00.RAM\[6\]\[2\] _1674_ _1752_ vssd1 vssd1 vccd1 vccd1 _1755_ sky130_fd_sc_hd__mux2_1
X_3655_ _1716_ vssd1 vssd1 vccd1 vccd1 _0382_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3844__A _1257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2606_ _0787_ _0994_ _0997_ vssd1 vssd1 vccd1 vccd1 _0998_ sky130_fd_sc_hd__a21oi_1
XANTENNA__3362__A1 _1456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3586_ _1224_ vssd1 vssd1 vccd1 vccd1 _1676_ sky130_fd_sc_hd__clkbuf_4
X_2537_ tms1x00.RAM\[70\]\[1\] tms1x00.RAM\[71\]\[1\] _0924_ vssd1 vssd1 vccd1 vccd1
+ _0929_ sky130_fd_sc_hd__mux2_1
X_2468_ _0859_ _0860_ _0783_ vssd1 vssd1 vccd1 vccd1 _0861_ sky130_fd_sc_hd__mux2_1
XFILLER_69_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4207_ _2072_ vssd1 vssd1 vccd1 vccd1 _0578_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2399_ tms1x00.RAM\[94\]\[0\] tms1x00.RAM\[95\]\[0\] _0788_ vssd1 vssd1 vccd1 vccd1
+ _0792_ sky130_fd_sc_hd__mux2_1
XFILLER_29_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4138_ tms1x00.P\[0\] _2007_ _2010_ _2014_ vssd1 vssd1 vccd1 vccd1 _0567_ sky130_fd_sc_hd__o22a_1
XFILLER_28_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4069_ net71 _1960_ vssd1 vssd1 vccd1 vccd1 _1965_ sky130_fd_sc_hd__or2_1
XFILLER_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2720__S0 _0816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2923__A _1283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4424__CLK clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2787__S0 _0923_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4574__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input38_A ram_val[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3592__A1 _1672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4917__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3440_ _1593_ vssd1 vssd1 vccd1 vccd1 _0290_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2778__S0 _0873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3371_ tms1x00.RAM\[36\]\[0\] _1456_ _1551_ vssd1 vssd1 vccd1 vccd1 _1552_ sky130_fd_sc_hd__mux2_1
XFILLER_69_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2322_ _0725_ vssd1 vssd1 vccd1 vccd1 _0726_ sky130_fd_sc_hd__buf_4
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5041_ clknet_leaf_4_wb_clk_i _0651_ vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__dfxtp_1
XFILLER_2_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2253_ _0694_ vssd1 vssd1 vccd1 vccd1 tms1x00.K_in\[2\] sky130_fd_sc_hd__clkbuf_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2184_ net25 wbs_o_buff\[1\] _0657_ vssd1 vssd1 vccd1 vccd1 _0659_ sky130_fd_sc_hd__mux2_1
XFILLER_81_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_0_wb_clk_i sky130_fd_sc_hd__clkbuf_16
XANTENNA__2219__S _0668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4057__C1 _1931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3558__B _1283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4447__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4825_ clknet_leaf_22_wb_clk_i _0439_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[7\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapped_tms1x00_168 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_168/HI io_oeb[29] sky130_fd_sc_hd__conb_1
Xwrapped_tms1x00_157 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_157/HI io_oeb[18] sky130_fd_sc_hd__conb_1
Xwrapped_tms1x00_179 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_179/HI io_out[2] sky130_fd_sc_hd__conb_1
X_4756_ clknet_leaf_11_wb_clk_i _0370_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[63\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_4687_ clknet_leaf_5_wb_clk_i _0301_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[44\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_3707_ _1745_ vssd1 vssd1 vccd1 vccd1 _0405_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4597__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3638_ _1034_ vssd1 vssd1 vccd1 vccd1 _1706_ sky130_fd_sc_hd__buf_2
X_3569_ _1665_ vssd1 vssd1 vccd1 vccd1 _0347_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3099__A0 _1366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2846__A0 _1130_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4048__C1 _1931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3468__B _1525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3574__A1 _1578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2940_ _1130_ tms1x00.RAM\[49\]\[2\] _1292_ vssd1 vssd1 vccd1 vccd1 _1295_ sky130_fd_sc_hd__mux2_1
XANTENNA__2563__A _0799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2871_ _1250_ _1251_ vssd1 vssd1 vccd1 vccd1 _1252_ sky130_fd_sc_hd__or2_2
X_4610_ clknet_leaf_11_wb_clk_i _0231_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[28\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4541_ clknet_leaf_14_wb_clk_i _0162_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[108\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_4472_ clknet_leaf_12_wb_clk_i _0093_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[19\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2773__C1 _0944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3317__A1 _1459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3423_ _1582_ vssd1 vssd1 vccd1 vccd1 _0284_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4002__B tms1x00.Y\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3354_ _1542_ vssd1 vssd1 vccd1 vccd1 _0255_ sky130_fd_sc_hd__clkbuf_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3285_ tms1x00.RAM\[25\]\[3\] _1463_ _1499_ vssd1 vssd1 vccd1 vccd1 _1503_ sky130_fd_sc_hd__mux2_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2305_ _0712_ vssd1 vssd1 vccd1 vccd1 _0027_ sky130_fd_sc_hd__clkbuf_1
X_5024_ clknet_leaf_2_wb_clk_i _0634_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[1\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2236_ net32 wbs_o_buff\[26\] _0679_ vssd1 vssd1 vccd1 vccd1 _0686_ sky130_fd_sc_hd__mux2_1
XFILLER_72_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_11_wb_clk_i_A clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_4808_ clknet_leaf_20_wb_clk_i _0422_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[76\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4739_ clknet_leaf_28_wb_clk_i _0353_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[58\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3556__A1 _1578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3308__A1 _1459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2648__A _0807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2383__A _0775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4762__CLK clknet_leaf_20_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2598__A2 _0989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3198__B _1430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3547__A1 _1578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output69_A net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3070_ _1364_ tms1x00.RAM\[114\]\[1\] _1376_ vssd1 vssd1 vccd1 vccd1 _1378_ sky130_fd_sc_hd__mux2_1
XFILLER_82_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2286__A1 net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3972_ net103 _1895_ vssd1 vssd1 vccd1 vccd1 _1896_ sky130_fd_sc_hd__or2_1
XANTENNA__2589__A2 _0974_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2923_ _1283_ vssd1 vssd1 vccd1 vccd1 _1284_ sky130_fd_sc_hd__clkbuf_8
X_2854_ tms1x00.ram_addr_buff\[1\] _1238_ _0717_ vssd1 vssd1 vccd1 vccd1 _1239_ sky130_fd_sc_hd__or3b_1
XFILLER_31_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2785_ _0821_ _1159_ _1163_ _0040_ _1174_ vssd1 vssd1 vccd1 vccd1 _1175_ sky130_fd_sc_hd__o311a_1
XANTENNA__3538__A1 _1578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4524_ clknet_leaf_16_wb_clk_i _0145_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[112\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4455_ clknet_leaf_12_wb_clk_i _0076_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[18\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_4386_ _2176_ vssd1 vssd1 vccd1 vccd1 _0653_ sky130_fd_sc_hd__clkbuf_1
X_3406_ _0911_ vssd1 vssd1 vccd1 vccd1 _1571_ sky130_fd_sc_hd__clkbuf_4
XFILLER_58_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4635__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3337_ _1488_ tms1x00.RAM\[31\]\[1\] _1531_ vssd1 vssd1 vccd1 vccd1 _1533_ sky130_fd_sc_hd__mux2_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3268_ _1493_ vssd1 vssd1 vccd1 vccd1 _0218_ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2277__A1 net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2219_ net23 wbs_o_buff\[18\] _0668_ vssd1 vssd1 vccd1 vccd1 _0677_ sky130_fd_sc_hd__mux2_1
XANTENNA__4785__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3199_ tms1x00.RAM\[120\]\[0\] _1324_ _1451_ vssd1 vssd1 vccd1 vccd1 _1452_ sky130_fd_sc_hd__mux2_1
X_5007_ clknet_leaf_1_wb_clk_i _0617_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[20\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_66_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3746__B _1286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3762__A _1129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2378__A _0738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input20_A ram_val[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2268__A1 _0701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output107_A net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4508__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2841__A _0914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2440__B2 _0807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3656__B _1236_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4193__A1 tms1x00.ins_in\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2570_ _0940_ _0961_ vssd1 vssd1 vccd1 vccd1 _0962_ sky130_fd_sc_hd__or2_1
XANTENNA__4658__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4240_ _0762_ _0738_ _0746_ _2058_ vssd1 vssd1 vccd1 vccd1 _2096_ sky130_fd_sc_hd__nor4_4
X_4171_ net148 _0721_ _2038_ _2040_ _2041_ vssd1 vssd1 vccd1 vccd1 _2042_ sky130_fd_sc_hd__a221o_1
XFILLER_68_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3122_ tms1x00.RAM\[10\]\[3\] _1334_ _1404_ vssd1 vssd1 vccd1 vccd1 _1408_ sky130_fd_sc_hd__mux2_1
XFILLER_67_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3053_ _1367_ vssd1 vssd1 vccd1 vccd1 _0129_ sky130_fd_sc_hd__clkbuf_1
XFILLER_36_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4008__A _0732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3955_ _1886_ vssd1 vssd1 vccd1 vccd1 _0512_ sky130_fd_sc_hd__clkbuf_1
X_2906_ _0912_ tms1x00.RAM\[18\]\[0\] _1274_ vssd1 vssd1 vccd1 vccd1 _1275_ sky130_fd_sc_hd__mux2_1
X_3886_ _1848_ vssd1 vssd1 vccd1 vccd1 _0481_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4184__A1 _0760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2837_ _1226_ vssd1 vssd1 vccd1 vccd1 _0054_ sky130_fd_sc_hd__clkbuf_1
X_2768_ _0798_ _1157_ vssd1 vssd1 vccd1 vccd1 _1158_ sky130_fd_sc_hd__or2_1
X_4507_ clknet_leaf_16_wb_clk_i _0128_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[96\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_2699_ _1086_ _1088_ _1089_ _0922_ _0942_ vssd1 vssd1 vccd1 vccd1 _1090_ sky130_fd_sc_hd__o221a_1
X_4438_ clknet_leaf_28_wb_clk_i _0059_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[69\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_4369_ tms1x00.RAM\[9\]\[1\] _1327_ _2166_ vssd1 vssd1 vccd1 vccd1 _2168_ sky130_fd_sc_hd__mux2_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2593__S1 _0791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2926__A _1284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3998__A1 _0701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4175__A1 tms1x00.PC\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4800__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2186__A0 net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input68_A wbs_we_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4950__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3686__A0 _1706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2489__A1 _0806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3989__A1 _0748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3740_ _1706_ tms1x00.RAM\[76\]\[1\] _1762_ vssd1 vssd1 vccd1 vccd1 _1764_ sky130_fd_sc_hd__mux2_1
X_3671_ _1725_ vssd1 vssd1 vccd1 vccd1 _0389_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__2290__B _0704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4166__A1 _0760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2622_ tms1x00.RAM\[36\]\[1\] tms1x00.RAM\[37\]\[1\] tms1x00.RAM\[38\]\[1\] tms1x00.RAM\[39\]\[1\]
+ _0808_ _0831_ vssd1 vssd1 vccd1 vccd1 _1014_ sky130_fd_sc_hd__mux4_2
Xoutput104 net104 vssd1 vssd1 vccd1 vccd1 ram_adrb[0] sky130_fd_sc_hd__buf_2
Xoutput115 net115 vssd1 vssd1 vccd1 vccd1 wbs_ack_o sky130_fd_sc_hd__buf_2
X_2553_ _0808_ vssd1 vssd1 vccd1 vccd1 _0945_ sky130_fd_sc_hd__buf_8
Xoutput126 net126 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[19] sky130_fd_sc_hd__buf_2
Xoutput137 net137 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[29] sky130_fd_sc_hd__buf_2
X_2484_ _0822_ _0876_ vssd1 vssd1 vccd1 vccd1 _0877_ sky130_fd_sc_hd__and2_1
XANTENNA__4010__B tms1x00.Y\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3677__A0 _1706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4223_ _0744_ _0904_ _2085_ _0750_ vssd1 vssd1 vccd1 vccd1 _2086_ sky130_fd_sc_hd__o22a_1
X_4154_ _2026_ _0744_ _0750_ _1975_ vssd1 vssd1 vccd1 vccd1 _2027_ sky130_fd_sc_hd__or4_4
X_4085_ tms1x00.status _0738_ _1972_ vssd1 vssd1 vccd1 vccd1 _1977_ sky130_fd_sc_hd__or3_1
X_3105_ _1361_ tms1x00.RAM\[110\]\[0\] _1397_ vssd1 vssd1 vccd1 vccd1 _1398_ sky130_fd_sc_hd__mux2_1
XFILLER_28_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3036_ _0912_ tms1x00.RAM\[97\]\[0\] _1356_ vssd1 vssd1 vccd1 vccd1 _1357_ sky130_fd_sc_hd__mux2_1
XFILLER_70_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4823__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3577__A _1284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4987_ clknet_leaf_35_wb_clk_i _0597_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[39\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3296__B _1409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3938_ _1877_ vssd1 vssd1 vccd1 vccd1 _0504_ sky130_fd_sc_hd__clkbuf_1
XFILLER_20_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3869_ tms1x00.RAM\[86\]\[3\] _1779_ _1835_ vssd1 vssd1 vccd1 vccd1 _1839_ sky130_fd_sc_hd__mux2_1
XANTENNA__4973__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3516__S _1634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3668__A0 _1706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_15_wb_clk_i clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_59_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput28 ram_val[22] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__clkbuf_1
Xinput17 ram_val[12] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4148__B2 _0732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput39 ram_val[3] vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3934__B _1403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3659__A0 _1706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4846__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4910_ clknet_leaf_8_wb_clk_i _0524_ vssd1 vssd1 vccd1 vccd1 tms1x00.ins_in\[4\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2634__A1 _0783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4841_ clknet_leaf_23_wb_clk_i _0455_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[84\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_61_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3397__A _1251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4387__A1 net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4772_ clknet_leaf_18_wb_clk_i _0386_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[67\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3723_ _1754_ vssd1 vssd1 vccd1 vccd1 _0412_ sky130_fd_sc_hd__clkbuf_1
X_3654_ _1710_ tms1x00.RAM\[60\]\[3\] _1712_ vssd1 vssd1 vccd1 vccd1 _1716_ sky130_fd_sc_hd__mux2_1
XFILLER_9_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3844__B _1273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2605_ _0928_ _0995_ _0996_ vssd1 vssd1 vccd1 vccd1 _0997_ sky130_fd_sc_hd__a21o_1
X_3585_ _1675_ vssd1 vssd1 vccd1 vccd1 _0353_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4021__A _0732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2536_ _0927_ vssd1 vssd1 vccd1 vccd1 _0928_ sky130_fd_sc_hd__buf_4
X_2467_ tms1x00.RAM\[20\]\[0\] tms1x00.RAM\[21\]\[0\] tms1x00.RAM\[22\]\[0\] tms1x00.RAM\[23\]\[0\]
+ _0830_ _0831_ vssd1 vssd1 vccd1 vccd1 _0860_ sky130_fd_sc_hd__mux4_2
XFILLER_69_863 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4206_ _0766_ _2071_ vssd1 vssd1 vccd1 vccd1 _2072_ sky130_fd_sc_hd__and2_1
XFILLER_68_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2398_ _0780_ vssd1 vssd1 vccd1 vccd1 _0791_ sky130_fd_sc_hd__buf_6
XFILLER_68_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4137_ tms1x00.ins_in\[4\] _1031_ _2011_ _2013_ vssd1 vssd1 vccd1 vccd1 _2014_ sky130_fd_sc_hd__a211o_1
XFILLER_28_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4068_ _0742_ tms1x00.A\[2\] vssd1 vssd1 vccd1 vccd1 _1964_ sky130_fd_sc_hd__and2b_1
X_3019_ _1347_ vssd1 vssd1 vccd1 vccd1 _0115_ sky130_fd_sc_hd__clkbuf_1
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2720__S1 _0977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5001__CLK clknet_leaf_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2787__S1 _0927_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4106__A net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4369__A1 _1327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2778__S1 _0977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3370_ _1337_ _1525_ vssd1 vssd1 vccd1 vccd1 _1551_ sky130_fd_sc_hd__nor2_2
X_2321_ _0718_ _0724_ vssd1 vssd1 vccd1 vccd1 _0725_ sky130_fd_sc_hd__nand2_2
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2252_ net4 K_override\[2\] net148 vssd1 vssd1 vccd1 vccd1 _0694_ sky130_fd_sc_hd__mux2_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5040_ clknet_leaf_4_wb_clk_i _0650_ vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__dfxtp_1
XFILLER_2_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2183_ _0658_ vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__clkbuf_1
XFILLER_66_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5024__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4016__A _0732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4824_ clknet_leaf_18_wb_clk_i _0438_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[80\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4755_ clknet_leaf_11_wb_clk_i _0369_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[63\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xwrapped_tms1x00_169 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_169/HI io_oeb[30] sky130_fd_sc_hd__conb_1
Xwrapped_tms1x00_158 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_158/HI io_oeb[19] sky130_fd_sc_hd__conb_1
XANTENNA__2466__S0 _0830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3706_ tms1x00.RAM\[71\]\[2\] _1674_ _1742_ vssd1 vssd1 vccd1 vccd1 _1745_ sky130_fd_sc_hd__mux2_1
X_4686_ clknet_leaf_4_wb_clk_i _0300_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[44\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_3637_ _1705_ vssd1 vssd1 vccd1 vccd1 _0375_ sky130_fd_sc_hd__clkbuf_1
XFILLER_1_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3568_ tms1x00.RAM\[5\]\[0\] _1571_ _1664_ vssd1 vssd1 vccd1 vccd1 _1665_ sky130_fd_sc_hd__mux2_1
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2519_ _0911_ vssd1 vssd1 vccd1 vccd1 _0912_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3499_ _1626_ vssd1 vssd1 vccd1 vccd1 _0316_ sky130_fd_sc_hd__clkbuf_1
XFILLER_57_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3765__A _1224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_30_wb_clk_i clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_4_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4691__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input50_A wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3005__A _0914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4039__B1 net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2870_ _0728_ _1228_ _0717_ vssd1 vssd1 vccd1 vccd1 _1251_ sky130_fd_sc_hd__or3b_4
XFILLER_31_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2448__S0 _0840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4270__S _2111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4540_ clknet_leaf_14_wb_clk_i _0161_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[108\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_4471_ clknet_leaf_12_wb_clk_i _0092_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[19\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_3422_ tms1x00.RAM\[40\]\[1\] _1574_ _1580_ vssd1 vssd1 vccd1 vccd1 _1582_ sky130_fd_sc_hd__mux2_1
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2620__S0 _0840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3353_ _1485_ tms1x00.RAM\[2\]\[0\] _1541_ vssd1 vssd1 vccd1 vccd1 _1542_ sky130_fd_sc_hd__mux2_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3284_ _1502_ vssd1 vssd1 vccd1 vccd1 _0225_ sky130_fd_sc_hd__clkbuf_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2304_ wbs_o_buff\[31\] _0699_ vssd1 vssd1 vccd1 vccd1 _0712_ sky130_fd_sc_hd__and2_1
XFILLER_57_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2828__A1 _0940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5023_ clknet_leaf_11_wb_clk_i _0633_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[1\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2235_ _0685_ vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__clkbuf_1
XFILLER_66_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4414__CLK clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4807_ clknet_leaf_18_wb_clk_i _0421_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[76\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2999_ _1223_ vssd1 vssd1 vccd1 vccd1 _1333_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__2439__S0 _0830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4738_ clknet_leaf_26_wb_clk_i _0352_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[58\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_4669_ clknet_leaf_10_wb_clk_i _0290_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[3\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_79_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_7_wb_clk_i_A clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_1_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4907__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3495__A _1337_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2603__S _0975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4103__B _0738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2755__B1 _0828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2839__A tms1x00.ram_addr_buff\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4437__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2286__A2 _0697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4587__CLK clknet_leaf_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4265__S _2106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3971_ _0742_ net6 _0724_ vssd1 vssd1 vccd1 vccd1 _1895_ sky130_fd_sc_hd__mux2_1
XFILLER_51_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2922_ tms1x00.ram_addr_buff\[6\] tms1x00.ram_addr_buff\[5\] tms1x00.ram_addr_buff\[4\]
+ vssd1 vssd1 vccd1 vccd1 _1283_ sky130_fd_sc_hd__nand3b_4
XFILLER_44_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2853_ tms1x00.ram_addr_buff\[3\] _0915_ tms1x00.ram_addr_buff\[2\] vssd1 vssd1 vccd1
+ vccd1 _1238_ sky130_fd_sc_hd__or3b_1
X_2784_ _0944_ _1167_ _1169_ _0804_ _1173_ vssd1 vssd1 vccd1 vccd1 _1174_ sky130_fd_sc_hd__a311o_1
X_4523_ clknet_leaf_14_wb_clk_i _0144_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[112\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_4454_ clknet_leaf_12_wb_clk_i _0075_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[18\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_3405_ _1570_ vssd1 vssd1 vccd1 vccd1 _0278_ sky130_fd_sc_hd__clkbuf_1
X_4385_ tms1x00.PA\[1\] net100 _2006_ vssd1 vssd1 vccd1 vccd1 _2176_ sky130_fd_sc_hd__mux2_1
XFILLER_59_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3336_ _1532_ vssd1 vssd1 vccd1 vccd1 _0247_ sky130_fd_sc_hd__clkbuf_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3267_ _1492_ tms1x00.RAM\[126\]\[3\] _1486_ vssd1 vssd1 vccd1 vccd1 _1493_ sky130_fd_sc_hd__mux2_1
XFILLER_39_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5006_ clknet_leaf_1_wb_clk_i _0616_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[20\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2218_ _0676_ vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__clkbuf_1
X_3198_ _1303_ _1430_ vssd1 vssd1 vccd1 vccd1 _1451_ sky130_fd_sc_hd__nor2_2
XFILLER_27_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2484__A _0822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2659__A _0798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2378__B _0760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input13_A oram_value[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2394__A _0786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2841__B _1229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4178__C1 _1966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2333__S _0726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2823__S0 _0816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output81_A net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4170_ _2038_ _2040_ vssd1 vssd1 vccd1 vccd1 _2041_ sky130_fd_sc_hd__nor2_1
XANTENNA__2900__A0 _1130_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3121_ _1407_ vssd1 vssd1 vccd1 vccd1 _0157_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3052_ _1366_ tms1x00.RAM\[96\]\[2\] _1362_ vssd1 vssd1 vccd1 vccd1 _1367_ sky130_fd_sc_hd__mux2_1
XFILLER_55_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4008__B _0730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3954_ tms1x00.Y\[1\] _0728_ _0726_ vssd1 vssd1 vccd1 vccd1 _1886_ sky130_fd_sc_hd__mux2_1
XFILLER_32_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2905_ _1250_ _1273_ vssd1 vssd1 vccd1 vccd1 _1274_ sky130_fd_sc_hd__or2_2
X_3885_ tms1x00.RAM\[88\]\[2\] _1777_ _1845_ vssd1 vssd1 vccd1 vccd1 _1848_ sky130_fd_sc_hd__mux2_1
XANTENNA__4024__A tms1x00.Y\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2836_ _1225_ tms1x00.RAM\[109\]\[3\] _0918_ vssd1 vssd1 vccd1 vccd1 _1226_ sky130_fd_sc_hd__mux2_1
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2814__S0 _0923_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2767_ tms1x00.RAM\[104\]\[3\] tms1x00.RAM\[105\]\[3\] tms1x00.RAM\[106\]\[3\] tms1x00.RAM\[107\]\[3\]
+ _0840_ _0813_ vssd1 vssd1 vccd1 vccd1 _1157_ sky130_fd_sc_hd__mux4_1
XANTENNA__4602__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4506_ clknet_leaf_16_wb_clk_i _0127_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[96\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_2698_ tms1x00.RAM\[88\]\[2\] tms1x00.RAM\[89\]\[2\] tms1x00.RAM\[90\]\[2\] tms1x00.RAM\[91\]\[2\]
+ _0931_ _0932_ vssd1 vssd1 vccd1 vccd1 _1089_ sky130_fd_sc_hd__mux4_1
X_4437_ clknet_leaf_16_wb_clk_i _0058_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[99\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4752__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input5_A io_in[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3695__A1 _1672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4368_ _2167_ vssd1 vssd1 vccd1 vccd1 _0644_ sky130_fd_sc_hd__clkbuf_1
XFILLER_58_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4299_ _1821_ tms1x00.RAM\[16\]\[2\] _2126_ vssd1 vssd1 vccd1 vccd1 _2129_ sky130_fd_sc_hd__mux2_1
X_3319_ tms1x00.RAM\[26\]\[2\] _1461_ _1519_ vssd1 vssd1 vccd1 vccd1 _1522_ sky130_fd_sc_hd__mux2_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2926__B _1286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3989__A2 _0724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4109__A net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2852__A _1236_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2949__A0 _1130_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4625__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3610__A1 _1672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3670_ _1708_ tms1x00.RAM\[66\]\[2\] _1722_ vssd1 vssd1 vccd1 vccd1 _1725_ sky130_fd_sc_hd__mux2_1
XANTENNA__3683__A _1236_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2621_ _0798_ _1012_ vssd1 vssd1 vccd1 vccd1 _1013_ sky130_fd_sc_hd__nor2_1
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2552_ _0775_ vssd1 vssd1 vccd1 vccd1 _0944_ sky130_fd_sc_hd__clkbuf_4
Xoutput105 net105 vssd1 vssd1 vccd1 vccd1 ram_adrb[1] sky130_fd_sc_hd__buf_2
Xoutput116 net116 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[0] sky130_fd_sc_hd__buf_2
Xoutput138 net138 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[2] sky130_fd_sc_hd__buf_2
Xoutput127 net127 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[1] sky130_fd_sc_hd__buf_2
XANTENNA__3126__A0 _1361_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4222_ _0743_ tms1x00.ins_in\[2\] tms1x00.ins_in\[1\] _0742_ vssd1 vssd1 vccd1 vccd1
+ _2085_ sky130_fd_sc_hd__or4_1
X_2483_ tms1x00.RAM\[6\]\[0\] tms1x00.RAM\[7\]\[0\] _0823_ vssd1 vssd1 vccd1 vccd1
+ _0876_ sky130_fd_sc_hd__mux2_1
XFILLER_68_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4153_ tms1x00.CL vssd1 vssd1 vccd1 vccd1 _2026_ sky130_fd_sc_hd__inv_2
X_3104_ _0913_ _1396_ vssd1 vssd1 vccd1 vccd1 _1397_ sky130_fd_sc_hd__or2_2
XFILLER_56_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4084_ tms1x00.CL _1973_ _1976_ _1966_ vssd1 vssd1 vccd1 vccd1 _0551_ sky130_fd_sc_hd__o211a_1
X_3035_ _0913_ _1251_ vssd1 vssd1 vccd1 vccd1 _1356_ sky130_fd_sc_hd__or2_2
XFILLER_37_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4019__A tms1x00.Y\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4986_ clknet_leaf_1_wb_clk_i _0596_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[39\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_3937_ tms1x00.RAM\[90\]\[1\] _1327_ _1875_ vssd1 vssd1 vccd1 vccd1 _1877_ sky130_fd_sc_hd__mux2_1
XANTENNA__3577__B _1403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3601__A1 _1672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3868_ _1838_ vssd1 vssd1 vccd1 vccd1 _0473_ sky130_fd_sc_hd__clkbuf_1
XFILLER_20_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3799_ _1798_ vssd1 vssd1 vccd1 vccd1 _0444_ sky130_fd_sc_hd__clkbuf_1
X_2819_ tms1x00.RAM\[55\]\[3\] _0931_ vssd1 vssd1 vccd1 vccd1 _1209_ sky130_fd_sc_hd__or2b_1
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4093__A1 tms1x00.PC\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4648__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3768__A _1237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput18 ram_val[13] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4798__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput29 ram_val[23] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2634__A2 _1025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4840_ clknet_leaf_23_wb_clk_i _0454_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[85\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_61_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4771_ clknet_leaf_18_wb_clk_i _0385_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[67\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3722_ tms1x00.RAM\[6\]\[1\] _1672_ _1752_ vssd1 vssd1 vccd1 vccd1 _1754_ sky130_fd_sc_hd__mux2_1
X_3653_ _1715_ vssd1 vssd1 vccd1 vccd1 _0381_ sky130_fd_sc_hd__clkbuf_1
X_2604_ _0794_ vssd1 vssd1 vccd1 vccd1 _0996_ sky130_fd_sc_hd__clkbuf_4
X_3584_ tms1x00.RAM\[58\]\[2\] _1674_ _1670_ vssd1 vssd1 vccd1 vccd1 _1675_ sky130_fd_sc_hd__mux2_1
X_2535_ _0850_ vssd1 vssd1 vccd1 vccd1 _0927_ sky130_fd_sc_hd__buf_4
X_2466_ tms1x00.RAM\[16\]\[0\] tms1x00.RAM\[17\]\[0\] tms1x00.RAM\[18\]\[0\] tms1x00.RAM\[19\]\[0\]
+ _0830_ _0831_ vssd1 vssd1 vccd1 vccd1 _0859_ sky130_fd_sc_hd__mux4_1
XFILLER_68_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4205_ tms1x00.Y\[1\] _2070_ _2063_ vssd1 vssd1 vccd1 vccd1 _2071_ sky130_fd_sc_hd__mux2_1
XFILLER_69_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4136_ _0743_ tms1x00.K_latch\[0\] _1956_ _2012_ tms1x00.Y\[0\] vssd1 vssd1 vccd1
+ vccd1 _2013_ sky130_fd_sc_hd__a32o_1
X_2397_ tms1x00.RAM\[92\]\[0\] tms1x00.RAM\[93\]\[0\] _0789_ vssd1 vssd1 vccd1 vccd1
+ _0790_ sky130_fd_sc_hd__mux2_1
X_4067_ _1958_ _1962_ _1963_ _1931_ vssd1 vssd1 vccd1 vccd1 _0547_ sky130_fd_sc_hd__o211a_1
XANTENNA_clkbuf_leaf_30_wb_clk_i_A clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_71_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3018_ _0912_ tms1x00.RAM\[0\]\[0\] _1346_ vssd1 vssd1 vccd1 vccd1 _1347_ sky130_fd_sc_hd__mux2_1
XFILLER_37_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4969_ clknet_leaf_9_wb_clk_i _0579_ vssd1 vssd1 vccd1 vccd1 tms1x00.Y\[2\] sky130_fd_sc_hd__dfxtp_2
XFILLER_20_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3527__S _1639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2431__S _0823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4470__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2320_ _0723_ vssd1 vssd1 vccd1 vccd1 _0724_ sky130_fd_sc_hd__clkbuf_4
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2251_ _0693_ vssd1 vssd1 vccd1 vccd1 tms1x00.K_in\[1\] sky130_fd_sc_hd__clkbuf_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4813__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4268__S _2111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2296__B _0704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2182_ net14 wbs_o_buff\[0\] _0657_ vssd1 vssd1 vccd1 vccd1 _0658_ sky130_fd_sc_hd__mux2_1
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4963__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_0_wb_clk_i clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_4823_ clknet_leaf_17_wb_clk_i _0437_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[80\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_34_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4754_ clknet_leaf_2_wb_clk_i _0368_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[63\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwrapped_tms1x00_159 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_159/HI io_oeb[20] sky130_fd_sc_hd__conb_1
XANTENNA__2466__S1 _0831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2240__A0 net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3705_ _1744_ vssd1 vssd1 vccd1 vccd1 _0404_ sky130_fd_sc_hd__clkbuf_1
X_4685_ clknet_leaf_3_wb_clk_i _0299_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[44\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_3636_ _1703_ tms1x00.RAM\[61\]\[0\] _1704_ vssd1 vssd1 vccd1 vccd1 _1705_ sky130_fd_sc_hd__mux2_1
X_3567_ _1240_ _1344_ vssd1 vssd1 vccd1 vccd1 _1664_ sky130_fd_sc_hd__nor2_2
XANTENNA__3740__A0 _1706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2518_ _0910_ vssd1 vssd1 vccd1 vccd1 _0911_ sky130_fd_sc_hd__buf_4
XANTENNA__3871__A _1303_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2543__A1 _0922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3498_ tms1x00.RAM\[4\]\[1\] _1574_ _1624_ vssd1 vssd1 vccd1 vccd1 _1626_ sky130_fd_sc_hd__mux2_1
X_2449_ tms1x00.RAM\[100\]\[0\] tms1x00.RAM\[101\]\[0\] tms1x00.RAM\[102\]\[0\] tms1x00.RAM\[103\]\[0\]
+ _0815_ _0779_ vssd1 vssd1 vccd1 vccd1 _0842_ sky130_fd_sc_hd__mux4_1
XFILLER_68_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4119_ tms1x00.PB\[1\] tms1x00.PA\[1\] _1996_ vssd1 vssd1 vccd1 vccd1 _1999_ sky130_fd_sc_hd__mux2_1
X_5099_ net52 vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__clkbuf_2
XFILLER_72_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3559__A0 _1585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input43_A ram_val[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4986__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3005__B _1337_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3798__A0 _1706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4117__A net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2448__S1 _0813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2773__A1 _0922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4470_ clknet_leaf_12_wb_clk_i _0091_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[19\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3421_ _1581_ vssd1 vssd1 vccd1 vccd1 _0283_ sky130_fd_sc_hd__clkbuf_1
X_3352_ _1273_ _1343_ vssd1 vssd1 vccd1 vccd1 _1541_ sky130_fd_sc_hd__or2_2
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2620__S1 _0813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2303_ _0711_ vssd1 vssd1 vccd1 vccd1 _0026_ sky130_fd_sc_hd__clkbuf_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3283_ tms1x00.RAM\[25\]\[2\] _1461_ _1499_ vssd1 vssd1 vccd1 vccd1 _1502_ sky130_fd_sc_hd__mux2_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5022_ clknet_leaf_2_wb_clk_i _0632_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[1\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2289__B1 _0704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2234_ net31 wbs_o_buff\[25\] _0679_ vssd1 vssd1 vccd1 vccd1 _0685_ sky130_fd_sc_hd__mux2_1
XFILLER_65_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4709__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2246__S net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4806_ clknet_leaf_17_wb_clk_i _0420_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[76\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2213__A0 net20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2439__S1 _0831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2998_ _1332_ vssd1 vssd1 vccd1 vccd1 _0109_ sky130_fd_sc_hd__clkbuf_1
X_4737_ clknet_leaf_28_wb_clk_i _0351_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[58\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_4668_ clknet_leaf_2_wb_clk_i _0289_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[3\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_3619_ _1588_ tms1x00.RAM\[63\]\[1\] _1693_ vssd1 vssd1 vccd1 vccd1 _1695_ sky130_fd_sc_hd__mux2_1
X_4599_ clknet_leaf_13_wb_clk_i _0220_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[125\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2683__B_N _0788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3495__B _1344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3952__A0 tms1x00.Y\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2755__A1 _0786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5014__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2839__B tms1x00.ram_addr_buff\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3970_ _1894_ vssd1 vssd1 vccd1 vccd1 _0519_ sky130_fd_sc_hd__clkbuf_1
XFILLER_50_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2921_ _1282_ vssd1 vssd1 vccd1 vccd1 _0082_ sky130_fd_sc_hd__clkbuf_1
X_2852_ _1236_ vssd1 vssd1 vccd1 vccd1 _1237_ sky130_fd_sc_hd__buf_4
X_2783_ _0940_ _1170_ _1172_ _0806_ vssd1 vssd1 vccd1 vccd1 _1173_ sky130_fd_sc_hd__o211a_1
X_4522_ clknet_leaf_15_wb_clk_i _0143_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[112\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_4453_ clknet_leaf_20_wb_clk_i _0074_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[79\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3404_ _1492_ tms1x00.RAM\[33\]\[3\] _1566_ vssd1 vssd1 vccd1 vccd1 _1570_ sky130_fd_sc_hd__mux2_1
X_4384_ _2175_ vssd1 vssd1 vccd1 vccd1 _0652_ sky130_fd_sc_hd__clkbuf_1
X_3335_ _1485_ tms1x00.RAM\[31\]\[0\] _1531_ vssd1 vssd1 vccd1 vccd1 _1532_ sky130_fd_sc_hd__mux2_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3266_ _1224_ vssd1 vssd1 vccd1 vccd1 _1492_ sky130_fd_sc_hd__buf_2
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5005_ clknet_leaf_20_wb_clk_i _0615_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[16\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_39_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2217_ net22 wbs_o_buff\[17\] _0668_ vssd1 vssd1 vccd1 vccd1 _0676_ sky130_fd_sc_hd__mux2_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3197_ _1450_ vssd1 vssd1 vccd1 vccd1 _0190_ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4681__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5037__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4220__A _0766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2659__B _1049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2673__B1 _0953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4114__B _0747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2823__S1 _0977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4130__A _0701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output74_A net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3153__A1 _1324_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4554__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3120_ tms1x00.RAM\[10\]\[2\] _1331_ _1404_ vssd1 vssd1 vccd1 vccd1 _1407_ sky130_fd_sc_hd__mux2_1
XFILLER_67_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3051_ _1129_ vssd1 vssd1 vccd1 vccd1 _1366_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__2585__A _0850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2664__B1 _0804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4008__C _0752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3953_ _1885_ vssd1 vssd1 vccd1 vccd1 _0511_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__2967__A1 _1235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2904_ _1228_ _0717_ _0728_ vssd1 vssd1 vccd1 vccd1 _1273_ sky130_fd_sc_hd__or3b_4
XFILLER_32_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3884_ _1847_ vssd1 vssd1 vccd1 vccd1 _0480_ sky130_fd_sc_hd__clkbuf_1
X_2835_ _1224_ vssd1 vssd1 vccd1 vccd1 _1225_ sky130_fd_sc_hd__clkbuf_4
X_2766_ tms1x00.RAM\[108\]\[3\] tms1x00.RAM\[109\]\[3\] tms1x00.RAM\[110\]\[3\] tms1x00.RAM\[111\]\[3\]
+ _0931_ _0932_ vssd1 vssd1 vccd1 vccd1 _1156_ sky130_fd_sc_hd__mux4_1
XANTENNA__2814__S1 _0791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4505_ clknet_leaf_16_wb_clk_i _0126_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[97\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_2697_ _0787_ _1087_ _0996_ vssd1 vssd1 vccd1 vccd1 _1088_ sky130_fd_sc_hd__a21o_1
X_4436_ clknet_leaf_16_wb_clk_i _0057_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[99\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2578__S0 _0945_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3144__A1 _1324_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4367_ tms1x00.RAM\[9\]\[0\] _1323_ _2166_ vssd1 vssd1 vccd1 vccd1 _2167_ sky130_fd_sc_hd__mux2_1
XFILLER_59_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3318_ _1521_ vssd1 vssd1 vccd1 vccd1 _0240_ sky130_fd_sc_hd__clkbuf_1
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4298_ _2128_ vssd1 vssd1 vccd1 vccd1 _0613_ sky130_fd_sc_hd__clkbuf_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3249_ _1481_ vssd1 vssd1 vccd1 vccd1 _0211_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__2655__B1 _0977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2750__S0 _0931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2434__S _0826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2958__A1 _1243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4577__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3135__A1 _1324_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2569__S0 _0945_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2609__S _0924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output112_A net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2620_ tms1x00.RAM\[32\]\[1\] tms1x00.RAM\[33\]\[1\] tms1x00.RAM\[34\]\[1\] tms1x00.RAM\[35\]\[1\]
+ _0840_ _0813_ vssd1 vssd1 vccd1 vccd1 _1012_ sky130_fd_sc_hd__mux4_1
XFILLER_9_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3683__B _1345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2551_ _0922_ _0936_ _0941_ _0942_ vssd1 vssd1 vccd1 vccd1 _0943_ sky130_fd_sc_hd__o211ai_1
Xoutput106 net106 vssd1 vssd1 vccd1 vccd1 ram_adrb[2] sky130_fd_sc_hd__buf_2
X_2482_ _0871_ _0872_ _0874_ _0818_ _0819_ vssd1 vssd1 vccd1 vccd1 _0875_ sky130_fd_sc_hd__a221o_1
XFILLER_5_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput139 net139 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[30] sky130_fd_sc_hd__buf_2
Xoutput117 net117 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[10] sky130_fd_sc_hd__buf_2
Xoutput128 net128 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[20] sky130_fd_sc_hd__buf_2
X_4221_ _2084_ vssd1 vssd1 vccd1 vccd1 _0580_ sky130_fd_sc_hd__clkbuf_1
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4152_ _2024_ vssd1 vssd1 vccd1 vccd1 _2025_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4083_ _0744_ _0750_ _1974_ _1975_ vssd1 vssd1 vccd1 vccd1 _1976_ sky130_fd_sc_hd__or4_1
X_3103_ _0717_ _0728_ _0916_ vssd1 vssd1 vccd1 vccd1 _1396_ sky130_fd_sc_hd__nand3b_4
XFILLER_28_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3034_ _1355_ vssd1 vssd1 vccd1 vccd1 _0122_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_20_wb_clk_i_A clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_52_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4985_ clknet_leaf_2_wb_clk_i _0595_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[119\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2254__S net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3062__A0 _1366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3936_ _1876_ vssd1 vssd1 vccd1 vccd1 _0503_ sky130_fd_sc_hd__clkbuf_1
XFILLER_23_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3867_ tms1x00.RAM\[86\]\[2\] _1777_ _1835_ vssd1 vssd1 vccd1 vccd1 _1838_ sky130_fd_sc_hd__mux2_1
X_3798_ _1706_ tms1x00.RAM\[78\]\[1\] _1796_ vssd1 vssd1 vccd1 vccd1 _1798_ sky130_fd_sc_hd__mux2_1
X_2818_ _0944_ _1201_ _1203_ _0821_ _1207_ vssd1 vssd1 vccd1 vccd1 _1208_ sky130_fd_sc_hd__a311o_1
X_2749_ _0787_ _1138_ _0953_ vssd1 vssd1 vccd1 vccd1 _1139_ sky130_fd_sc_hd__a21o_1
XFILLER_11_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4419_ clknet_leaf_26_wb_clk_i _0018_ vssd1 vssd1 vccd1 vccd1 wbs_o_buff\[23\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__2876__A0 _1130_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2628__B1 _0038_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3768__B _1261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_24_wb_clk_i clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_23_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput19 ram_val[14] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2339__S _0726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2619__B1 _0802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4770_ clknet_leaf_18_wb_clk_i _0384_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[67\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4742__CLK clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3721_ _1753_ vssd1 vssd1 vccd1 vccd1 _0411_ sky130_fd_sc_hd__clkbuf_1
X_3652_ _1708_ tms1x00.RAM\[60\]\[2\] _1712_ vssd1 vssd1 vccd1 vccd1 _1715_ sky130_fd_sc_hd__mux2_1
X_3583_ _1129_ vssd1 vssd1 vccd1 vccd1 _1674_ sky130_fd_sc_hd__buf_2
X_2603_ tms1x00.RAM\[6\]\[1\] tms1x00.RAM\[7\]\[1\] _0975_ vssd1 vssd1 vccd1 vccd1
+ _0995_ sky130_fd_sc_hd__mux2_1
X_2534_ _0787_ _0925_ vssd1 vssd1 vccd1 vccd1 _0926_ sky130_fd_sc_hd__nand2_1
XFILLER_69_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2465_ _0773_ _0805_ _0834_ _0835_ _0857_ vssd1 vssd1 vccd1 vccd1 _0858_ sky130_fd_sc_hd__a311o_2
X_4204_ _2068_ _2069_ vssd1 vssd1 vccd1 vccd1 _2070_ sky130_fd_sc_hd__xnor2_1
X_2396_ _0788_ vssd1 vssd1 vccd1 vccd1 _0789_ sky130_fd_sc_hd__buf_4
XFILLER_69_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4135_ _0770_ _1975_ vssd1 vssd1 vccd1 vccd1 _2012_ sky130_fd_sc_hd__or2_1
XFILLER_29_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4066_ net70 _1960_ vssd1 vssd1 vccd1 vccd1 _1963_ sky130_fd_sc_hd__or2_1
XFILLER_25_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3017_ _1344_ _1345_ vssd1 vssd1 vccd1 vccd1 _1346_ sky130_fd_sc_hd__or2_2
XFILLER_36_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4968_ clknet_leaf_8_wb_clk_i _0578_ vssd1 vssd1 vccd1 vccd1 tms1x00.Y\[1\] sky130_fd_sc_hd__dfxtp_2
X_3919_ _1819_ tms1x00.RAM\[92\]\[1\] _1865_ vssd1 vssd1 vccd1 vccd1 _1867_ sky130_fd_sc_hd__mux2_1
X_4899_ clknet_leaf_12_wb_clk_i _0513_ vssd1 vssd1 vccd1 vccd1 tms1x00.ram_addr_buff\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4615__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3274__A0 _1490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4765__CLK clknet_leaf_20_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3453__S _1599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2250_ net3 K_override\[1\] net148 vssd1 vssd1 vccd1 vccd1 _0693_ sky130_fd_sc_hd__mux2_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2181_ net49 vssd1 vssd1 vccd1 vccd1 _0657_ sky130_fd_sc_hd__clkbuf_4
XFILLER_65_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4822_ clknet_leaf_17_wb_clk_i _0436_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[80\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_4753_ clknet_leaf_2_wb_clk_i _0367_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[63\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3568__A1 _1571_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwrapped_tms1x00_149 vssd1 vssd1 vccd1 vccd1 wrapped_tms1x00_149/HI io_oeb[10] sky130_fd_sc_hd__conb_1
X_3704_ tms1x00.RAM\[71\]\[1\] _1672_ _1742_ vssd1 vssd1 vccd1 vccd1 _1744_ sky130_fd_sc_hd__mux2_1
X_4684_ clknet_leaf_5_wb_clk_i _0298_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[45\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_3635_ _0917_ _1283_ vssd1 vssd1 vccd1 vccd1 _1704_ sky130_fd_sc_hd__or2_2
X_3566_ _1663_ vssd1 vssd1 vccd1 vccd1 _0346_ sky130_fd_sc_hd__clkbuf_1
X_2517_ _0771_ _0907_ _0909_ tms1x00.A\[0\] vssd1 vssd1 vccd1 vccd1 _0910_ sky130_fd_sc_hd__a22o_1
XANTENNA__2768__A _0798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3871__B _1344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3497_ _1625_ vssd1 vssd1 vccd1 vccd1 _0315_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4638__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2448_ tms1x00.RAM\[96\]\[0\] tms1x00.RAM\[97\]\[0\] tms1x00.RAM\[98\]\[0\] tms1x00.RAM\[99\]\[0\]
+ _0840_ _0813_ vssd1 vssd1 vccd1 vccd1 _0841_ sky130_fd_sc_hd__mux4_2
XFILLER_69_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2379_ _0747_ _0748_ vssd1 vssd1 vccd1 vccd1 _0772_ sky130_fd_sc_hd__or2_1
XANTENNA__4788__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4118_ _1998_ vssd1 vssd1 vccd1 vccd1 _0563_ sky130_fd_sc_hd__clkbuf_1
XFILLER_29_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5098_ net51 vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__clkbuf_2
X_4049_ _0733_ _0730_ _0763_ _1915_ vssd1 vssd1 vccd1 vccd1 _1950_ sky130_fd_sc_hd__and4_1
XFILLER_44_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3731__A1 _1672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input36_A ram_val[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3972__A net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2773__A2 _1160_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3420_ tms1x00.RAM\[40\]\[0\] _1571_ _1580_ vssd1 vssd1 vccd1 vccd1 _1581_ sky130_fd_sc_hd__mux2_1
X_3351_ _1540_ vssd1 vssd1 vccd1 vccd1 _0254_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__3722__A1 _1672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2302_ wbs_o_buff\[30\] _0699_ vssd1 vssd1 vccd1 vccd1 _0711_ sky130_fd_sc_hd__and2_1
XANTENNA__4930__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3282_ _1501_ vssd1 vssd1 vccd1 vccd1 _0224_ sky130_fd_sc_hd__clkbuf_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5021_ clknet_leaf_21_wb_clk_i _0631_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[15\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2289__A1 net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2233_ _0684_ vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__clkbuf_1
XFILLER_65_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3789__A1 _1775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4805_ clknet_leaf_17_wb_clk_i _0419_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[76\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_22_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4043__A _0718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2997_ tms1x00.RAM\[101\]\[2\] _1331_ _1325_ vssd1 vssd1 vccd1 vccd1 _1332_ sky130_fd_sc_hd__mux2_1
XFILLER_21_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4736_ clknet_leaf_28_wb_clk_i _0350_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[5\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_4667_ clknet_leaf_3_wb_clk_i _0288_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[3\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4460__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3618_ _1694_ vssd1 vssd1 vccd1 vccd1 _0367_ sky130_fd_sc_hd__clkbuf_1
X_4598_ clknet_leaf_13_wb_clk_i _0219_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[125\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3713__A1 _1672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3549_ _1284_ _1337_ vssd1 vssd1 vccd1 vccd1 _1654_ sky130_fd_sc_hd__nor2_2
XFILLER_29_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4803__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4953__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3704__A1 _1672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4128__A _0738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2871__A _1250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2920_ K_override\[3\] net61 _0715_ vssd1 vssd1 vccd1 vccd1 _1282_ sky130_fd_sc_hd__mux2_1
X_2851_ tms1x00.ram_addr_buff\[4\] tms1x00.ram_addr_buff\[5\] tms1x00.ram_addr_buff\[6\]
+ vssd1 vssd1 vccd1 vccd1 _1236_ sky130_fd_sc_hd__or3b_4
XFILLER_31_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2782_ _0783_ _1171_ vssd1 vssd1 vccd1 vccd1 _1172_ sky130_fd_sc_hd__or2_1
X_4521_ clknet_leaf_15_wb_clk_i _0142_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[113\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4452_ clknet_leaf_17_wb_clk_i _0073_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[79\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_3403_ _1569_ vssd1 vssd1 vccd1 vccd1 _0277_ sky130_fd_sc_hd__clkbuf_1
X_4383_ tms1x00.PA\[0\] net99 _2006_ vssd1 vssd1 vccd1 vccd1 _2175_ sky130_fd_sc_hd__mux2_1
XANTENNA__3207__A _1323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3334_ _1249_ _1267_ vssd1 vssd1 vccd1 vccd1 _1531_ sky130_fd_sc_hd__or2_2
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3265_ _1491_ vssd1 vssd1 vccd1 vccd1 _0217_ sky130_fd_sc_hd__clkbuf_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5004_ clknet_leaf_15_wb_clk_i _0614_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[16\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_2216_ _0675_ vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__clkbuf_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3196_ tms1x00.RAM\[121\]\[3\] _1334_ _1446_ vssd1 vssd1 vccd1 vccd1 _1450_ sky130_fd_sc_hd__mux2_1
XFILLER_82_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4826__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4976__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4187__A1 tms1x00.PC\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2198__A0 net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2737__A2 _1126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4719_ clknet_leaf_29_wb_clk_i _0333_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[54\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3816__S _1806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2370__B1 net77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2673__A1 _0818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4178__A1 _0760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4130__B _2006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3050_ _1365_ vssd1 vssd1 vccd1 vccd1 _0128_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_10_wb_clk_i_A clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4849__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2664__A1 _0776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2805__S _0778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3952_ tms1x00.Y\[0\] _0717_ _0726_ vssd1 vssd1 vccd1 vccd1 _1885_ sky130_fd_sc_hd__mux2_1
XFILLER_32_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4999__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2903_ _1272_ vssd1 vssd1 vccd1 vccd1 _0074_ sky130_fd_sc_hd__clkbuf_1
XFILLER_32_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3883_ tms1x00.RAM\[88\]\[1\] _1775_ _1845_ vssd1 vssd1 vccd1 vccd1 _1847_ sky130_fd_sc_hd__mux2_1
XANTENNA__4169__A1 tms1x00.PC\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2834_ _1223_ vssd1 vssd1 vccd1 vccd1 _1224_ sky130_fd_sc_hd__clkbuf_4
X_4504_ clknet_leaf_16_wb_clk_i _0125_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[97\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_2765_ _0920_ _1135_ _1141_ _1154_ _0773_ vssd1 vssd1 vccd1 vccd1 _1155_ sky130_fd_sc_hd__o311a_1
XANTENNA__4321__A _1267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2696_ tms1x00.RAM\[92\]\[2\] tms1x00.RAM\[93\]\[2\] _0975_ vssd1 vssd1 vccd1 vccd1
+ _1087_ sky130_fd_sc_hd__mux2_1
X_4435_ clknet_leaf_16_wb_clk_i _0056_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[99\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2578__S1 _0956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4366_ _1261_ _1344_ vssd1 vssd1 vccd1 vccd1 _2166_ sky130_fd_sc_hd__nor2_2
XFILLER_59_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3317_ tms1x00.RAM\[26\]\[1\] _1459_ _1519_ vssd1 vssd1 vccd1 vccd1 _1521_ sky130_fd_sc_hd__mux2_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4297_ _1819_ tms1x00.RAM\[16\]\[1\] _2126_ vssd1 vssd1 vccd1 vccd1 _2128_ sky130_fd_sc_hd__mux2_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3248_ _1361_ tms1x00.RAM\[115\]\[0\] _1480_ vssd1 vssd1 vccd1 vccd1 _1481_ sky130_fd_sc_hd__mux2_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2655__A1 _0975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3179_ _1440_ vssd1 vssd1 vccd1 vccd1 _0182_ sky130_fd_sc_hd__clkbuf_1
XFILLER_26_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2750__S1 _0932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2569__S1 _0791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4377__S _2006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output105_A net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2550_ _0802_ vssd1 vssd1 vccd1 vccd1 _0942_ sky130_fd_sc_hd__clkbuf_4
XFILLER_5_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput107 net107 vssd1 vssd1 vccd1 vccd1 ram_adrb[3] sky130_fd_sc_hd__buf_2
X_2481_ tms1x00.RAM\[12\]\[0\] tms1x00.RAM\[13\]\[0\] _0873_ vssd1 vssd1 vccd1 vccd1
+ _0874_ sky130_fd_sc_hd__mux2_1
XFILLER_5_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput118 net118 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[11] sky130_fd_sc_hd__buf_2
Xoutput129 net129 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[21] sky130_fd_sc_hd__buf_2
X_4220_ _0766_ _2083_ vssd1 vssd1 vccd1 vccd1 _2084_ sky130_fd_sc_hd__and2_1
XFILLER_5_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4151_ _0701_ _0720_ tms1x00.PC\[0\] vssd1 vssd1 vccd1 vccd1 _2024_ sky130_fd_sc_hd__and3b_1
XANTENNA__2596__A _0818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3102_ _1395_ vssd1 vssd1 vccd1 vccd1 _0150_ sky130_fd_sc_hd__clkbuf_1
X_4082_ tms1x00.ins_in\[1\] tms1x00.ins_in\[0\] vssd1 vssd1 vccd1 vccd1 _1975_ sky130_fd_sc_hd__nand2_1
X_3033_ _1225_ tms1x00.RAM\[98\]\[3\] _1351_ vssd1 vssd1 vccd1 vccd1 _1355_ sky130_fd_sc_hd__mux2_1
XFILLER_49_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2637__A1 _0040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5027__CLK clknet_leaf_20_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4984_ clknet_leaf_2_wb_clk_i _0594_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[119\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3220__A _1317_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4035__B _0730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3935_ tms1x00.RAM\[90\]\[0\] _1323_ _1875_ vssd1 vssd1 vccd1 vccd1 _1876_ sky130_fd_sc_hd__mux2_1
XFILLER_20_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3866_ _1837_ vssd1 vssd1 vccd1 vccd1 _0472_ sky130_fd_sc_hd__clkbuf_1
X_3797_ _1797_ vssd1 vssd1 vccd1 vccd1 _0443_ sky130_fd_sc_hd__clkbuf_1
X_2817_ _0940_ _1204_ _1206_ _0806_ vssd1 vssd1 vccd1 vccd1 _1207_ sky130_fd_sc_hd__o211a_1
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2748_ tms1x00.RAM\[92\]\[3\] tms1x00.RAM\[93\]\[3\] _0789_ vssd1 vssd1 vccd1 vccd1
+ _1138_ sky130_fd_sc_hd__mux2_1
X_2679_ _0785_ _1069_ _0793_ vssd1 vssd1 vccd1 vccd1 _1070_ sky130_fd_sc_hd__a21o_1
X_4418_ clknet_leaf_26_wb_clk_i _0017_ vssd1 vssd1 vccd1 vccd1 wbs_o_buff\[22\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__2350__A_N net76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4349_ _1235_ tms1x00.RAM\[13\]\[0\] _2156_ vssd1 vssd1 vccd1 vccd1 _2157_ sky130_fd_sc_hd__mux2_1
XTAP_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2628__A1 _0794_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2487__S0 _0830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4544__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4694__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input66_A wbs_dat_i[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3305__A _1250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2619__A1 _0807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3292__A1 _1461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3975__A net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3720_ tms1x00.RAM\[6\]\[0\] _1669_ _1752_ vssd1 vssd1 vccd1 vccd1 _1753_ sky130_fd_sc_hd__mux2_1
XFILLER_41_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3651_ _1714_ vssd1 vssd1 vccd1 vccd1 _0380_ sky130_fd_sc_hd__clkbuf_1
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3582_ _1673_ vssd1 vssd1 vccd1 vccd1 _0352_ sky130_fd_sc_hd__clkbuf_1
X_2602_ tms1x00.RAM\[4\]\[1\] tms1x00.RAM\[5\]\[1\] _0924_ vssd1 vssd1 vccd1 vccd1
+ _0994_ sky130_fd_sc_hd__mux2_1
XFILLER_6_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2533_ tms1x00.RAM\[68\]\[1\] tms1x00.RAM\[69\]\[1\] _0924_ vssd1 vssd1 vccd1 vccd1
+ _0925_ sky130_fd_sc_hd__mux2_1
XANTENNA__2650__S0 _0955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2464_ _0821_ _0839_ _0844_ _0856_ _0040_ vssd1 vssd1 vccd1 vccd1 _0857_ sky130_fd_sc_hd__o311a_1
XFILLER_69_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4203_ tms1x00.P\[0\] _2059_ _2060_ vssd1 vssd1 vccd1 vccd1 _2069_ sky130_fd_sc_hd__a21bo_1
X_2395_ _0777_ vssd1 vssd1 vccd1 vccd1 _0788_ sky130_fd_sc_hd__buf_6
XFILLER_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4134_ _0701_ _2006_ vssd1 vssd1 vccd1 vccd1 _2011_ sky130_fd_sc_hd__or2_1
XANTENNA__3807__A0 _1706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4065_ _0742_ tms1x00.A\[1\] vssd1 vssd1 vccd1 vccd1 _1962_ sky130_fd_sc_hd__and2b_1
XFILLER_49_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3016_ _0717_ _0728_ _1228_ vssd1 vssd1 vccd1 vccd1 _1345_ sky130_fd_sc_hd__or3_4
XFILLER_37_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3283__A1 _1461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4967_ clknet_leaf_8_wb_clk_i _0577_ vssd1 vssd1 vccd1 vccd1 tms1x00.Y\[0\] sky130_fd_sc_hd__dfxtp_2
X_3918_ _1866_ vssd1 vssd1 vccd1 vccd1 _0495_ sky130_fd_sc_hd__clkbuf_1
X_4898_ clknet_leaf_3_wb_clk_i _0512_ vssd1 vssd1 vccd1 vccd1 tms1x00.ram_addr_buff\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3849_ _1821_ tms1x00.RAM\[82\]\[2\] _1825_ vssd1 vssd1 vccd1 vccd1 _1828_ sky130_fd_sc_hd__mux2_1
XANTENNA__3991__C1 _1901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2546__B1 _0932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4299__A0 _1821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3125__A _0913_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2482__C1 _0819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3795__A _1236_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3982__C1 _1901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2785__B1 _0040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2204__A _0669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3035__A _0913_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2180_ _0656_ vssd1 vssd1 vccd1 vccd1 valid sky130_fd_sc_hd__clkbuf_2
XFILLER_66_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4821_ clknet_leaf_18_wb_clk_i _0435_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[80\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_34_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4752_ clknet_leaf_28_wb_clk_i _0366_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[55\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_4683_ clknet_leaf_5_wb_clk_i _0297_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[45\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_3703_ _1743_ vssd1 vssd1 vccd1 vccd1 _0403_ sky130_fd_sc_hd__clkbuf_1
X_3634_ _0911_ vssd1 vssd1 vccd1 vccd1 _1703_ sky130_fd_sc_hd__clkbuf_4
X_3565_ _1592_ tms1x00.RAM\[51\]\[3\] _1659_ vssd1 vssd1 vccd1 vccd1 _1663_ sky130_fd_sc_hd__mux2_1
X_2516_ _0771_ _0908_ vssd1 vssd1 vccd1 vccd1 _0909_ sky130_fd_sc_hd__and2b_1
XANTENNA__2768__B _1157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3496_ tms1x00.RAM\[4\]\[0\] _1571_ _1624_ vssd1 vssd1 vccd1 vccd1 _1625_ sky130_fd_sc_hd__mux2_1
X_2447_ _0815_ vssd1 vssd1 vccd1 vccd1 _0840_ sky130_fd_sc_hd__buf_8
XFILLER_57_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2378_ _0738_ _0760_ _0767_ _0770_ vssd1 vssd1 vccd1 vccd1 _0771_ sky130_fd_sc_hd__or4_2
XFILLER_29_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4117_ net103 _1997_ vssd1 vssd1 vccd1 vccd1 _1998_ sky130_fd_sc_hd__or2_1
X_5097_ net50 vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__clkbuf_2
XFILLER_17_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4048_ _0753_ _1948_ _1949_ _1931_ vssd1 vssd1 vccd1 vccd1 _0542_ sky130_fd_sc_hd__o211a_1
XFILLER_56_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2464__C1 _0040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4205__A0 tms1x00.Y\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3008__A1 _1328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4732__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4385__S _2006_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input29_A ram_val[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4882__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2869__A _1249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output97_A net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3350_ _1492_ tms1x00.RAM\[30\]\[3\] _1536_ vssd1 vssd1 vccd1 vccd1 _1540_ sky130_fd_sc_hd__mux2_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2301_ _0710_ vssd1 vssd1 vccd1 vccd1 _0024_ sky130_fd_sc_hd__clkbuf_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3281_ tms1x00.RAM\[25\]\[1\] _1459_ _1499_ vssd1 vssd1 vccd1 vccd1 _1501_ sky130_fd_sc_hd__mux2_1
X_5020_ clknet_leaf_21_wb_clk_i _0630_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[15\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_66_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2289__A2 _0697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2232_ net30 wbs_o_buff\[24\] _0679_ vssd1 vssd1 vccd1 vccd1 _0684_ sky130_fd_sc_hd__mux2_1
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2446__C1 _0802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4804_ clknet_leaf_24_wb_clk_i _0418_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[68\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2749__B1 _0953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4735_ clknet_leaf_28_wb_clk_i _0349_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[5\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2996_ _1330_ vssd1 vssd1 vccd1 vccd1 _1331_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__4605__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4666_ clknet_leaf_3_wb_clk_i _0287_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[3\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_4597_ clknet_leaf_12_wb_clk_i _0218_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[126\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2779__A _0921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3617_ _1585_ tms1x00.RAM\[63\]\[0\] _1693_ vssd1 vssd1 vccd1 vccd1 _1694_ sky130_fd_sc_hd__mux2_1
X_3548_ _1653_ vssd1 vssd1 vccd1 vccd1 _0338_ sky130_fd_sc_hd__clkbuf_1
XFILLER_77_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3479_ _1615_ vssd1 vssd1 vccd1 vccd1 _0307_ sky130_fd_sc_hd__clkbuf_1
XFILLER_76_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3165__A0 _1364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2912__A0 _1225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4128__B _0760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4628__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2871__B _1251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2850_ _0911_ vssd1 vssd1 vccd1 vccd1 _1235_ sky130_fd_sc_hd__clkbuf_4
XFILLER_31_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2826__S0 _0826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2781_ tms1x00.RAM\[120\]\[3\] tms1x00.RAM\[121\]\[3\] tms1x00.RAM\[122\]\[3\] tms1x00.RAM\[123\]\[3\]
+ _0823_ _0850_ vssd1 vssd1 vccd1 vccd1 _1171_ sky130_fd_sc_hd__mux4_1
X_4520_ clknet_leaf_16_wb_clk_i _0141_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[113\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2600__C1 _0806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4451_ clknet_leaf_17_wb_clk_i _0072_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[79\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3402_ _1490_ tms1x00.RAM\[33\]\[2\] _1566_ vssd1 vssd1 vccd1 vccd1 _1569_ sky130_fd_sc_hd__mux2_1
X_4382_ _2174_ vssd1 vssd1 vccd1 vccd1 _0651_ sky130_fd_sc_hd__clkbuf_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3333_ _1530_ vssd1 vssd1 vccd1 vccd1 _0246_ sky130_fd_sc_hd__clkbuf_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3264_ _1490_ tms1x00.RAM\[126\]\[2\] _1486_ vssd1 vssd1 vccd1 vccd1 _1491_ sky130_fd_sc_hd__mux2_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5003_ clknet_leaf_12_wb_clk_i _0613_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[16\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_38_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2215_ net21 wbs_o_buff\[16\] _0668_ vssd1 vssd1 vccd1 vccd1 _0675_ sky130_fd_sc_hd__mux2_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3195_ _1449_ vssd1 vssd1 vccd1 vccd1 _0189_ sky130_fd_sc_hd__clkbuf_1
XFILLER_82_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4038__B _0730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3395__A0 _1492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2198__A1 wbs_o_buff\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2979_ _1319_ vssd1 vssd1 vccd1 vccd1 _0103_ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4718_ clknet_leaf_29_wb_clk_i _0332_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[54\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_4649_ clknet_leaf_8_wb_clk_i _0270_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[35\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_18_wb_clk_i clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_29_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4920__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3386__A0 _1492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2649__C1 _0942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4450__CLK clknet_leaf_20_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_6_wb_clk_i_A clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__3978__A net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2882__A tms1x00.ram_addr_buff\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3951_ _1884_ vssd1 vssd1 vccd1 vccd1 _0510_ sky130_fd_sc_hd__clkbuf_1
XFILLER_17_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2902_ _1225_ tms1x00.RAM\[79\]\[3\] _1268_ vssd1 vssd1 vccd1 vccd1 _1272_ sky130_fd_sc_hd__mux2_1
XFILLER_16_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3882_ _1846_ vssd1 vssd1 vccd1 vccd1 _0479_ sky130_fd_sc_hd__clkbuf_1
X_2833_ tms1x00.A\[3\] _0909_ _1221_ _1222_ vssd1 vssd1 vccd1 vccd1 _1223_ sky130_fd_sc_hd__a22o_1
XFILLER_32_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2764_ _0821_ _1147_ _1153_ vssd1 vssd1 vccd1 vccd1 _1154_ sky130_fd_sc_hd__or3_1
XANTENNA__2821__S _0975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4503_ clknet_leaf_16_wb_clk_i _0124_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[97\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4321__B _1375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2695_ _0928_ _1085_ vssd1 vssd1 vccd1 vccd1 _1086_ sky130_fd_sc_hd__and2_1
X_4434_ clknet_leaf_17_wb_clk_i _0055_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[99\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_4365_ _2165_ vssd1 vssd1 vccd1 vccd1 _0643_ sky130_fd_sc_hd__clkbuf_1
X_3316_ _1520_ vssd1 vssd1 vccd1 vccd1 _0239_ sky130_fd_sc_hd__clkbuf_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4296_ _2127_ vssd1 vssd1 vccd1 vccd1 _0612_ sky130_fd_sc_hd__clkbuf_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3247_ _1229_ _1375_ vssd1 vssd1 vccd1 vccd1 _1480_ sky130_fd_sc_hd__or2_2
XANTENNA__3301__A0 _1490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3178_ tms1x00.RAM\[123\]\[3\] _1334_ _1436_ vssd1 vssd1 vccd1 vccd1 _1440_ sky130_fd_sc_hd__mux2_1
XFILLER_54_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3827__S _1811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4473__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input11_A oram_value[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3359__A0 _1492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2480_ _0815_ vssd1 vssd1 vccd1 vccd1 _0873_ sky130_fd_sc_hd__buf_6
Xoutput119 net119 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[12] sky130_fd_sc_hd__buf_2
Xoutput108 net108 vssd1 vssd1 vccd1 vccd1 ram_adrb[4] sky130_fd_sc_hd__buf_2
XFILLER_68_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4150_ tms1x00.P\[3\] _2007_ _2021_ _2023_ vssd1 vssd1 vccd1 vccd1 _0570_ sky130_fd_sc_hd__o22a_1
Xoutput90 net90 vssd1 vssd1 vccd1 vccd1 io_out[31] sky130_fd_sc_hd__buf_2
X_3101_ _1368_ tms1x00.RAM\[111\]\[3\] _1391_ vssd1 vssd1 vccd1 vccd1 _1395_ sky130_fd_sc_hd__mux2_1
XFILLER_1_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4081_ _0760_ _1971_ vssd1 vssd1 vccd1 vccd1 _1974_ sky130_fd_sc_hd__or2_1
X_3032_ _1354_ vssd1 vssd1 vccd1 vccd1 _0121_ sky130_fd_sc_hd__clkbuf_1
XFILLER_49_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4983_ clknet_leaf_2_wb_clk_i _0593_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[119\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3220__B _1430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3934_ _1258_ _1403_ vssd1 vssd1 vccd1 vccd1 _1875_ sky130_fd_sc_hd__nor2_2
XFILLER_32_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3865_ tms1x00.RAM\[86\]\[1\] _1775_ _1835_ vssd1 vssd1 vccd1 vccd1 _1837_ sky130_fd_sc_hd__mux2_1
X_2816_ _0783_ _1205_ vssd1 vssd1 vccd1 vccd1 _1206_ sky130_fd_sc_hd__or2_1
XFILLER_31_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3796_ _1703_ tms1x00.RAM\[78\]\[0\] _1796_ vssd1 vssd1 vccd1 vccd1 _1797_ sky130_fd_sc_hd__mux2_1
X_2747_ _0928_ _1136_ vssd1 vssd1 vccd1 vccd1 _1137_ sky130_fd_sc_hd__and2_1
XFILLER_11_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2678_ tms1x00.RAM\[4\]\[2\] tms1x00.RAM\[5\]\[2\] _0823_ vssd1 vssd1 vccd1 vccd1
+ _1069_ sky130_fd_sc_hd__mux2_1
X_4417_ clknet_leaf_27_wb_clk_i _0016_ vssd1 vssd1 vccd1 vccd1 wbs_o_buff\[21\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_input3_A io_in[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4348_ _0917_ _1343_ vssd1 vssd1 vccd1 vccd1 _2156_ sky130_fd_sc_hd__or2_2
X_4279_ _1819_ tms1x00.RAM\[29\]\[1\] _2116_ vssd1 vssd1 vccd1 vccd1 _2118_ sky130_fd_sc_hd__mux2_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3825__A1 _1775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4250__A1 _1323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2487__S1 _0831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input59_A wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_33_wb_clk_i clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_33_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__4989__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3305__B _1286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3816__A1 _1775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3650_ _1706_ tms1x00.RAM\[60\]\[1\] _1712_ vssd1 vssd1 vccd1 vccd1 _1714_ sky130_fd_sc_hd__mux2_1
X_2601_ _0944_ _0986_ _0992_ _0920_ vssd1 vssd1 vccd1 vccd1 _0993_ sky130_fd_sc_hd__a211oi_1
X_3581_ tms1x00.RAM\[58\]\[1\] _1672_ _1670_ vssd1 vssd1 vccd1 vccd1 _1673_ sky130_fd_sc_hd__mux2_1
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2532_ _0923_ vssd1 vssd1 vccd1 vccd1 _0924_ sky130_fd_sc_hd__buf_6
XANTENNA__2650__S1 _0956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4202_ _2066_ _2067_ vssd1 vssd1 vccd1 vccd1 _2068_ sky130_fd_sc_hd__nand2_1
X_2463_ _0846_ _0848_ _0853_ _0855_ _0804_ vssd1 vssd1 vccd1 vccd1 _0856_ sky130_fd_sc_hd__a221o_1
XFILLER_69_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2394_ _0786_ vssd1 vssd1 vccd1 vccd1 _0787_ sky130_fd_sc_hd__buf_4
X_4133_ _2008_ _2009_ vssd1 vssd1 vccd1 vccd1 _2010_ sky130_fd_sc_hd__nor2_1
X_4064_ _1958_ _1959_ _1961_ _1931_ vssd1 vssd1 vccd1 vccd1 _0546_ sky130_fd_sc_hd__o211a_1
XFILLER_56_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3015_ _1343_ vssd1 vssd1 vccd1 vccd1 _1344_ sky130_fd_sc_hd__buf_6
XFILLER_52_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4966_ clknet_leaf_7_wb_clk_i _0576_ vssd1 vssd1 vccd1 vccd1 tms1x00.PC\[5\] sky130_fd_sc_hd__dfxtp_1
X_3917_ _1816_ tms1x00.RAM\[92\]\[0\] _1865_ vssd1 vssd1 vccd1 vccd1 _1866_ sky130_fd_sc_hd__mux2_1
X_4897_ clknet_leaf_3_wb_clk_i _0511_ vssd1 vssd1 vccd1 vccd1 tms1x00.ram_addr_buff\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3848_ _1827_ vssd1 vssd1 vccd1 vccd1 _0464_ sky130_fd_sc_hd__clkbuf_1
XFILLER_20_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3779_ _1787_ vssd1 vssd1 vccd1 vccd1 _0435_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__2546__A1 _0924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3406__A _0911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3125__B _1409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3795__B _1396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2234__A0 net31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2785__A1 _0821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3982__B1 _1902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5017__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3035__B _1251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3051__A _1129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3986__A net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4820_ clknet_leaf_24_wb_clk_i _0434_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[73\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_4751_ clknet_leaf_21_wb_clk_i _0365_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[55\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_4682_ clknet_leaf_4_wb_clk_i _0296_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[45\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_3702_ tms1x00.RAM\[71\]\[0\] _1669_ _1742_ vssd1 vssd1 vccd1 vccd1 _1743_ sky130_fd_sc_hd__mux2_1
X_3633_ _1702_ vssd1 vssd1 vccd1 vccd1 _0374_ sky130_fd_sc_hd__clkbuf_1
X_3564_ _1662_ vssd1 vssd1 vccd1 vccd1 _0345_ sky130_fd_sc_hd__clkbuf_1
X_2515_ tms1x00.ins_in\[1\] _0742_ vssd1 vssd1 vccd1 vccd1 _0908_ sky130_fd_sc_hd__nor2_1
X_3495_ _1337_ _1344_ vssd1 vssd1 vccd1 vccd1 _1624_ sky130_fd_sc_hd__nor2_2
X_2446_ _0819_ _0836_ _0838_ _0802_ vssd1 vssd1 vccd1 vccd1 _0839_ sky130_fd_sc_hd__o211a_1
XFILLER_69_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2377_ tms1x00.ins_in\[3\] _0768_ _0769_ vssd1 vssd1 vccd1 vccd1 _0770_ sky130_fd_sc_hd__or3b_1
X_4116_ tms1x00.PB\[0\] tms1x00.PA\[0\] _1996_ vssd1 vssd1 vccd1 vccd1 _1997_ sky130_fd_sc_hd__mux2_1
XFILLER_57_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4047_ _0764_ _1947_ net89 vssd1 vssd1 vccd1 vccd1 _1949_ sky130_fd_sc_hd__a21o_1
XFILLER_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4684__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4949_ clknet_leaf_6_wb_clk_i _0559_ vssd1 vssd1 vccd1 vccd1 tms1x00.PB\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_33_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3192__A1 _1328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2455__B1 _0038_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2914__S _0715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2207__A0 net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3183__A1 _1328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3280_ _1500_ vssd1 vssd1 vccd1 vccd1 _0223_ sky130_fd_sc_hd__clkbuf_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2300_ wbs_o_buff\[29\] _0704_ vssd1 vssd1 vccd1 vccd1 _0710_ sky130_fd_sc_hd__and2_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2231_ _0683_ vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__clkbuf_1
XFILLER_2_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2885__A _1258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2541__S0 _0931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2997__A1 _1331_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4803_ clknet_leaf_22_wb_clk_i _0417_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[68\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2749__A1 _0787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2995_ _1128_ vssd1 vssd1 vccd1 vccd1 _1330_ sky130_fd_sc_hd__clkbuf_4
X_4734_ clknet_leaf_28_wb_clk_i _0348_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[5\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4665_ clknet_leaf_27_wb_clk_i _0286_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[40\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_4596_ clknet_leaf_10_wb_clk_i _0217_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[126\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_3616_ _1267_ _1283_ vssd1 vssd1 vccd1 vccd1 _1693_ sky130_fd_sc_hd__or2_2
XANTENNA__3174__A1 _1328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3547_ tms1x00.RAM\[53\]\[3\] _1578_ _1649_ vssd1 vssd1 vccd1 vccd1 _1653_ sky130_fd_sc_hd__mux2_1
X_3478_ tms1x00.RAM\[42\]\[0\] _1571_ _1614_ vssd1 vssd1 vccd1 vccd1 _1615_ sky130_fd_sc_hd__mux2_1
X_2429_ _0812_ vssd1 vssd1 vccd1 vccd1 _0822_ sky130_fd_sc_hd__buf_6
XANTENNA__2780__S0 _0923_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4234__B _2007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3937__A0 tms1x00.RAM\[90\]\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2599__S0 _0945_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4362__A0 _1245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input41_A ram_val[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2771__S0 _0873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2780_ tms1x00.RAM\[124\]\[3\] tms1x00.RAM\[125\]\[3\] tms1x00.RAM\[126\]\[3\] tms1x00.RAM\[127\]\[3\]
+ _0923_ _0927_ vssd1 vssd1 vccd1 vccd1 _1170_ sky130_fd_sc_hd__mux4_1
XANTENNA__2826__S1 _0850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2600__B1 _0991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4450_ clknet_leaf_20_wb_clk_i _0071_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[79\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3401_ _1568_ vssd1 vssd1 vccd1 vccd1 _0276_ sky130_fd_sc_hd__clkbuf_1
X_4381_ tms1x00.PC\[5\] net98 _2006_ vssd1 vssd1 vccd1 vccd1 _2174_ sky130_fd_sc_hd__mux2_1
XANTENNA__4353__A0 _1245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3332_ _1492_ tms1x00.RAM\[32\]\[3\] _1526_ vssd1 vssd1 vccd1 vccd1 _1530_ sky130_fd_sc_hd__mux2_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3263_ _1129_ vssd1 vssd1 vccd1 vccd1 _1490_ sky130_fd_sc_hd__buf_2
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5002_ clknet_leaf_12_wb_clk_i _0612_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[16\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3504__A _1284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2214_ _0674_ vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__clkbuf_1
X_3194_ tms1x00.RAM\[121\]\[2\] _1331_ _1446_ vssd1 vssd1 vccd1 vccd1 _1449_ sky130_fd_sc_hd__mux2_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3092__A0 _1368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3919__A0 _1819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4722__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2978_ tms1x00.RAM\[102\]\[0\] _1235_ _1318_ vssd1 vssd1 vccd1 vccd1 _1319_ sky130_fd_sc_hd__mux2_1
XFILLER_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4717_ clknet_leaf_29_wb_clk_i _0331_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[54\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_4648_ clknet_leaf_6_wb_clk_i _0269_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[35\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4070__A _0718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4344__A0 _1245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4579_ clknet_leaf_2_wb_clk_i _0200_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[118\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2302__B _0699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3083__A0 _1368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4335__A0 _1245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4139__B _1030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3310__A1 _1461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3074__A0 _1368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3950_ tms1x00.RAM\[23\]\[3\] _1333_ _1880_ vssd1 vssd1 vccd1 vccd1 _1884_ sky130_fd_sc_hd__mux2_1
XFILLER_17_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2901_ _1271_ vssd1 vssd1 vccd1 vccd1 _0073_ sky130_fd_sc_hd__clkbuf_1
XFILLER_32_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4745__CLK clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3994__A _0701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3881_ tms1x00.RAM\[88\]\[0\] _1772_ _1845_ vssd1 vssd1 vccd1 vccd1 _1846_ sky130_fd_sc_hd__mux2_1
XANTENNA__4023__C1 _1931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2832_ _0747_ _0748_ vssd1 vssd1 vccd1 vccd1 _1222_ sky130_fd_sc_hd__nand2_1
X_2763_ _0798_ _1148_ _1152_ _0802_ vssd1 vssd1 vccd1 vccd1 _1153_ sky130_fd_sc_hd__o211a_1
XANTENNA__4895__CLK clknet_leaf_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3377__A1 _1463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4502_ clknet_leaf_16_wb_clk_i _0123_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[97\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4326__A0 _1821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2694_ tms1x00.RAM\[94\]\[2\] tms1x00.RAM\[95\]\[2\] _0789_ vssd1 vssd1 vccd1 vccd1
+ _1085_ sky130_fd_sc_hd__mux2_1
XFILLER_8_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4433_ clknet_leaf_14_wb_clk_i _0054_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[109\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4364_ _1247_ tms1x00.RAM\[14\]\[3\] _2161_ vssd1 vssd1 vccd1 vccd1 _2165_ sky130_fd_sc_hd__mux2_1
XFILLER_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4295_ _1816_ tms1x00.RAM\[16\]\[0\] _2126_ vssd1 vssd1 vccd1 vccd1 _2127_ sky130_fd_sc_hd__mux2_1
X_3315_ tms1x00.RAM\[26\]\[0\] _1456_ _1519_ vssd1 vssd1 vccd1 vccd1 _1520_ sky130_fd_sc_hd__mux2_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3246_ _1479_ vssd1 vssd1 vccd1 vccd1 _0210_ sky130_fd_sc_hd__clkbuf_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4049__B _0730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3177_ _1439_ vssd1 vssd1 vccd1 vccd1 _0181_ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3368__A1 _1463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2576__C1 _0942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4317__A0 _1821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2459__S _0788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4618__CLK clknet_leaf_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4768__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4005__C1 _1901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2567__C1 _0920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2223__A net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput109 net109 vssd1 vssd1 vccd1 vccd1 ram_adrb[5] sky130_fd_sc_hd__buf_2
XANTENNA_output72_A net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput91 net91 vssd1 vssd1 vccd1 vccd1 io_out[32] sky130_fd_sc_hd__buf_2
Xoutput80 net80 vssd1 vssd1 vccd1 vccd1 io_out[21] sky130_fd_sc_hd__buf_2
XFILLER_68_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3100_ _1394_ vssd1 vssd1 vccd1 vccd1 _0149_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__3054__A _1224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4080_ tms1x00.status _0747_ _0748_ _1972_ vssd1 vssd1 vccd1 vccd1 _1973_ sky130_fd_sc_hd__and4_2
X_3031_ _1130_ tms1x00.RAM\[98\]\[2\] _1351_ vssd1 vssd1 vccd1 vccd1 _1354_ sky130_fd_sc_hd__mux2_1
XFILLER_48_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4982_ clknet_leaf_2_wb_clk_i _0592_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[119\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_3_wb_clk_i clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_16_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3933_ _1874_ vssd1 vssd1 vccd1 vccd1 _0502_ sky130_fd_sc_hd__clkbuf_1
X_3864_ _1836_ vssd1 vssd1 vccd1 vccd1 _0471_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__2270__B2 wbs_o_buff\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2270__A1 net76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2815_ tms1x00.RAM\[40\]\[3\] tms1x00.RAM\[41\]\[3\] tms1x00.RAM\[42\]\[3\] tms1x00.RAM\[43\]\[3\]
+ _0826_ _0780_ vssd1 vssd1 vccd1 vccd1 _1205_ sky130_fd_sc_hd__mux4_1
X_3795_ _1236_ _1396_ vssd1 vssd1 vccd1 vccd1 _1796_ sky130_fd_sc_hd__or2_2
XANTENNA__3229__A _1240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2746_ tms1x00.RAM\[94\]\[3\] tms1x00.RAM\[95\]\[3\] _0923_ vssd1 vssd1 vccd1 vccd1
+ _1136_ sky130_fd_sc_hd__mux2_1
XFILLER_11_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2677_ _0813_ _1067_ vssd1 vssd1 vccd1 vccd1 _1068_ sky130_fd_sc_hd__and2_1
X_4416_ clknet_leaf_27_wb_clk_i _0015_ vssd1 vssd1 vccd1 vccd1 wbs_o_buff\[20\] sky130_fd_sc_hd__dfxtp_1
X_4347_ _2155_ vssd1 vssd1 vccd1 vccd1 _0635_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4910__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4278_ _2117_ vssd1 vssd1 vccd1 vccd1 _0604_ sky130_fd_sc_hd__clkbuf_1
XTAP_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3229_ _1240_ _1430_ vssd1 vssd1 vccd1 vccd1 _1470_ sky130_fd_sc_hd__nor2_2
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3038__A0 _1035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2308__A net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2549__C1 _0940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4440__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3029__A0 _1035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output110_A net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2252__A1 K_override\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2600_ _0988_ _0990_ _0991_ _0948_ _0806_ vssd1 vssd1 vccd1 vccd1 _0992_ sky130_fd_sc_hd__o221a_1
X_3580_ _1034_ vssd1 vssd1 vccd1 vccd1 _1672_ sky130_fd_sc_hd__clkbuf_4
X_2531_ _0826_ vssd1 vssd1 vccd1 vccd1 _0923_ sky130_fd_sc_hd__buf_6
X_4201_ tms1x00.P\[1\] tms1x00.N\[1\] vssd1 vssd1 vccd1 vccd1 _2067_ sky130_fd_sc_hd__or2_1
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2462_ _0797_ _0854_ _0774_ vssd1 vssd1 vccd1 vccd1 _0855_ sky130_fd_sc_hd__o21a_1
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2393_ _0785_ vssd1 vssd1 vccd1 vccd1 _0786_ sky130_fd_sc_hd__clkbuf_4
XFILLER_68_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4132_ _0743_ _0768_ _0769_ _0908_ vssd1 vssd1 vccd1 vccd1 _2009_ sky130_fd_sc_hd__and4_1
XFILLER_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4063_ net69 _1960_ vssd1 vssd1 vccd1 vccd1 _1961_ sky130_fd_sc_hd__or2_1
XFILLER_56_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3014_ tms1x00.ram_addr_buff\[4\] tms1x00.ram_addr_buff\[5\] tms1x00.ram_addr_buff\[6\]
+ vssd1 vssd1 vccd1 vccd1 _1343_ sky130_fd_sc_hd__or3_4
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4965_ clknet_leaf_6_wb_clk_i _0575_ vssd1 vssd1 vccd1 vccd1 tms1x00.PC\[4\] sky130_fd_sc_hd__dfxtp_2
XFILLER_24_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3916_ _1257_ _1409_ vssd1 vssd1 vccd1 vccd1 _1865_ sky130_fd_sc_hd__or2_2
XFILLER_60_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4896_ clknet_leaf_0_wb_clk_i _0510_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[23\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3991__A1 _0747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3847_ _1819_ tms1x00.RAM\[82\]\[1\] _1825_ vssd1 vssd1 vccd1 vccd1 _1827_ sky130_fd_sc_hd__mux2_1
XANTENNA__4463__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3778_ _1703_ tms1x00.RAM\[80\]\[0\] _1786_ vssd1 vssd1 vccd1 vccd1 _1787_ sky130_fd_sc_hd__mux2_1
X_2729_ tms1x00.RAM\[108\]\[2\] tms1x00.RAM\[109\]\[2\] tms1x00.RAM\[110\]\[2\] tms1x00.RAM\[111\]\[2\]
+ _0816_ _0977_ vssd1 vssd1 vccd1 vccd1 _1120_ sky130_fd_sc_hd__mux4_1
XFILLER_4_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2482__B2 _0818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4806__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4956__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2374__D_N net75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4147__B _1221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3670__A0 _1708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4750_ clknet_leaf_28_wb_clk_i _0364_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[55\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_4681_ clknet_leaf_4_wb_clk_i _0295_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[45\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_3701_ _1237_ _1310_ vssd1 vssd1 vccd1 vccd1 _1742_ sky130_fd_sc_hd__nor2_2
X_3632_ _1592_ tms1x00.RAM\[62\]\[3\] _1698_ vssd1 vssd1 vccd1 vccd1 _1702_ sky130_fd_sc_hd__mux2_1
X_3563_ _1590_ tms1x00.RAM\[51\]\[2\] _1659_ vssd1 vssd1 vccd1 vccd1 _1662_ sky130_fd_sc_hd__mux2_1
X_2514_ _0772_ _0858_ _0903_ _0906_ vssd1 vssd1 vccd1 vccd1 _0907_ sky130_fd_sc_hd__a31o_1
X_3494_ _1623_ vssd1 vssd1 vccd1 vccd1 _0314_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__2411__A _0039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3489__A0 _1588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2445_ _0797_ _0837_ vssd1 vssd1 vccd1 vccd1 _0838_ sky130_fd_sc_hd__or2_1
XFILLER_69_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2557__S _0948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4115_ tms1x00.CL _1974_ _1995_ _1976_ vssd1 vssd1 vccd1 vccd1 _1996_ sky130_fd_sc_hd__o31a_2
X_2376_ tms1x00.ins_in\[5\] tms1x00.ins_in\[4\] tms1x00.ins_in\[7\] tms1x00.ins_in\[6\]
+ vssd1 vssd1 vccd1 vccd1 _0769_ sky130_fd_sc_hd__and4b_1
XFILLER_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4046_ _1947_ vssd1 vssd1 vccd1 vccd1 _1948_ sky130_fd_sc_hd__inv_2
XFILLER_17_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3661__A0 _1708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4829__CLK clknet_leaf_20_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2464__A1 _0821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4979__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4073__A net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4948_ clknet_leaf_7_wb_clk_i _0558_ vssd1 vssd1 vccd1 vccd1 tms1x00.SR\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_33_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4879_ clknet_leaf_17_wb_clk_i _0493_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[93\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2321__A _0718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4141__A1 tms1x00.ins_in\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3152__A _0914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3652__A0 _1708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2455__A1 _0794_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3404__A0 _1492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2230_ net29 wbs_o_buff\[23\] _0679_ vssd1 vssd1 vccd1 vccd1 _0683_ sky130_fd_sc_hd__mux2_1
XFILLER_2_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2885__B _1261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3997__A net76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2446__A1 _0819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2541__S1 _0932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2406__A _0777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2994_ _1329_ vssd1 vssd1 vccd1 vccd1 _0108_ sky130_fd_sc_hd__clkbuf_1
X_4802_ clknet_leaf_22_wb_clk_i _0416_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[68\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4733_ clknet_leaf_27_wb_clk_i _0347_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[5\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3946__A1 _1327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4664_ clknet_leaf_28_wb_clk_i _0285_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[40\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_4595_ clknet_leaf_9_wb_clk_i _0216_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[126\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_3615_ _1692_ vssd1 vssd1 vccd1 vccd1 _0366_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4501__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4371__A1 _1330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3546_ _1652_ vssd1 vssd1 vccd1 vccd1 _0337_ sky130_fd_sc_hd__clkbuf_1
X_3477_ _1403_ _1525_ vssd1 vssd1 vccd1 vccd1 _1614_ sky130_fd_sc_hd__nor2_2
X_2428_ _0039_ vssd1 vssd1 vccd1 vccd1 _0821_ sky130_fd_sc_hd__clkbuf_4
X_2359_ tms1x00.Y\[3\] vssd1 vssd1 vccd1 vccd1 _0754_ sky130_fd_sc_hd__inv_2
XFILLER_57_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4651__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2780__S1 _0927_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4029_ _0754_ _0763_ _1935_ net84 vssd1 vssd1 vccd1 vccd1 _1936_ sky130_fd_sc_hd__a31o_1
XFILLER_71_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5007__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3937__A1 _1327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2599__S1 _0791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input34_A ram_val[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2771__S1 _0977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3928__A1 _1775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4524__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2600__B2 _0948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3057__A _1258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3400_ _1488_ tms1x00.RAM\[33\]\[1\] _1566_ vssd1 vssd1 vccd1 vccd1 _1568_ sky130_fd_sc_hd__mux2_1
X_4380_ _2173_ vssd1 vssd1 vccd1 vccd1 _0650_ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4674__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3331_ _1529_ vssd1 vssd1 vccd1 vccd1 _0245_ sky130_fd_sc_hd__clkbuf_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3262_ _1489_ vssd1 vssd1 vccd1 vccd1 _0216_ sky130_fd_sc_hd__clkbuf_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3504__B _1345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5001_ clknet_leaf_0_wb_clk_i _0611_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[21\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_2213_ net20 wbs_o_buff\[15\] _0668_ vssd1 vssd1 vccd1 vccd1 _0674_ sky130_fd_sc_hd__mux2_1
X_3193_ _1448_ vssd1 vssd1 vccd1 vccd1 _0188_ sky130_fd_sc_hd__clkbuf_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4041__B1 net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2977_ _0914_ _1317_ vssd1 vssd1 vccd1 vccd1 _1318_ sky130_fd_sc_hd__nor2_2
X_4716_ clknet_leaf_3_wb_clk_i _0330_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[46\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_4647_ clknet_leaf_6_wb_clk_i _0268_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[35\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_4578_ clknet_leaf_2_wb_clk_i _0199_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[118\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3529_ _1592_ tms1x00.RAM\[46\]\[3\] _1639_ vssd1 vssd1 vccd1 vccd1 _1643_ sky130_fd_sc_hd__mux2_1
XFILLER_39_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_27_wb_clk_i clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__4547__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2830__A1 _0040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4697__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2649__A1 _0940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2900_ _1130_ tms1x00.RAM\[79\]\[2\] _1268_ vssd1 vssd1 vccd1 vccd1 _1271_ sky130_fd_sc_hd__mux2_1
XFILLER_44_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3880_ _1258_ _1303_ vssd1 vssd1 vccd1 vccd1 _1845_ sky130_fd_sc_hd__nor2_2
X_2831_ _0835_ _1155_ _1175_ _1199_ _1220_ vssd1 vssd1 vccd1 vccd1 _1221_ sky130_fd_sc_hd__o32a_2
XFILLER_31_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2762_ _1149_ _1150_ _1151_ _0786_ _0828_ vssd1 vssd1 vccd1 vccd1 _1152_ sky130_fd_sc_hd__a221o_1
X_4501_ clknet_leaf_16_wb_clk_i _0122_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[98\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2376__A_N tms1x00.ins_in\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2714__B_N _0945_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4432_ clknet_leaf_14_wb_clk_i _0053_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[109\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2680__S0 _0808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2693_ _0922_ _1081_ _1083_ _0944_ vssd1 vssd1 vccd1 vccd1 _1084_ sky130_fd_sc_hd__o211a_1
X_4363_ _2164_ vssd1 vssd1 vccd1 vccd1 _0642_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__2888__A1 _1243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4294_ _1249_ _1345_ vssd1 vssd1 vccd1 vccd1 _2126_ sky130_fd_sc_hd__or2_2
X_3314_ _1250_ _1403_ vssd1 vssd1 vccd1 vccd1 _1519_ sky130_fd_sc_hd__nor2_2
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3245_ tms1x00.RAM\[116\]\[3\] _1463_ _1475_ vssd1 vssd1 vccd1 vccd1 _1479_ sky130_fd_sc_hd__mux2_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4049__C _0763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3176_ tms1x00.RAM\[123\]\[2\] _1331_ _1436_ vssd1 vssd1 vccd1 vccd1 _1439_ sky130_fd_sc_hd__mux2_1
XFILLER_27_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4081__A _0760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2882__C_N tms1x00.ram_addr_buff\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4308__A1 _1330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput70 net70 vssd1 vssd1 vccd1 vccd1 io_out[11] sky130_fd_sc_hd__buf_2
Xoutput92 net92 vssd1 vssd1 vccd1 vccd1 io_out[33] sky130_fd_sc_hd__buf_2
Xoutput81 net81 vssd1 vssd1 vccd1 vccd1 io_out[22] sky130_fd_sc_hd__buf_2
XFILLER_68_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3030_ _1353_ vssd1 vssd1 vccd1 vccd1 _0120_ sky130_fd_sc_hd__clkbuf_1
XFILLER_49_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4712__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4981_ clknet_leaf_8_wb_clk_i _0591_ vssd1 vssd1 vccd1 vccd1 tms1x00.A\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_17_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4862__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3932_ tms1x00.RAM\[91\]\[3\] _1779_ _1870_ vssd1 vssd1 vccd1 vccd1 _1874_ sky130_fd_sc_hd__mux2_1
XFILLER_32_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3863_ tms1x00.RAM\[86\]\[0\] _1772_ _1835_ vssd1 vssd1 vccd1 vccd1 _1836_ sky130_fd_sc_hd__mux2_1
X_2814_ tms1x00.RAM\[44\]\[3\] tms1x00.RAM\[45\]\[3\] tms1x00.RAM\[46\]\[3\] tms1x00.RAM\[47\]\[3\]
+ _0923_ _0791_ vssd1 vssd1 vccd1 vccd1 _1204_ sky130_fd_sc_hd__mux4_2
XFILLER_20_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3229__B _1430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3794_ _1795_ vssd1 vssd1 vccd1 vccd1 _0442_ sky130_fd_sc_hd__clkbuf_1
X_2745_ _0922_ _1132_ _1134_ _0776_ vssd1 vssd1 vccd1 vccd1 _1135_ sky130_fd_sc_hd__o211a_1
XANTENNA__3944__S _1880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2676_ tms1x00.RAM\[6\]\[2\] tms1x00.RAM\[7\]\[2\] _0815_ vssd1 vssd1 vccd1 vccd1
+ _1067_ sky130_fd_sc_hd__mux2_1
X_4415_ clknet_leaf_27_wb_clk_i _0013_ vssd1 vssd1 vccd1 vccd1 wbs_o_buff\[19\] sky130_fd_sc_hd__dfxtp_1
X_4346_ _1247_ tms1x00.RAM\[1\]\[3\] _2151_ vssd1 vssd1 vccd1 vccd1 _2155_ sky130_fd_sc_hd__mux2_1
XFILLER_59_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4277_ _1816_ tms1x00.RAM\[29\]\[0\] _2116_ vssd1 vssd1 vccd1 vccd1 _2117_ sky130_fd_sc_hd__mux2_1
XTAP_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3228_ _1469_ vssd1 vssd1 vccd1 vccd1 _0202_ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4076__A net73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3159_ tms1x00.RAM\[105\]\[3\] _1334_ _1425_ vssd1 vssd1 vccd1 vccd1 _1429_ sky130_fd_sc_hd__mux2_1
XFILLER_27_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4735__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4885__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output103_A net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3201__A1 _1328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2530_ _0921_ vssd1 vssd1 vccd1 vccd1 _0922_ sky130_fd_sc_hd__clkbuf_4
XFILLER_10_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2461_ tms1x00.RAM\[112\]\[0\] tms1x00.RAM\[113\]\[0\] tms1x00.RAM\[114\]\[0\] tms1x00.RAM\[115\]\[0\]
+ _0815_ _0812_ vssd1 vssd1 vccd1 vccd1 _0854_ sky130_fd_sc_hd__mux4_2
XFILLER_5_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4200_ tms1x00.P\[1\] tms1x00.N\[1\] vssd1 vssd1 vccd1 vccd1 _2066_ sky130_fd_sc_hd__nand2_1
XFILLER_68_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2392_ _0036_ vssd1 vssd1 vccd1 vccd1 _0785_ sky130_fd_sc_hd__inv_2
XFILLER_68_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4131_ _0858_ _0903_ vssd1 vssd1 vccd1 vccd1 _2008_ sky130_fd_sc_hd__nand2_1
XFILLER_68_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4062_ _0761_ _1957_ vssd1 vssd1 vccd1 vccd1 _1960_ sky130_fd_sc_hd__and2_1
X_3013_ _1342_ vssd1 vssd1 vccd1 vccd1 _0114_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__2409__A _0038_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4964_ clknet_leaf_7_wb_clk_i _0574_ vssd1 vssd1 vccd1 vccd1 tms1x00.PC\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5040__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3915_ _1864_ vssd1 vssd1 vccd1 vccd1 _0494_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4608__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4895_ clknet_leaf_0_wb_clk_i _0509_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[23\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3991__A2 _0724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3846_ _1826_ vssd1 vssd1 vccd1 vccd1 _0463_ sky130_fd_sc_hd__clkbuf_1
X_3777_ _1258_ _1345_ vssd1 vssd1 vccd1 vccd1 _1786_ sky130_fd_sc_hd__or2_2
X_2728_ _0921_ _1118_ vssd1 vssd1 vccd1 vccd1 _1119_ sky130_fd_sc_hd__or2_1
XANTENNA__4758__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2951__A0 _1225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2659_ _0798_ _1049_ vssd1 vssd1 vccd1 vccd1 _1050_ sky130_fd_sc_hd__or2_1
XANTENNA__2703__B1 _0794_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4329_ _2145_ vssd1 vssd1 vccd1 vccd1 _0627_ sky130_fd_sc_hd__clkbuf_1
XFILLER_47_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3982__A2 _0724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2942__A0 _1225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input64_A wbs_dat_i[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3498__A1 _1574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3422__A1 _1574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3700_ _1741_ vssd1 vssd1 vccd1 vccd1 _0402_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4900__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4680_ clknet_leaf_1_wb_clk_i _0294_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[38\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_3631_ _1701_ vssd1 vssd1 vccd1 vccd1 _0373_ sky130_fd_sc_hd__clkbuf_1
X_3562_ _1661_ vssd1 vssd1 vccd1 vccd1 _0344_ sky130_fd_sc_hd__clkbuf_1
X_2513_ tms1x00.ins_in\[2\] _0905_ vssd1 vssd1 vccd1 vccd1 _0906_ sky130_fd_sc_hd__nor2_1
X_3493_ _1592_ tms1x00.RAM\[50\]\[3\] _1619_ vssd1 vssd1 vccd1 vccd1 _1623_ sky130_fd_sc_hd__mux2_1
X_2444_ tms1x00.RAM\[104\]\[0\] tms1x00.RAM\[105\]\[0\] tms1x00.RAM\[106\]\[0\] tms1x00.RAM\[107\]\[0\]
+ _0777_ _0779_ vssd1 vssd1 vccd1 vccd1 _0837_ sky130_fd_sc_hd__mux4_1
XFILLER_68_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4150__A2 _2007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2375_ tms1x00.ins_in\[2\] vssd1 vssd1 vccd1 vccd1 _0768_ sky130_fd_sc_hd__inv_2
XFILLER_69_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4114_ tms1x00.status _0747_ vssd1 vssd1 vccd1 vccd1 _1995_ sky130_fd_sc_hd__nand2_4
XFILLER_69_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4045_ tms1x00.Y\[3\] tms1x00.Y\[2\] _0740_ vssd1 vssd1 vccd1 vccd1 _1947_ sky130_fd_sc_hd__and3_1
XFILLER_56_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4947_ clknet_leaf_7_wb_clk_i _0557_ vssd1 vssd1 vccd1 vccd1 tms1x00.SR\[4\] sky130_fd_sc_hd__dfxtp_1
X_4878_ clknet_leaf_17_wb_clk_i _0492_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[93\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4580__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3829_ tms1x00.RAM\[84\]\[3\] _1779_ _1811_ vssd1 vssd1 vccd1 vccd1 _1815_ sky130_fd_sc_hd__mux2_1
XFILLER_3_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2321__B _0724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2748__S _0789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3152__B _1261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3101__A0 _1368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2483__S _0823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2478__B_N _0789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3343__A _1249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4453__CLK clknet_leaf_20_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3997__B net75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4801_ clknet_leaf_24_wb_clk_i _0415_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[68\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2993_ tms1x00.RAM\[101\]\[1\] _1328_ _1325_ vssd1 vssd1 vccd1 vccd1 _1329_ sky130_fd_sc_hd__mux2_1
XFILLER_22_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4732_ clknet_leaf_3_wb_clk_i _0346_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[51\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4663_ clknet_leaf_27_wb_clk_i _0284_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[40\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_3614_ tms1x00.RAM\[55\]\[3\] _1676_ _1688_ vssd1 vssd1 vccd1 vccd1 _1692_ sky130_fd_sc_hd__mux2_1
XANTENNA__2906__A0 _0912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4594_ clknet_leaf_13_wb_clk_i _0215_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[126\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3952__S _0726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3545_ tms1x00.RAM\[53\]\[2\] _1576_ _1649_ vssd1 vssd1 vccd1 vccd1 _1652_ sky130_fd_sc_hd__mux2_1
X_3476_ _1613_ vssd1 vssd1 vccd1 vccd1 _0306_ sky130_fd_sc_hd__clkbuf_1
X_2427_ _0811_ _0814_ _0817_ _0818_ _0819_ vssd1 vssd1 vccd1 vccd1 _0820_ sky130_fd_sc_hd__a221o_1
X_2358_ _0752_ vssd1 vssd1 vccd1 vccd1 _0753_ sky130_fd_sc_hd__buf_2
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2289_ net92 _0697_ _0704_ wbs_o_buff\[23\] vssd1 vssd1 vccd1 vccd1 _0018_ sky130_fd_sc_hd__a22o_1
XFILLER_71_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4028_ _0739_ _1921_ vssd1 vssd1 vccd1 vccd1 _1935_ sky130_fd_sc_hd__nor2_1
XFILLER_71_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2316__B net75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3398__A0 _1485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3428__A _0911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2332__A _0732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2373__A1 chip_sel_override vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4476__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input27_A ram_val[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3389__A0 _1485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3057__B _1267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output95_A net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3330_ _1490_ tms1x00.RAM\[32\]\[2\] _1526_ vssd1 vssd1 vccd1 vccd1 _1529_ sky130_fd_sc_hd__mux2_1
XANTENNA__3561__A0 _1588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3261_ _1488_ tms1x00.RAM\[126\]\[1\] _1486_ vssd1 vssd1 vccd1 vccd1 _1489_ sky130_fd_sc_hd__mux2_1
X_5000_ clknet_leaf_0_wb_clk_i _0610_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[21\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_3_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4969__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2212_ _0673_ vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__clkbuf_1
X_3192_ tms1x00.RAM\[121\]\[1\] _1328_ _1446_ vssd1 vssd1 vccd1 vccd1 _1448_ sky130_fd_sc_hd__mux2_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2417__A _0807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4041__A1 _0732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2976_ _1316_ vssd1 vssd1 vccd1 vccd1 _1317_ sky130_fd_sc_hd__buf_4
X_4715_ clknet_leaf_5_wb_clk_i _0329_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[46\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_4646_ clknet_leaf_5_wb_clk_i _0267_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[35\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_4577_ clknet_leaf_2_wb_clk_i _0198_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[11\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_3528_ _1642_ vssd1 vssd1 vccd1 vccd1 _0329_ sky130_fd_sc_hd__clkbuf_1
XFILLER_77_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4079__A _0760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3459_ _1409_ _1524_ vssd1 vssd1 vccd1 vccd1 _1604_ sky130_fd_sc_hd__or2_2
XFILLER_58_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2761__S _0826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2594__A1 _0985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4099__A1 tms1x00.PC\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2649__A2 _1037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2806__C1 _0794_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2282__B1 _0703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2830_ _0040_ _1208_ _1219_ _0041_ vssd1 vssd1 vccd1 vccd1 _1220_ sky130_fd_sc_hd__a31o_1
XFILLER_32_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4023__A1 net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2761_ tms1x00.RAM\[76\]\[3\] tms1x00.RAM\[77\]\[3\] _0826_ vssd1 vssd1 vccd1 vccd1
+ _1151_ sky130_fd_sc_hd__mux2_1
XFILLER_31_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4641__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3782__A0 _1708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4500_ clknet_leaf_16_wb_clk_i _0121_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[98\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_2692_ _0953_ _1082_ vssd1 vssd1 vccd1 vccd1 _1083_ sky130_fd_sc_hd__or2_1
X_4431_ clknet_leaf_14_wb_clk_i _0052_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[109\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2680__S1 _0831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4362_ _1245_ tms1x00.RAM\[14\]\[2\] _2161_ vssd1 vssd1 vccd1 vccd1 _2164_ sky130_fd_sc_hd__mux2_1
XANTENNA__4791__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3313_ _1518_ vssd1 vssd1 vccd1 vccd1 _0238_ sky130_fd_sc_hd__clkbuf_1
X_4293_ _2125_ vssd1 vssd1 vccd1 vccd1 _0611_ sky130_fd_sc_hd__clkbuf_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3244_ _1478_ vssd1 vssd1 vccd1 vccd1 _0209_ sky130_fd_sc_hd__clkbuf_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3531__A _1284_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3175_ _1438_ vssd1 vssd1 vccd1 vccd1 _0180_ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2959_ _1306_ vssd1 vssd1 vccd1 vccd1 _0096_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__2576__A1 _0940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4629_ clknet_leaf_10_wb_clk_i _0250_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[31\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3525__A0 _1588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3441__A _1317_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4664__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4005__A1 net78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2567__A1 _0944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3516__A0 _1588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3616__A _1267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput93 net93 vssd1 vssd1 vccd1 vccd1 io_out[36] sky130_fd_sc_hd__buf_2
Xoutput82 net82 vssd1 vssd1 vccd1 vccd1 io_out[23] sky130_fd_sc_hd__buf_2
Xoutput71 net71 vssd1 vssd1 vccd1 vccd1 io_out[12] sky130_fd_sc_hd__buf_2
XFILLER_1_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4980_ clknet_leaf_8_wb_clk_i _0590_ vssd1 vssd1 vccd1 vccd1 tms1x00.A\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_23_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3931_ _1873_ vssd1 vssd1 vccd1 vccd1 _0501_ sky130_fd_sc_hd__clkbuf_1
X_3862_ _1258_ _1317_ vssd1 vssd1 vccd1 vccd1 _1835_ sky130_fd_sc_hd__nor2_2
X_2813_ _0921_ _1202_ vssd1 vssd1 vccd1 vccd1 _1203_ sky130_fd_sc_hd__or2_1
XFILLER_32_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3793_ tms1x00.RAM\[7\]\[3\] _1779_ _1791_ vssd1 vssd1 vccd1 vccd1 _1795_ sky130_fd_sc_hd__mux2_1
X_2744_ _0953_ _1133_ vssd1 vssd1 vccd1 vccd1 _1134_ sky130_fd_sc_hd__or2_1
XFILLER_9_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2675_ _1062_ _1064_ _1065_ _0948_ _0942_ vssd1 vssd1 vccd1 vccd1 _1066_ sky130_fd_sc_hd__o221a_1
XANTENNA__3507__A0 _1588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4414_ clknet_leaf_26_wb_clk_i _0012_ vssd1 vssd1 vccd1 vccd1 wbs_o_buff\[18\] sky130_fd_sc_hd__dfxtp_1
X_4345_ _2154_ vssd1 vssd1 vccd1 vccd1 _0634_ sky130_fd_sc_hd__clkbuf_1
X_4276_ _0917_ _1249_ vssd1 vssd1 vccd1 vccd1 _2116_ sky130_fd_sc_hd__or2_2
XTAP_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4357__A _1343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3227_ tms1x00.RAM\[118\]\[3\] _1463_ _1465_ vssd1 vssd1 vccd1 vccd1 _1469_ sky130_fd_sc_hd__mux2_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3158_ _1428_ vssd1 vssd1 vccd1 vccd1 _0173_ sky130_fd_sc_hd__clkbuf_1
XFILLER_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4687__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3089_ _1388_ vssd1 vssd1 vccd1 vccd1 _0144_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__2246__A0 net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2308__C valid vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2549__B2 _0787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_5_wb_clk_i_A clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_2_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3171__A _1286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4267__A _1250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5098__A net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2515__A tms1x00.ins_in\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3985__A0 tms1x00.ins_in\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_11_wb_clk_i clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_13_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2460_ _0849_ _0851_ _0852_ _0786_ _0828_ vssd1 vssd1 vccd1 vccd1 _0853_ sky130_fd_sc_hd__a221o_1
XFILLER_5_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2960__A1 _1245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4130_ _0701_ _2006_ vssd1 vssd1 vccd1 vccd1 _2007_ sky130_fd_sc_hd__nor2_2
X_2391_ _0781_ _0782_ _0783_ vssd1 vssd1 vccd1 vccd1 _0784_ sky130_fd_sc_hd__mux2_1
XFILLER_68_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4177__A tms1x00.PC\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4061_ _0742_ tms1x00.A\[0\] vssd1 vssd1 vccd1 vccd1 _1959_ sky130_fd_sc_hd__and2b_1
XFILLER_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3012_ tms1x00.RAM\[100\]\[3\] _1334_ _1338_ vssd1 vssd1 vccd1 vccd1 _1342_ sky130_fd_sc_hd__mux2_1
XANTENNA__2571__S0 _0945_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4963_ clknet_leaf_8_wb_clk_i _0573_ vssd1 vssd1 vccd1 vccd1 tms1x00.PC\[2\] sky130_fd_sc_hd__dfxtp_2
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2228__A0 net28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3914_ _1823_ tms1x00.RAM\[93\]\[3\] _1860_ vssd1 vssd1 vccd1 vccd1 _1864_ sky130_fd_sc_hd__mux2_1
XFILLER_60_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4894_ clknet_leaf_1_wb_clk_i _0508_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[23\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_3845_ _1816_ tms1x00.RAM\[82\]\[0\] _1825_ vssd1 vssd1 vccd1 vccd1 _1826_ sky130_fd_sc_hd__mux2_1
XFILLER_20_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3776_ _1785_ vssd1 vssd1 vccd1 vccd1 _0434_ sky130_fd_sc_hd__clkbuf_1
X_2727_ tms1x00.RAM\[96\]\[2\] tms1x00.RAM\[97\]\[2\] tms1x00.RAM\[98\]\[2\] tms1x00.RAM\[99\]\[2\]
+ _0873_ _0822_ vssd1 vssd1 vccd1 vccd1 _1118_ sky130_fd_sc_hd__mux4_2
XANTENNA__3256__A _0911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2658_ tms1x00.RAM\[48\]\[2\] tms1x00.RAM\[49\]\[2\] tms1x00.RAM\[50\]\[2\] tms1x00.RAM\[51\]\[2\]
+ _0799_ _0800_ vssd1 vssd1 vccd1 vccd1 _1049_ sky130_fd_sc_hd__mux4_2
XFILLER_59_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2589_ _0948_ _0974_ _0980_ _0776_ vssd1 vssd1 vccd1 vccd1 _0981_ sky130_fd_sc_hd__o211a_1
XANTENNA__2703__A1 _0786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4328_ _1823_ tms1x00.RAM\[127\]\[3\] _2141_ vssd1 vssd1 vccd1 vccd1 _2145_ sky130_fd_sc_hd__mux2_1
XANTENNA_input1_A io_in[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4087__A _0718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4259_ tms1x00.RAM\[39\]\[0\] _1323_ _2106_ vssd1 vssd1 vccd1 vccd1 _2107_ sky130_fd_sc_hd__mux2_1
XFILLER_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4852__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input57_A wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2458__B1 _0850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2630__B1 _0780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3630_ _1590_ tms1x00.RAM\[62\]\[2\] _1698_ vssd1 vssd1 vccd1 vccd1 _1701_ sky130_fd_sc_hd__mux2_1
X_3561_ _1588_ tms1x00.RAM\[51\]\[1\] _1659_ vssd1 vssd1 vccd1 vccd1 _1661_ sky130_fd_sc_hd__mux2_1
XANTENNA__4383__A0 tms1x00.PA\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3076__A _1251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2512_ tms1x00.ins_in\[3\] _0738_ _0746_ _0904_ vssd1 vssd1 vccd1 vccd1 _0905_ sky130_fd_sc_hd__or4_1
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2933__A1 _1247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3492_ _1622_ vssd1 vssd1 vccd1 vccd1 _0313_ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2443_ tms1x00.RAM\[108\]\[0\] tms1x00.RAM\[109\]\[0\] tms1x00.RAM\[110\]\[0\] tms1x00.RAM\[111\]\[0\]
+ _0799_ _0800_ vssd1 vssd1 vccd1 vccd1 _0836_ sky130_fd_sc_hd__mux4_1
XANTENNA__3804__A _0917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2374_ net76 net74 tms1x00.ins_in\[1\] net75 vssd1 vssd1 vccd1 vccd1 _0767_ sky130_fd_sc_hd__or4b_1
XANTENNA__2697__B1 _0996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4113_ _1994_ vssd1 vssd1 vccd1 vccd1 _0562_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4044_ _1946_ vssd1 vssd1 vccd1 vccd1 _0541_ sky130_fd_sc_hd__clkbuf_1
XFILLER_37_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2544__S0 _0924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4071__C1 _1966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4946_ clknet_leaf_7_wb_clk_i _0556_ vssd1 vssd1 vccd1 vccd1 tms1x00.SR\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4725__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4877_ clknet_leaf_18_wb_clk_i _0491_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[93\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_3828_ _1814_ vssd1 vssd1 vccd1 vccd1 _0457_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4875__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3759_ _1034_ vssd1 vssd1 vccd1 vccd1 _1775_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2512__B _0738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5030__CLK clknet_leaf_20_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3343__B _1396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4748__CLK clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4800_ clknet_leaf_22_wb_clk_i _0414_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[6\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2992_ _1327_ vssd1 vssd1 vccd1 vccd1 _1328_ sky130_fd_sc_hd__buf_2
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4731_ clknet_leaf_5_wb_clk_i _0345_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[51\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4898__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4662_ clknet_leaf_32_wb_clk_i _0283_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[40\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3159__A1 _1334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3613_ _1691_ vssd1 vssd1 vccd1 vccd1 _0365_ sky130_fd_sc_hd__clkbuf_1
X_4593_ clknet_leaf_15_wb_clk_i _0214_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[115\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_3544_ _1651_ vssd1 vssd1 vccd1 vccd1 _0336_ sky130_fd_sc_hd__clkbuf_1
X_3475_ tms1x00.RAM\[43\]\[3\] _1578_ _1609_ vssd1 vssd1 vccd1 vccd1 _1613_ sky130_fd_sc_hd__mux2_1
XFILLER_69_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2426_ _0793_ vssd1 vssd1 vccd1 vccd1 _0819_ sky130_fd_sc_hd__clkbuf_4
X_2357_ tms1x00.ins_in\[1\] _0742_ _0744_ _0751_ vssd1 vssd1 vccd1 vccd1 _0752_ sky130_fd_sc_hd__or4_4
XFILLER_29_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2288_ net91 _0697_ _0704_ wbs_o_buff\[22\] vssd1 vssd1 vccd1 vccd1 _0017_ sky130_fd_sc_hd__a22o_1
XANTENNA__3095__A0 _1361_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4027_ net83 _1933_ _1934_ _1931_ vssd1 vssd1 vccd1 vccd1 _0536_ sky130_fd_sc_hd__o211a_1
XFILLER_56_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2842__A0 _0912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4929_ clknet_leaf_9_wb_clk_i _0539_ vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__dfxtp_2
XFILLER_60_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3570__A1 _1574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2756__S0 _0830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3086__A0 _1361_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2833__B1 _1221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output88_A net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4420__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3260_ _1034_ vssd1 vssd1 vccd1 vccd1 _1488_ sky130_fd_sc_hd__buf_2
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2211_ net19 wbs_o_buff\[14\] _0668_ vssd1 vssd1 vccd1 vccd1 _0673_ sky130_fd_sc_hd__mux2_1
X_3191_ _1447_ vssd1 vssd1 vccd1 vccd1 _0187_ sky130_fd_sc_hd__clkbuf_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4570__CLK clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3077__A0 _1361_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4041__A2 _0763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4714_ clknet_leaf_4_wb_clk_i _0328_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[46\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_2975_ _1238_ tms1x00.ram_addr_buff\[0\] _0728_ vssd1 vssd1 vccd1 vccd1 _1316_ sky130_fd_sc_hd__or3b_1
XANTENNA__2588__C1 _0819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4645_ clknet_leaf_1_wb_clk_i _0266_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[36\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_4576_ clknet_leaf_1_wb_clk_i _0197_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[11\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_3527_ _1590_ tms1x00.RAM\[46\]\[2\] _1639_ vssd1 vssd1 vccd1 vccd1 _1642_ sky130_fd_sc_hd__mux2_1
XFILLER_2_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3552__A1 _1574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4913__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3458_ _1603_ vssd1 vssd1 vccd1 vccd1 _0298_ sky130_fd_sc_hd__clkbuf_1
XFILLER_76_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3389_ _1485_ tms1x00.RAM\[34\]\[0\] _1561_ vssd1 vssd1 vccd1 vccd1 _1562_ sky130_fd_sc_hd__mux2_1
X_2409_ _0038_ vssd1 vssd1 vccd1 vccd1 _0802_ sky130_fd_sc_hd__clkbuf_4
XFILLER_69_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3068__A0 _1361_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4443__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3791__A1 _1777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3543__A1 _1574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2751__C1 _0942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2729__S0 _0816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2282__A1 net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2760_ _0778_ tms1x00.RAM\[78\]\[3\] _0812_ vssd1 vssd1 vccd1 vccd1 _1150_ sky130_fd_sc_hd__o21a_1
XFILLER_8_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2691_ tms1x00.RAM\[84\]\[2\] tms1x00.RAM\[85\]\[2\] tms1x00.RAM\[86\]\[2\] tms1x00.RAM\[87\]\[2\]
+ _0873_ _0977_ vssd1 vssd1 vccd1 vccd1 _1082_ sky130_fd_sc_hd__mux4_1
XFILLER_8_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4430_ clknet_leaf_14_wb_clk_i _0051_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[109\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4936__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2399__S _0788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3534__A1 _1574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4361_ _2163_ vssd1 vssd1 vccd1 vccd1 _0641_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3312_ tms1x00.RAM\[27\]\[3\] _1463_ _1514_ vssd1 vssd1 vccd1 vccd1 _1518_ sky130_fd_sc_hd__mux2_1
X_4292_ tms1x00.RAM\[21\]\[3\] _1333_ _2121_ vssd1 vssd1 vccd1 vccd1 _2125_ sky130_fd_sc_hd__mux2_1
XFILLER_4_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3243_ tms1x00.RAM\[116\]\[2\] _1461_ _1475_ vssd1 vssd1 vccd1 vccd1 _1478_ sky130_fd_sc_hd__mux2_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3531__B _1317_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3174_ tms1x00.RAM\[123\]\[1\] _1328_ _1436_ vssd1 vssd1 vccd1 vccd1 _1438_ sky130_fd_sc_hd__mux2_1
XFILLER_81_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2428__A _0039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4466__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2958_ tms1x00.RAM\[104\]\[1\] _1243_ _1304_ vssd1 vssd1 vccd1 vccd1 _1306_ sky130_fd_sc_hd__mux2_1
XFILLER_22_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3773__A1 _1777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4628_ clknet_leaf_8_wb_clk_i _0249_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[31\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_2889_ _1264_ vssd1 vssd1 vccd1 vccd1 _0068_ sky130_fd_sc_hd__clkbuf_1
X_4559_ clknet_leaf_35_wb_clk_i _0180_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[123\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_77_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3441__B _1525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4809__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2264__A1 net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4959__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3616__B _1283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput94 net94 vssd1 vssd1 vccd1 vccd1 io_out[37] sky130_fd_sc_hd__buf_2
Xoutput83 net83 vssd1 vssd1 vccd1 vccd1 io_out[24] sky130_fd_sc_hd__buf_2
Xoutput72 net72 vssd1 vssd1 vccd1 vccd1 io_out[13] sky130_fd_sc_hd__buf_2
XFILLER_68_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4229__C1 _0766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3930_ tms1x00.RAM\[91\]\[2\] _1777_ _1870_ vssd1 vssd1 vccd1 vccd1 _1873_ sky130_fd_sc_hd__mux2_1
XFILLER_32_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3861_ _1834_ vssd1 vssd1 vccd1 vccd1 _0470_ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2812_ tms1x00.RAM\[32\]\[3\] tms1x00.RAM\[33\]\[3\] tms1x00.RAM\[34\]\[3\] tms1x00.RAM\[35\]\[3\]
+ _0816_ _0927_ vssd1 vssd1 vccd1 vccd1 _1202_ sky130_fd_sc_hd__mux4_2
XFILLER_32_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3792_ _1794_ vssd1 vssd1 vccd1 vccd1 _0441_ sky130_fd_sc_hd__clkbuf_1
X_2743_ tms1x00.RAM\[84\]\[3\] tms1x00.RAM\[85\]\[3\] tms1x00.RAM\[86\]\[3\] tms1x00.RAM\[87\]\[3\]
+ _0840_ _0813_ vssd1 vssd1 vccd1 vccd1 _1133_ sky130_fd_sc_hd__mux4_1
X_2674_ tms1x00.RAM\[24\]\[2\] tms1x00.RAM\[25\]\[2\] tms1x00.RAM\[26\]\[2\] tms1x00.RAM\[27\]\[2\]
+ _0955_ _0956_ vssd1 vssd1 vccd1 vccd1 _1065_ sky130_fd_sc_hd__mux4_2
X_4413_ clknet_leaf_28_wb_clk_i _0011_ vssd1 vssd1 vccd1 vccd1 wbs_o_buff\[17\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__4180__A1 _0748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4344_ _1245_ tms1x00.RAM\[1\]\[2\] _2151_ vssd1 vssd1 vccd1 vccd1 _2154_ sky130_fd_sc_hd__mux2_1
X_4275_ _2115_ vssd1 vssd1 vccd1 vccd1 _0603_ sky130_fd_sc_hd__clkbuf_1
XTAP_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3226_ _1468_ vssd1 vssd1 vccd1 vccd1 _0201_ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4357__B _1396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3157_ tms1x00.RAM\[105\]\[2\] _1331_ _1425_ vssd1 vssd1 vccd1 vccd1 _1428_ sky130_fd_sc_hd__mux2_1
XFILLER_55_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3088_ _1364_ tms1x00.RAM\[112\]\[1\] _1386_ vssd1 vssd1 vccd1 vccd1 _1388_ sky130_fd_sc_hd__mux2_1
XFILLER_42_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2621__A _0798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4171__A1 net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2182__A0 net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4267__B _1317_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4631__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3171__B _1430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2515__B _0742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2531__A _0826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output70_A net70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2390_ _0037_ vssd1 vssd1 vccd1 vccd1 _0783_ sky130_fd_sc_hd__clkbuf_4
XFILLER_69_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4060_ _0761_ _1957_ vssd1 vssd1 vccd1 vccd1 _1958_ sky130_fd_sc_hd__nand2_1
XFILLER_37_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3011_ _1341_ vssd1 vssd1 vccd1 vccd1 _0113_ sky130_fd_sc_hd__clkbuf_1
XFILLER_64_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2571__S1 _0791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4962_ clknet_leaf_7_wb_clk_i _0572_ vssd1 vssd1 vccd1 vccd1 tms1x00.PC\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3913_ _1863_ vssd1 vssd1 vccd1 vccd1 _0493_ sky130_fd_sc_hd__clkbuf_1
X_4893_ clknet_leaf_0_wb_clk_i _0507_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[23\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_60_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3844_ _1257_ _1273_ vssd1 vssd1 vccd1 vccd1 _1825_ sky130_fd_sc_hd__or2_2
XFILLER_32_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3775_ tms1x00.RAM\[73\]\[3\] _1779_ _1781_ vssd1 vssd1 vccd1 vccd1 _1785_ sky130_fd_sc_hd__mux2_1
XANTENNA__4504__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2726_ _0953_ _1116_ vssd1 vssd1 vccd1 vccd1 _1117_ sky130_fd_sc_hd__or2_1
X_2657_ _1045_ _1046_ _1047_ _0818_ _0953_ vssd1 vssd1 vccd1 vccd1 _1048_ sky130_fd_sc_hd__a221o_1
XANTENNA__3971__S _0724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4654__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2588_ _0976_ _0978_ _0979_ _0818_ _0819_ vssd1 vssd1 vccd1 vccd1 _0980_ sky130_fd_sc_hd__a221o_1
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4327_ _2144_ vssd1 vssd1 vccd1 vccd1 _0626_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__2587__S _0923_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4258_ _1310_ _1525_ vssd1 vssd1 vccd1 vccd1 _2106_ sky130_fd_sc_hd__nor2_2
XFILLER_74_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3209_ tms1x00.RAM\[11\]\[0\] _1456_ _1457_ vssd1 vssd1 vccd1 vccd1 _1458_ sky130_fd_sc_hd__mux2_1
X_4189_ tms1x00.PC\[5\] _1908_ _0766_ vssd1 vssd1 vccd1 vccd1 _2057_ sky130_fd_sc_hd__o21a_1
XFILLER_55_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2458__A1 _0808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3958__A1 tms1x00.ram_addr_buff\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2630__A1 _0840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3560_ _1660_ vssd1 vssd1 vccd1 vccd1 _0343_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__2261__A _0699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3076__B _1375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2511_ _0747_ _0762_ _0748_ tms1x00.ins_in\[5\] vssd1 vssd1 vccd1 vccd1 _0904_ sky130_fd_sc_hd__or4b_1
XFILLER_6_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4677__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3491_ _1590_ tms1x00.RAM\[50\]\[2\] _1619_ vssd1 vssd1 vccd1 vccd1 _1622_ sky130_fd_sc_hd__mux2_1
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2442_ _0041_ vssd1 vssd1 vccd1 vccd1 _0835_ sky130_fd_sc_hd__inv_2
XANTENNA__3804__B _1236_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2373_ chip_sel_override _0714_ _0716_ net64 vssd1 vssd1 vccd1 vccd1 _0050_ sky130_fd_sc_hd__a22o_1
XANTENNA__2697__A1 _0787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4112_ net103 _1993_ vssd1 vssd1 vccd1 vccd1 _1994_ sky130_fd_sc_hd__or2_1
X_4043_ _0718_ _1944_ _1945_ vssd1 vssd1 vccd1 vccd1 _1946_ sky130_fd_sc_hd__and3_1
XFILLER_65_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2544__S1 _0928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4945_ clknet_leaf_7_wb_clk_i _0555_ vssd1 vssd1 vccd1 vccd1 tms1x00.SR\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_52_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4876_ clknet_leaf_17_wb_clk_i _0490_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[94\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3827_ tms1x00.RAM\[84\]\[2\] _1777_ _1811_ vssd1 vssd1 vccd1 vccd1 _1814_ sky130_fd_sc_hd__mux2_1
X_3758_ _1774_ vssd1 vssd1 vccd1 vccd1 _0427_ sky130_fd_sc_hd__clkbuf_1
X_2709_ tms1x00.RAM\[76\]\[2\] tms1x00.RAM\[77\]\[2\] _0788_ vssd1 vssd1 vccd1 vccd1
+ _1100_ sky130_fd_sc_hd__mux2_1
XFILLER_4_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3689_ _1735_ vssd1 vssd1 vccd1 vccd1 _0397_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2860__A1 _1243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2612__A1 _0928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3628__A0 _1588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2991_ _1033_ vssd1 vssd1 vccd1 vccd1 _1327_ sky130_fd_sc_hd__clkbuf_4
XFILLER_15_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4730_ clknet_leaf_3_wb_clk_i _0344_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[51\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3800__A0 _1708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4661_ clknet_leaf_27_wb_clk_i _0282_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[41\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_3612_ tms1x00.RAM\[55\]\[2\] _1674_ _1688_ vssd1 vssd1 vccd1 vccd1 _1691_ sky130_fd_sc_hd__mux2_1
X_4592_ clknet_leaf_15_wb_clk_i _0213_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[115\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_29_wb_clk_i_A clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_3543_ tms1x00.RAM\[53\]\[1\] _1574_ _1649_ vssd1 vssd1 vccd1 vccd1 _1651_ sky130_fd_sc_hd__mux2_1
X_3474_ _1612_ vssd1 vssd1 vccd1 vccd1 _0305_ sky130_fd_sc_hd__clkbuf_1
X_2425_ _0785_ vssd1 vssd1 vccd1 vccd1 _0818_ sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_2_2__f_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_0_wb_clk_i_A wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2356_ _0746_ _0750_ vssd1 vssd1 vccd1 vccd1 _0751_ sky130_fd_sc_hd__or2_1
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3619__A0 _1588_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2287_ net90 _0697_ _0704_ wbs_o_buff\[21\] vssd1 vssd1 vccd1 vccd1 _0016_ sky130_fd_sc_hd__a22o_1
X_4026_ _0732_ _0753_ _1932_ vssd1 vssd1 vccd1 vccd1 _1934_ sky130_fd_sc_hd__or3_1
XFILLER_37_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4928_ clknet_leaf_9_wb_clk_i _0538_ vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__dfxtp_2
XFILLER_12_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4859_ clknet_leaf_23_wb_clk_i _0473_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[86\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4992__CLK clknet_leaf_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3858__A0 _1821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2756__S1 _0831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4283__A0 _1823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2523__B tms1x00.ram_addr_buff\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3010__A1 _1331_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2444__S0 _0777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3635__A _0917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3849__A0 _1821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4715__CLK clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2210_ _0672_ vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__clkbuf_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3190_ tms1x00.RAM\[121\]\[0\] _1324_ _1446_ vssd1 vssd1 vccd1 vccd1 _1447_ sky130_fd_sc_hd__mux2_1
XANTENNA__2685__S _0823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3370__A _1337_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4865__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2974_ _1315_ vssd1 vssd1 vccd1 vccd1 _0102_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_6_wb_clk_i clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_4713_ clknet_leaf_4_wb_clk_i _0327_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[46\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4644_ clknet_leaf_1_wb_clk_i _0265_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[36\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_4575_ clknet_leaf_2_wb_clk_i _0196_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[11\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3001__A1 _1334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3526_ _1641_ vssd1 vssd1 vccd1 vccd1 _0328_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__2760__B1 _0812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3457_ _1592_ tms1x00.RAM\[45\]\[3\] _1599_ vssd1 vssd1 vccd1 vccd1 _1603_ sky130_fd_sc_hd__mux2_1
XFILLER_39_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3388_ _1273_ _1524_ vssd1 vssd1 vccd1 vccd1 _1561_ sky130_fd_sc_hd__or2_2
X_2408_ tms1x00.RAM\[88\]\[0\] tms1x00.RAM\[89\]\[0\] tms1x00.RAM\[90\]\[0\] tms1x00.RAM\[91\]\[0\]
+ _0799_ _0800_ vssd1 vssd1 vccd1 vccd1 _0801_ sky130_fd_sc_hd__mux4_1
XFILLER_58_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2339_ tms1x00.X\[1\] tms1x00.ram_addr_buff\[6\] _0726_ vssd1 vssd1 vccd1 vccd1 _0737_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__2595__S _0873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4009_ net79 _1919_ _1920_ _1901_ vssd1 vssd1 vccd1 vccd1 _0532_ sky130_fd_sc_hd__o211a_1
XFILLER_44_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4017__B1 net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5020__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2674__S0 _0955_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2343__B valid vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4738__CLK clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2729__S1 _0977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2503__B1 _0812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input32_A ram_val[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4888__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2806__B2 _0786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2534__A _0787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2690_ tms1x00.RAM\[80\]\[2\] tms1x00.RAM\[81\]\[2\] tms1x00.RAM\[82\]\[2\] tms1x00.RAM\[83\]\[2\]
+ _0931_ _0932_ vssd1 vssd1 vccd1 vccd1 _1081_ sky130_fd_sc_hd__mux4_2
X_4360_ _1243_ tms1x00.RAM\[14\]\[1\] _2161_ vssd1 vssd1 vccd1 vccd1 _2163_ sky130_fd_sc_hd__mux2_1
XFILLER_6_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3311_ _1517_ vssd1 vssd1 vccd1 vccd1 _0237_ sky130_fd_sc_hd__clkbuf_1
X_4291_ _2124_ vssd1 vssd1 vccd1 vccd1 _0610_ sky130_fd_sc_hd__clkbuf_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3242_ _1477_ vssd1 vssd1 vccd1 vccd1 _0208_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4196__A tms1x00.ins_in\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3173_ _1437_ vssd1 vssd1 vccd1 vccd1 _0179_ sky130_fd_sc_hd__clkbuf_1
XFILLER_66_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5043__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3974__S _0724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2957_ _1305_ vssd1 vssd1 vccd1 vccd1 _0095_ sky130_fd_sc_hd__clkbuf_1
X_2888_ tms1x00.RAM\[89\]\[1\] _1243_ _1262_ vssd1 vssd1 vccd1 vccd1 _1264_ sky130_fd_sc_hd__mux2_1
X_4627_ clknet_leaf_10_wb_clk_i _0248_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[31\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2408__S0 _0799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4558_ clknet_leaf_31_wb_clk_i _0179_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[123\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2733__B1 _0821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3509_ _1590_ tms1x00.RAM\[48\]\[2\] _1629_ vssd1 vssd1 vccd1 vccd1 _1632_ sky130_fd_sc_hd__mux2_1
X_4489_ clknet_leaf_29_wb_clk_i _0110_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[101\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_66_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2497__C1 _0775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2500__A3 tms1x00.RAM\[63\]\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2354__A _0747_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4410__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2647__S0 _0830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2724__B1 _0804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput84 net84 vssd1 vssd1 vccd1 vccd1 io_out[25] sky130_fd_sc_hd__buf_2
Xoutput73 net73 vssd1 vssd1 vccd1 vccd1 io_out[14] sky130_fd_sc_hd__buf_2
XFILLER_49_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput95 net95 vssd1 vssd1 vccd1 vccd1 oram_addr[0] sky130_fd_sc_hd__buf_2
XFILLER_0_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2488__C1 _0775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4903__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3860_ _1823_ tms1x00.RAM\[81\]\[3\] _1830_ vssd1 vssd1 vccd1 vccd1 _1834_ sky130_fd_sc_hd__mux2_1
XFILLER_31_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2811_ _0996_ _1200_ vssd1 vssd1 vccd1 vccd1 _1201_ sky130_fd_sc_hd__or2_1
X_3791_ tms1x00.RAM\[7\]\[2\] _1777_ _1791_ vssd1 vssd1 vccd1 vccd1 _1794_ sky130_fd_sc_hd__mux2_1
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2742_ tms1x00.RAM\[80\]\[3\] tms1x00.RAM\[81\]\[3\] tms1x00.RAM\[82\]\[3\] tms1x00.RAM\[83\]\[3\]
+ _0931_ _0932_ vssd1 vssd1 vccd1 vccd1 _1132_ sky130_fd_sc_hd__mux4_1
XFILLER_9_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2412__C1 _0804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2673_ _0818_ _1063_ _0953_ vssd1 vssd1 vccd1 vccd1 _1064_ sky130_fd_sc_hd__a21o_1
XANTENNA__2203__S _0668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4412_ clknet_leaf_26_wb_clk_i _0010_ vssd1 vssd1 vccd1 vccd1 wbs_o_buff\[16\] sky130_fd_sc_hd__dfxtp_1
X_4343_ _2153_ vssd1 vssd1 vccd1 vccd1 _0633_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__2810__S0 _0816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2715__B1 _0927_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4274_ tms1x00.RAM\[22\]\[3\] _1333_ _2111_ vssd1 vssd1 vccd1 vccd1 _2115_ sky130_fd_sc_hd__mux2_1
X_3225_ tms1x00.RAM\[118\]\[2\] _1461_ _1465_ vssd1 vssd1 vccd1 vccd1 _1468_ sky130_fd_sc_hd__mux2_1
XFILLER_67_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3969__S _0738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3156_ _1427_ vssd1 vssd1 vccd1 vccd1 _0172_ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3087_ _1387_ vssd1 vssd1 vccd1 vccd1 _0143_ sky130_fd_sc_hd__clkbuf_1
XFILLER_54_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4583__CLK clknet_leaf_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3989_ _0748_ _0724_ _1906_ _1901_ vssd1 vssd1 vccd1 vccd1 _0526_ sky130_fd_sc_hd__o211a_1
XFILLER_10_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2621__B _1012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4156__C1 _0701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2945__A0 _0912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4456__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_20_wb_clk_i clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2259__A _0697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3010_ tms1x00.RAM\[100\]\[2\] _1331_ _1338_ vssd1 vssd1 vccd1 vccd1 _1341_ sky130_fd_sc_hd__mux2_1
XFILLER_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4961_ clknet_leaf_7_wb_clk_i _0571_ vssd1 vssd1 vccd1 vccd1 tms1x00.PC\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_52_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3912_ _1821_ tms1x00.RAM\[93\]\[2\] _1860_ vssd1 vssd1 vccd1 vccd1 _1863_ sky130_fd_sc_hd__mux2_1
X_4892_ clknet_leaf_29_wb_clk_i _0506_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[90\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_3843_ _1824_ vssd1 vssd1 vccd1 vccd1 _0462_ sky130_fd_sc_hd__clkbuf_1
XFILLER_32_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2722__A _0783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2936__A0 _0912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3774_ _1784_ vssd1 vssd1 vccd1 vccd1 _0433_ sky130_fd_sc_hd__clkbuf_1
X_2725_ tms1x00.RAM\[100\]\[2\] tms1x00.RAM\[101\]\[2\] tms1x00.RAM\[102\]\[2\] tms1x00.RAM\[103\]\[2\]
+ _0873_ _0822_ vssd1 vssd1 vccd1 vccd1 _1116_ sky130_fd_sc_hd__mux4_1
X_2656_ tms1x00.RAM\[52\]\[2\] tms1x00.RAM\[53\]\[2\] _0923_ vssd1 vssd1 vccd1 vccd1
+ _1047_ sky130_fd_sc_hd__mux2_1
X_2587_ tms1x00.RAM\[116\]\[1\] tms1x00.RAM\[117\]\[1\] _0923_ vssd1 vssd1 vccd1 vccd1
+ _0979_ sky130_fd_sc_hd__mux2_1
X_4326_ _1821_ tms1x00.RAM\[127\]\[2\] _2141_ vssd1 vssd1 vccd1 vccd1 _2144_ sky130_fd_sc_hd__mux2_1
XFILLER_75_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4257_ _2105_ vssd1 vssd1 vccd1 vccd1 _0595_ sky130_fd_sc_hd__clkbuf_1
Xfanout148 net94 vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__buf_4
X_4188_ tms1x00.PC\[4\] _2048_ _2054_ _0760_ vssd1 vssd1 vccd1 vccd1 _2056_ sky130_fd_sc_hd__a31o_1
XFILLER_55_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4949__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3208_ _1286_ _1344_ vssd1 vssd1 vccd1 vccd1 _1457_ sky130_fd_sc_hd__nor2_2
XFILLER_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3139_ tms1x00.RAM\[107\]\[2\] _1331_ _1415_ vssd1 vssd1 vccd1 vccd1 _1418_ sky130_fd_sc_hd__mux2_1
XFILLER_27_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2624__C1 _0804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3728__A _1237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4294__A _1249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output101_A net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2615__C1 _0920_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3638__A _1034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2918__A0 K_override\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3490_ _1621_ vssd1 vssd1 vccd1 vccd1 _0312_ sky130_fd_sc_hd__clkbuf_1
X_2510_ _0773_ _0868_ _0882_ _0902_ _0041_ vssd1 vssd1 vccd1 vccd1 _0903_ sky130_fd_sc_hd__a311o_1
XANTENNA_clkbuf_leaf_19_wb_clk_i_A clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_2441_ _0806_ _0810_ _0820_ _0821_ _0833_ vssd1 vssd1 vccd1 vccd1 _0834_ sky130_fd_sc_hd__a311o_1
XFILLER_6_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2372_ _0733_ _0741_ _0753_ _0765_ _0766_ vssd1 vssd1 vccd1 vccd1 _0049_ sky130_fd_sc_hd__o311a_1
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3894__A1 _1777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4111_ tms1x00.PA\[3\] _1973_ _1987_ tms1x00.PB\[3\] vssd1 vssd1 vccd1 vccd1 _1993_
+ sky130_fd_sc_hd__a22o_1
XFILLER_68_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4042_ _0754_ _0752_ _1922_ vssd1 vssd1 vccd1 vccd1 _1945_ sky130_fd_sc_hd__or3b_1
XFILLER_65_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3312__S _1514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4944_ clknet_leaf_7_wb_clk_i _0554_ vssd1 vssd1 vccd1 vccd1 tms1x00.SR\[1\] sky130_fd_sc_hd__dfxtp_1
X_4875_ clknet_leaf_17_wb_clk_i _0489_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[94\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3826_ _1813_ vssd1 vssd1 vccd1 vccd1 _0456_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4621__CLK clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3757_ tms1x00.RAM\[74\]\[0\] _1772_ _1773_ vssd1 vssd1 vccd1 vccd1 _1774_ sky130_fd_sc_hd__mux2_1
X_2708_ _0830_ tms1x00.RAM\[78\]\[2\] _0850_ vssd1 vssd1 vccd1 vccd1 _1099_ sky130_fd_sc_hd__o21a_1
X_3688_ _1708_ tms1x00.RAM\[64\]\[2\] _1732_ vssd1 vssd1 vccd1 vccd1 _1735_ sky130_fd_sc_hd__mux2_1
X_2639_ _0747_ _0748_ vssd1 vssd1 vccd1 vccd1 _1031_ sky130_fd_sc_hd__and2b_1
XFILLER_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3885__A1 _1777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4309_ _2134_ vssd1 vssd1 vccd1 vccd1 _0618_ sky130_fd_sc_hd__clkbuf_1
XFILLER_75_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input62_A wbs_dat_i[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3876__A1 _1777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3628__A1 tms1x00.RAM\[62\]\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2990_ _1326_ vssd1 vssd1 vccd1 vccd1 _0107_ sky130_fd_sc_hd__clkbuf_1
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4644__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4660_ clknet_leaf_31_wb_clk_i _0281_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[41\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_3611_ _1690_ vssd1 vssd1 vccd1 vccd1 _0364_ sky130_fd_sc_hd__clkbuf_1
X_4591_ clknet_leaf_14_wb_clk_i _0212_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[115\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_3542_ _1650_ vssd1 vssd1 vccd1 vccd1 _0335_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4794__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3473_ tms1x00.RAM\[43\]\[2\] _1576_ _1609_ vssd1 vssd1 vccd1 vccd1 _1612_ sky130_fd_sc_hd__mux2_1
XFILLER_69_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2424_ tms1x00.RAM\[76\]\[0\] tms1x00.RAM\[77\]\[0\] _0816_ vssd1 vssd1 vccd1 vccd1
+ _0817_ sky130_fd_sc_hd__mux2_1
XANTENNA__2211__S _0668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3867__A1 _1777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2355_ tms1x00.ins_in\[4\] _0749_ vssd1 vssd1 vccd1 vccd1 _0750_ sky130_fd_sc_hd__or2_1
XFILLER_69_466 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3831__A _0911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3619__A1 tms1x00.RAM\[63\]\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2286_ net89 _0697_ _0704_ wbs_o_buff\[20\] vssd1 vssd1 vccd1 vccd1 _0015_ sky130_fd_sc_hd__a22o_1
X_4025_ _1932_ _0755_ _0764_ vssd1 vssd1 vccd1 vccd1 _1933_ sky130_fd_sc_hd__and3b_1
XANTENNA__2447__A _0815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4292__A1 _1333_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4927_ clknet_leaf_9_wb_clk_i _0537_ vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__dfxtp_2
XFILLER_52_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3278__A _1250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4858_ clknet_leaf_23_wb_clk_i _0472_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[86\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3809_ _1708_ tms1x00.RAM\[77\]\[2\] _1801_ vssd1 vssd1 vccd1 vccd1 _1804_ sky130_fd_sc_hd__mux2_1
X_4789_ clknet_leaf_24_wb_clk_i _0403_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[71\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2357__A tms1x00.ins_in\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4667__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2523__C tms1x00.ram_addr_buff\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3916__A _1257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2444__S1 _0779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3635__B _1283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2267__A net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3370__B _1525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2809__C1 _0773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4274__A1 _1333_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2973_ tms1x00.RAM\[103\]\[3\] _1247_ _1311_ vssd1 vssd1 vccd1 vccd1 _1315_ sky130_fd_sc_hd__mux2_1
X_4712_ clknet_leaf_5_wb_clk_i _0326_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[47\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2588__B2 _0818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4643_ clknet_leaf_1_wb_clk_i _0264_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[36\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_4574_ clknet_leaf_1_wb_clk_i _0195_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[11\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_3525_ _1588_ tms1x00.RAM\[46\]\[1\] _1639_ vssd1 vssd1 vccd1 vccd1 _1641_ sky130_fd_sc_hd__mux2_1
XANTENNA__2760__A1 _0778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3456_ _1602_ vssd1 vssd1 vccd1 vccd1 _0297_ sky130_fd_sc_hd__clkbuf_1
X_3387_ _1560_ vssd1 vssd1 vccd1 vccd1 _0270_ sky130_fd_sc_hd__clkbuf_1
X_2407_ _0779_ vssd1 vssd1 vccd1 vccd1 _0800_ sky130_fd_sc_hd__buf_6
XFILLER_69_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2338_ _0736_ vssd1 vssd1 vccd1 vccd1 _0047_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2269_ net75 _0698_ _0700_ wbs_o_buff\[6\] vssd1 vssd1 vccd1 vccd1 _0031_ sky130_fd_sc_hd__a22o_1
X_4008_ _0732_ _0730_ _0752_ _1918_ vssd1 vssd1 vccd1 vccd1 _1920_ sky130_fd_sc_hd__or4b_1
XANTENNA__4265__A1 _1333_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2276__B1 _0703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2905__A _1250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2674__S1 _0956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2200__A0 net45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2751__B2 _0922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2503__A1 _0778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2707__B_N _0830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input25_A ram_val[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4256__A1 _1333_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2550__A _0802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output93_A net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3310_ tms1x00.RAM\[27\]\[2\] _1461_ _1514_ vssd1 vssd1 vccd1 vccd1 _1517_ sky130_fd_sc_hd__mux2_1
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4290_ tms1x00.RAM\[21\]\[2\] _1330_ _2121_ vssd1 vssd1 vccd1 vccd1 _2124_ sky130_fd_sc_hd__mux2_1
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2696__S _0975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4832__CLK clknet_leaf_20_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3241_ tms1x00.RAM\[116\]\[1\] _1459_ _1475_ vssd1 vssd1 vccd1 vccd1 _1477_ sky130_fd_sc_hd__mux2_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3172_ tms1x00.RAM\[123\]\[0\] _1324_ _1436_ vssd1 vssd1 vccd1 vccd1 _1437_ sky130_fd_sc_hd__mux2_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4982__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5101__A net54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2956_ tms1x00.RAM\[104\]\[0\] _1235_ _1304_ vssd1 vssd1 vccd1 vccd1 _1305_ sky130_fd_sc_hd__mux2_1
X_2887_ _1263_ vssd1 vssd1 vccd1 vccd1 _0067_ sky130_fd_sc_hd__clkbuf_1
X_4626_ clknet_leaf_10_wb_clk_i _0247_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[31\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2408__S1 _0800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4557_ clknet_leaf_13_wb_clk_i _0178_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[124\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2733__A1 _0776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3508_ _1631_ vssd1 vssd1 vccd1 vccd1 _0320_ sky130_fd_sc_hd__clkbuf_1
XFILLER_1_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4488_ clknet_leaf_29_wb_clk_i _0109_ vssd1 vssd1 vccd1 vccd1 tms1x00.RAM\[101\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_58_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3439_ _1592_ tms1x00.RAM\[3\]\[3\] _1586_ vssd1 vssd1 vccd1 vccd1 _1593_ sky130_fd_sc_hd__mux2_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2592__S0 _0975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2354__B _0748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4705__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2647__S1 _0831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2421__B1 _0813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4855__CLK clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3921__A0 _1821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2724__A1 _0944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput85 net85 vssd1 vssd1 vccd1 vccd1 io_out[26] sky130_fd_sc_hd__buf_2
Xoutput74 net74 vssd1 vssd1 vccd1 vccd1 io_out[15] sky130_fd_sc_hd__buf_2
Xoutput96 net96 vssd1 vssd1 vccd1 vccd1 oram_addr[1] sky130_fd_sc_hd__buf_2
XFILLER_1_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3790_ _1793_ vssd1 vssd1 vccd1 vccd1 _0440_ sky130_fd_sc_hd__clkbuf_1
X_2810_ tms1x00.RAM\[36\]\[3\] tms1x00.RAM\[37\]\[3\] tms1x00.RAM\[38\]\[3\] tms1x00.RAM\[39\]\[3\]
+ _0816_ _0927_ vssd1 vssd1 vccd1 vccd1 _1200_ sky130_fd_sc_hd__mux4_1
X_2741_ _1131_ vssd1 vssd1 vccd1 vccd1 _0053_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2672_ tms1x00.RAM\[28\]\[2\] tms1x00.RAM\[29\]\[2\] _0789_ vssd1 vssd1 vccd1 vccd1
+ _1063_ sky130_fd_sc_hd__mux2_1
XFILLER_8_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4411_ clknet_leaf_27_wb_clk_i _0009_ vssd1 vssd1 vccd1 vccd1 wbs_o_buff\[15\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__3912__A0 _1821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2715__A1 _0945_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4342_ _1243_ tms1x00.RAM\[1\]\[1\] _2151_ vssd1 vssd1 vccd1 vccd1 _2153_ sky130_fd_sc_hd__mux2_1
XANTENNA__2810__S1 _0927_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4273_ _2114_ vssd1 vssd1 vccd1 vccd1 _0602_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5010__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3224_ _1467_ vssd1 vssd1 vccd1 vccd1 _0200_ sky130_fd_sc_hd__clkbuf_1
XTAP_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3315__S _1519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
.ends

