* NGSPICE file created from tms1x00_ram.ext - technology: sky130B

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

.subckt tms1x00_ram clk r_val[0] r_val[1] r_val[2] r_val[3] ram_addr[0] ram_addr[1]
+ ram_addr[2] ram_addr[3] ram_addr[4] ram_addr[5] ram_addr[6] vccd1 vssd1 w_val[0]
+ w_val[1] w_val[2] w_val[3] wen
XTAP_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2106_ _2367_/CLK _2106_/D vssd1 vssd1 vccd1 vccd1 _2106_/Q sky130_fd_sc_hd__dfxtp_1
X_2037_ _2049_/CLK _2037_/D vssd1 vssd1 vccd1 vccd1 _2037_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1270_ _2185_/Q _2225_/Q _1270_/S vssd1 vssd1 vccd1 vccd1 _1270_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1606_ _1646_/A _1926_/B vssd1 vssd1 vccd1 vccd1 _1610_/S sky130_fd_sc_hd__nor2_2
X_1537_ _2138_/Q _1582_/A0 _1540_/S vssd1 vssd1 vccd1 vccd1 _2138_/D sky130_fd_sc_hd__mux2_1
Xfanout127 input10/X vssd1 vssd1 vccd1 vccd1 fanout127/X sky130_fd_sc_hd__buf_4
Xfanout138 fanout148/X vssd1 vssd1 vccd1 vccd1 _1285_/S0 sky130_fd_sc_hd__buf_8
Xfanout105 _1740_/A0 vssd1 vssd1 vccd1 vccd1 _1935_/A0 sky130_fd_sc_hd__buf_4
Xfanout116 _1784_/A0 vssd1 vssd1 vccd1 vccd1 _1824_/A0 sky130_fd_sc_hd__buf_4
X_1468_ _2084_/Q _1809_/A0 _1469_/S vssd1 vssd1 vccd1 vccd1 _2084_/D sky130_fd_sc_hd__mux2_1
X_1399_ _1966_/B _1981_/B vssd1 vssd1 vccd1 vccd1 _1403_/S sky130_fd_sc_hd__nor2_2
XFILLER_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_283 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2440_ _2448_/CLK _2440_/D vssd1 vssd1 vccd1 vccd1 _2440_/Q sky130_fd_sc_hd__dfxtp_1
X_2371_ _2433_/CLK _2371_/D vssd1 vssd1 vccd1 vccd1 _2371_/Q sky130_fd_sc_hd__dfxtp_1
X_1322_ _1322_/A _1385_/B vssd1 vssd1 vccd1 vccd1 _1806_/A sky130_fd_sc_hd__or2_4
X_1253_ _2373_/Q _2377_/Q _2381_/Q _2021_/Q _1253_/S0 _1253_/S1 vssd1 vssd1 vccd1
+ vccd1 _1253_/X sky130_fd_sc_hd__mux4_1
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1184_ _0992_/A _1182_/X _1183_/X vssd1 vssd1 vccd1 vccd1 _1184_/X sky130_fd_sc_hd__a21o_1
XFILLER_64_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1940_ _1940_/A0 _2461_/Q _1940_/S vssd1 vssd1 vccd1 vccd1 _2461_/D sky130_fd_sc_hd__mux2_1
XFILLER_14_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1871_ _1951_/A _1901_/B vssd1 vssd1 vccd1 vccd1 _1875_/S sky130_fd_sc_hd__nand2_4
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2423_ _2495_/CLK _2423_/D vssd1 vssd1 vccd1 vccd1 _2423_/Q sky130_fd_sc_hd__dfxtp_1
X_2354_ _2369_/CLK _2354_/D vssd1 vssd1 vccd1 vccd1 _2354_/Q sky130_fd_sc_hd__dfxtp_1
X_1305_ _1023_/X _1303_/X _1304_/X _1305_/B2 vssd1 vssd1 vccd1 vccd1 _1305_/X sky130_fd_sc_hd__a22o_1
X_2285_ _2416_/CLK _2285_/D vssd1 vssd1 vccd1 vccd1 _2285_/Q sky130_fd_sc_hd__dfxtp_1
X_1236_ _2245_/Q _2249_/Q _2253_/Q _2257_/Q _1245_/S0 _1174_/A vssd1 vssd1 vccd1 vccd1
+ _1237_/B sky130_fd_sc_hd__mux4_1
XFILLER_37_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1167_ _1453_/C _1165_/X _1166_/X _1464_/C vssd1 vssd1 vccd1 vccd1 _1167_/X sky130_fd_sc_hd__o22a_1
XFILLER_52_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1098_ input5/X _1096_/Y _1097_/Y vssd1 vssd1 vccd1 vccd1 _1098_/X sky130_fd_sc_hd__a21o_1
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2070_ _2337_/CLK _2070_/D vssd1 vssd1 vccd1 vccd1 _2070_/Q sky130_fd_sc_hd__dfxtp_1
X_1021_ _1220_/A _1024_/B vssd1 vssd1 vccd1 vccd1 _1475_/C sky130_fd_sc_hd__nand2b_4
XFILLER_46_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1923_ _1978_/A0 _2447_/Q _1925_/S vssd1 vssd1 vccd1 vccd1 _2447_/D sky130_fd_sc_hd__mux2_1
X_1854_ _1969_/A0 _2392_/Q _1855_/S vssd1 vssd1 vccd1 vccd1 _2392_/D sky130_fd_sc_hd__mux2_1
X_1785_ _1800_/A0 _2337_/Q _1785_/S vssd1 vssd1 vccd1 vccd1 _2337_/D sky130_fd_sc_hd__mux2_1
X_2406_ _2481_/CLK _2406_/D vssd1 vssd1 vccd1 vccd1 _2406_/Q sky130_fd_sc_hd__dfxtp_1
X_2337_ _2337_/CLK _2337_/D vssd1 vssd1 vccd1 vccd1 _2337_/Q sky130_fd_sc_hd__dfxtp_1
X_2268_ _2301_/CLK _2268_/D vssd1 vssd1 vccd1 vccd1 _2268_/Q sky130_fd_sc_hd__dfxtp_1
X_1219_ _2148_/Q _2152_/Q _2156_/Q _2160_/Q _1292_/S _1291_/A vssd1 vssd1 vccd1 vccd1
+ _1220_/B sky130_fd_sc_hd__mux4_1
XFILLER_37_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2199_ _2461_/CLK _2199_/D vssd1 vssd1 vccd1 vccd1 _2199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1570_ _2165_/Q _1585_/A0 _1570_/S vssd1 vssd1 vccd1 vccd1 _2165_/D sky130_fd_sc_hd__mux2_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2122_ _2232_/CLK _2122_/D vssd1 vssd1 vccd1 vccd1 _2122_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2053_ _2094_/CLK _2053_/D vssd1 vssd1 vccd1 vccd1 _2053_/Q sky130_fd_sc_hd__dfxtp_1
X_1004_ _2298_/Q _2010_/Q _1240_/S vssd1 vssd1 vccd1 vccd1 _1004_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1906_ _1966_/A _1906_/B vssd1 vssd1 vccd1 vccd1 _1910_/S sky130_fd_sc_hd__nor2_2
X_1837_ _2378_/Q _1972_/A0 _1840_/S vssd1 vssd1 vccd1 vccd1 _2378_/D sky130_fd_sc_hd__mux2_1
X_1768_ _2323_/Q _1783_/A0 _1770_/S vssd1 vssd1 vccd1 vccd1 _2323_/D sky130_fd_sc_hd__mux2_1
X_1699_ _2268_/Q _1739_/A0 _1700_/S vssd1 vssd1 vccd1 vccd1 _2268_/D sky130_fd_sc_hd__mux2_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1622_ _1917_/A1 _2206_/Q _1625_/S vssd1 vssd1 vccd1 vccd1 _2206_/D sky130_fd_sc_hd__mux2_1
X_1553_ _2151_/Q _1918_/A1 _1555_/S vssd1 vssd1 vccd1 vccd1 _2151_/D sky130_fd_sc_hd__mux2_1
X_1484_ _1824_/A0 _2096_/Q _1485_/S vssd1 vssd1 vccd1 vccd1 _2096_/D sky130_fd_sc_hd__mux2_1
XFILLER_39_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2105_ _2385_/CLK _2105_/D vssd1 vssd1 vccd1 vccd1 _2105_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2036_ _2049_/CLK _2036_/D vssd1 vssd1 vccd1 vccd1 _2036_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1605_ _1765_/A0 _2193_/Q _1605_/S vssd1 vssd1 vccd1 vccd1 _2193_/D sky130_fd_sc_hd__mux2_1
X_1536_ _1566_/A _1936_/B vssd1 vssd1 vccd1 vccd1 _1540_/S sky130_fd_sc_hd__nor2_4
Xfanout128 _1420_/A vssd1 vssd1 vccd1 vccd1 _1297_/S0 sky130_fd_sc_hd__buf_8
Xfanout117 _1784_/A0 vssd1 vssd1 vccd1 vccd1 _1809_/A0 sky130_fd_sc_hd__buf_4
Xfanout106 _1845_/A1 vssd1 vssd1 vccd1 vccd1 _1985_/A1 sky130_fd_sc_hd__clkbuf_4
X_1467_ _2083_/Q _1778_/A0 _1469_/S vssd1 vssd1 vccd1 vccd1 _2083_/D sky130_fd_sc_hd__mux2_1
Xfanout139 fanout148/X vssd1 vssd1 vccd1 vccd1 _1453_/A sky130_fd_sc_hd__clkbuf_4
X_1398_ _1398_/A _1398_/B vssd1 vssd1 vccd1 vccd1 _1691_/A sky130_fd_sc_hd__or2_4
XFILLER_82_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2019_ _2485_/CLK _2019_/D vssd1 vssd1 vccd1 vccd1 _2019_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2370_ _2482_/CLK _2370_/D vssd1 vssd1 vccd1 vccd1 _2370_/Q sky130_fd_sc_hd__dfxtp_1
X_1321_ _1322_/A _1385_/B vssd1 vssd1 vccd1 vccd1 _1821_/A sky130_fd_sc_hd__nor2_8
XFILLER_68_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1252_ _2389_/Q _2393_/Q _2397_/Q _2401_/Q _1253_/S0 _1256_/S1 vssd1 vssd1 vccd1
+ vccd1 _1252_/X sky130_fd_sc_hd__mux4_1
XFILLER_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1183_ _1475_/B _1181_/X _1258_/A vssd1 vssd1 vccd1 vccd1 _1183_/X sky130_fd_sc_hd__a21o_1
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1519_ _2124_/Q _1579_/A0 _1520_/S vssd1 vssd1 vccd1 vccd1 _2124_/D sky130_fd_sc_hd__mux2_1
XFILLER_28_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1870_ _2405_/Q _1905_/A0 _1870_/S vssd1 vssd1 vccd1 vccd1 _2405_/D sky130_fd_sc_hd__mux2_1
XFILLER_80_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2422_ _2495_/CLK _2422_/D vssd1 vssd1 vccd1 vccd1 _2422_/Q sky130_fd_sc_hd__dfxtp_1
X_2353_ _2369_/CLK _2353_/D vssd1 vssd1 vccd1 vccd1 _2353_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1304_ _2053_/Q _2057_/Q _2061_/Q _2009_/Q _1304_/S0 _1304_/S1 vssd1 vssd1 vccd1
+ vccd1 _1304_/X sky130_fd_sc_hd__mux4_1
X_2284_ _2481_/CLK _2284_/D vssd1 vssd1 vccd1 vccd1 _2284_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1235_ _1174_/A _1232_/X _1234_/X vssd1 vssd1 vccd1 vccd1 _1235_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_25_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1166_ _2468_/Q _2472_/Q _2476_/Q _2480_/Q _1475_/A _1464_/B vssd1 vssd1 vccd1 vccd1
+ _1166_/X sky130_fd_sc_hd__mux4_2
XFILLER_64_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1097_ input5/X _1090_/X input6/X vssd1 vssd1 vccd1 vccd1 _1097_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_52_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1999_ _2241_/CLK _1999_/D vssd1 vssd1 vccd1 vccd1 _1999_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1020_ _1020_/A _1023_/B vssd1 vssd1 vccd1 vccd1 _1020_/X sky130_fd_sc_hd__and2_4
XFILLER_19_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1922_ _1977_/A0 _2446_/Q _1925_/S vssd1 vssd1 vccd1 vccd1 _2446_/D sky130_fd_sc_hd__mux2_1
X_1853_ _1903_/A0 _2391_/Q _1855_/S vssd1 vssd1 vccd1 vccd1 _2391_/D sky130_fd_sc_hd__mux2_1
X_1784_ _1784_/A0 _2336_/Q _1785_/S vssd1 vssd1 vccd1 vccd1 _2336_/D sky130_fd_sc_hd__mux2_1
X_2405_ _2432_/CLK _2405_/D vssd1 vssd1 vccd1 vccd1 _2405_/Q sky130_fd_sc_hd__dfxtp_1
X_2336_ _2337_/CLK _2336_/D vssd1 vssd1 vccd1 vccd1 _2336_/Q sky130_fd_sc_hd__dfxtp_1
X_2267_ _2301_/CLK _2267_/D vssd1 vssd1 vccd1 vccd1 _2267_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1218_ _2164_/Q _2168_/Q _2172_/Q _2176_/Q _1297_/S0 _1297_/S1 vssd1 vssd1 vccd1
+ vccd1 _1218_/X sky130_fd_sc_hd__mux4_1
XFILLER_72_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2198_ _2461_/CLK _2198_/D vssd1 vssd1 vccd1 vccd1 _2198_/Q sky130_fd_sc_hd__dfxtp_1
X_1149_ _2323_/Q _2327_/Q _2331_/Q _2335_/Q _1275_/S0 _1065_/A vssd1 vssd1 vccd1 vccd1
+ _1149_/X sky130_fd_sc_hd__mux4_2
XFILLER_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2121_ _2449_/CLK _2121_/D vssd1 vssd1 vccd1 vccd1 _2121_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2052_ _2094_/CLK _2052_/D vssd1 vssd1 vccd1 vccd1 _2052_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1003_ _2290_/Q _2294_/Q _1240_/S vssd1 vssd1 vccd1 vccd1 _1003_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1905_ _1905_/A0 _2433_/Q _1905_/S vssd1 vssd1 vccd1 vccd1 _2433_/D sky130_fd_sc_hd__mux2_1
X_1836_ _1886_/A _1916_/B vssd1 vssd1 vccd1 vccd1 _1840_/S sky130_fd_sc_hd__nor2_2
X_1767_ _2322_/Q _1842_/A1 _1770_/S vssd1 vssd1 vccd1 vccd1 _2322_/D sky130_fd_sc_hd__mux2_1
X_1698_ _2267_/Q _1793_/A1 _1700_/S vssd1 vssd1 vccd1 vccd1 _2267_/D sky130_fd_sc_hd__mux2_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2319_ _2363_/CLK _2319_/D vssd1 vssd1 vccd1 vccd1 _2319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1621_ _1661_/A _1861_/A vssd1 vssd1 vccd1 vccd1 _1625_/S sky130_fd_sc_hd__nand2_2
X_1552_ _2150_/Q _1977_/A0 _1555_/S vssd1 vssd1 vccd1 vccd1 _2150_/D sky130_fd_sc_hd__mux2_1
X_1483_ _1778_/A0 _2095_/Q _1485_/S vssd1 vssd1 vccd1 vccd1 _2095_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2104_ _2496_/CLK _2104_/D vssd1 vssd1 vccd1 vccd1 _2104_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2035_ _2049_/CLK _2035_/D vssd1 vssd1 vccd1 vccd1 _2035_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1819_ _1824_/A0 _2364_/Q _1820_/S vssd1 vssd1 vccd1 vccd1 _2364_/D sky130_fd_sc_hd__mux2_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1604_ _1814_/A0 _2192_/Q _1605_/S vssd1 vssd1 vccd1 vccd1 _2192_/D sky130_fd_sc_hd__mux2_1
X_1535_ _2137_/Q _1660_/A0 _1535_/S vssd1 vssd1 vccd1 vccd1 _2137_/D sky130_fd_sc_hd__mux2_1
Xfanout129 _1420_/A vssd1 vssd1 vccd1 vccd1 _1292_/S sky130_fd_sc_hd__buf_6
Xfanout118 fanout127/X vssd1 vssd1 vccd1 vccd1 _1784_/A0 sky130_fd_sc_hd__clkbuf_4
Xfanout107 _1740_/A0 vssd1 vssd1 vccd1 vccd1 _1845_/A1 sky130_fd_sc_hd__buf_4
X_1466_ _2082_/Q _1777_/A0 _1469_/S vssd1 vssd1 vccd1 vccd1 _2082_/D sky130_fd_sc_hd__mux2_1
X_1397_ _1398_/A _1398_/B vssd1 vssd1 vccd1 vccd1 _1941_/B sky130_fd_sc_hd__nor2_8
XFILLER_82_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2018_ _2477_/CLK _2018_/D vssd1 vssd1 vccd1 vccd1 _2018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1320_ _1366_/A _1475_/C vssd1 vssd1 vccd1 vccd1 _1981_/A sky130_fd_sc_hd__or2_4
XFILLER_78_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1251_ _1420_/C _1247_/X _1250_/X _1246_/X vssd1 vssd1 vccd1 vccd1 _1251_/X sky130_fd_sc_hd__o211a_1
XFILLER_83_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1182_ _2300_/Q _2012_/Q _1182_/S vssd1 vssd1 vccd1 vccd1 _1182_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1518_ _2123_/Q _1583_/A0 _1520_/S vssd1 vssd1 vccd1 vccd1 _2123_/D sky130_fd_sc_hd__mux2_1
X_1449_ _2070_/Q _1822_/A0 _1452_/S vssd1 vssd1 vccd1 vccd1 _2070_/D sky130_fd_sc_hd__mux2_1
XFILLER_28_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2421_ _2421_/CLK _2421_/D vssd1 vssd1 vccd1 vccd1 _2421_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2352_ _2457_/CLK _2352_/D vssd1 vssd1 vccd1 vccd1 _2352_/Q sky130_fd_sc_hd__dfxtp_1
X_2283_ _2481_/CLK _2283_/D vssd1 vssd1 vccd1 vccd1 _2283_/Q sky130_fd_sc_hd__dfxtp_1
X_1303_ _2101_/Q _2017_/Q _2109_/Q _2113_/Q _1303_/S0 _1304_/S1 vssd1 vssd1 vccd1
+ vccd1 _1303_/X sky130_fd_sc_hd__mux4_1
XFILLER_56_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1234_ _1234_/A1 _1233_/X _1241_/B1 vssd1 vssd1 vccd1 vccd1 _1234_/X sky130_fd_sc_hd__a21o_1
XFILLER_84_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1165_ _2452_/Q _2456_/Q _2460_/Q _2028_/Q _1475_/A _1464_/B vssd1 vssd1 vccd1 vccd1
+ _1165_/X sky130_fd_sc_hd__mux4_1
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1096_ _1396_/C _1094_/X _1095_/X _1420_/C _1093_/X vssd1 vssd1 vccd1 vccd1 _1096_/Y
+ sky130_fd_sc_hd__o221ai_4
XFILLER_52_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1998_ _2241_/CLK _1998_/D vssd1 vssd1 vccd1 vccd1 _1998_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1921_ _1921_/A _1976_/A vssd1 vssd1 vccd1 vccd1 _1925_/S sky130_fd_sc_hd__nand2_2
XFILLER_42_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1852_ _1902_/A0 _2390_/Q _1855_/S vssd1 vssd1 vccd1 vccd1 _2390_/D sky130_fd_sc_hd__mux2_1
X_1783_ _1783_/A0 _2335_/Q _1785_/S vssd1 vssd1 vccd1 vccd1 _2335_/D sky130_fd_sc_hd__mux2_1
XFILLER_6_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2404_ _2416_/CLK _2404_/D vssd1 vssd1 vccd1 vccd1 _2404_/Q sky130_fd_sc_hd__dfxtp_1
X_2335_ _2335_/CLK _2335_/D vssd1 vssd1 vccd1 vccd1 _2335_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2266_ _2343_/CLK _2266_/D vssd1 vssd1 vccd1 vccd1 _2266_/Q sky130_fd_sc_hd__dfxtp_1
X_1217_ _1298_/B2 _1215_/X _1216_/X _1295_/B2 vssd1 vssd1 vccd1 vccd1 _1217_/X sky130_fd_sc_hd__a22o_1
X_2197_ _2368_/CLK _2197_/D vssd1 vssd1 vccd1 vccd1 _2197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1148_ _1037_/X _1147_/X _1139_/X vssd1 vssd1 vccd1 vccd1 _1148_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_80_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1079_ _1298_/B2 _1077_/X _1078_/X _1020_/X vssd1 vssd1 vccd1 vccd1 _1079_/X sky130_fd_sc_hd__a22o_1
XFILLER_52_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2120_ _2176_/CLK _2120_/D vssd1 vssd1 vccd1 vccd1 _2120_/Q sky130_fd_sc_hd__dfxtp_1
X_2051_ _2094_/CLK _2051_/D vssd1 vssd1 vccd1 vccd1 _2051_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1002_ _2274_/Q _2278_/Q _2282_/Q _2286_/Q _1181_/S _0992_/A vssd1 vssd1 vccd1 vccd1
+ _1002_/X sky130_fd_sc_hd__mux4_1
XFILLER_47_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1904_ _1904_/A0 _2432_/Q _1905_/S vssd1 vssd1 vccd1 vccd1 _2432_/D sky130_fd_sc_hd__mux2_1
XFILLER_30_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1835_ _2377_/Q _1975_/A0 _1835_/S vssd1 vssd1 vccd1 vccd1 _2377_/D sky130_fd_sc_hd__mux2_1
X_1766_ _1806_/A _1926_/B vssd1 vssd1 vccd1 vccd1 _1770_/S sky130_fd_sc_hd__nor2_2
X_1697_ _2266_/Q _1792_/A1 _1700_/S vssd1 vssd1 vccd1 vccd1 _2266_/D sky130_fd_sc_hd__mux2_1
XFILLER_85_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2318_ _2320_/CLK _2318_/D vssd1 vssd1 vccd1 vccd1 _2318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2249_ _2343_/CLK _2249_/D vssd1 vssd1 vccd1 vccd1 _2249_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1620_ _1765_/A0 _2205_/Q _1620_/S vssd1 vssd1 vccd1 vccd1 _2205_/D sky130_fd_sc_hd__mux2_1
X_1551_ _1981_/A _1566_/A vssd1 vssd1 vccd1 vccd1 _1555_/S sky130_fd_sc_hd__nor2_4
X_1482_ _1777_/A0 _2094_/Q _1485_/S vssd1 vssd1 vccd1 vccd1 _2094_/D sky130_fd_sc_hd__mux2_1
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2103_ _2385_/CLK _2103_/D vssd1 vssd1 vccd1 vccd1 _2103_/Q sky130_fd_sc_hd__dfxtp_1
X_2034_ _2049_/CLK _2034_/D vssd1 vssd1 vccd1 vccd1 _2034_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1818_ _1823_/A0 _2363_/Q _1820_/S vssd1 vssd1 vccd1 vccd1 _2363_/D sky130_fd_sc_hd__mux2_1
X_1749_ _2308_/Q _1814_/A0 _1750_/S vssd1 vssd1 vccd1 vccd1 _2308_/D sky130_fd_sc_hd__mux2_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_283 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1603_ _1663_/A0 _2191_/Q _1605_/S vssd1 vssd1 vccd1 vccd1 _2191_/D sky130_fd_sc_hd__mux2_1
X_1534_ _2136_/Q _1579_/A0 _1535_/S vssd1 vssd1 vccd1 vccd1 _2136_/D sky130_fd_sc_hd__mux2_1
Xfanout119 _1884_/A0 vssd1 vssd1 vccd1 vccd1 _1969_/A0 sky130_fd_sc_hd__buf_4
Xfanout108 fanout109/X vssd1 vssd1 vccd1 vccd1 _1740_/A0 sky130_fd_sc_hd__clkbuf_4
X_1465_ _1486_/A _1946_/B vssd1 vssd1 vccd1 vccd1 _1469_/S sky130_fd_sc_hd__nor2_2
X_1396_ _1464_/A _1442_/B _1396_/C vssd1 vssd1 vccd1 vccd1 _1966_/B sky130_fd_sc_hd__or3_4
X_2017_ _2367_/CLK _2017_/D vssd1 vssd1 vccd1 vccd1 _2017_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1250_ _1464_/C _1248_/X _1249_/X _1396_/C vssd1 vssd1 vccd1 vccd1 _1250_/X sky130_fd_sc_hd__o22a_1
X_1181_ _2292_/Q _2296_/Q _1181_/S vssd1 vssd1 vccd1 vccd1 _1181_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1517_ _2122_/Q _1582_/A0 _1520_/S vssd1 vssd1 vccd1 vccd1 _2122_/D sky130_fd_sc_hd__mux2_1
X_2497_ _2497_/CLK _2497_/D vssd1 vssd1 vccd1 vccd1 _2497_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1448_ _1641_/A _1486_/A vssd1 vssd1 vccd1 vccd1 _1452_/S sky130_fd_sc_hd__nor2_2
X_1379_ _1971_/A _1901_/B vssd1 vssd1 vccd1 vccd1 _1383_/S sky130_fd_sc_hd__nand2_2
XFILLER_82_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout90 fanout94/X vssd1 vssd1 vccd1 vccd1 _1409_/B sky130_fd_sc_hd__clkbuf_8
X_2420_ _2421_/CLK _2420_/D vssd1 vssd1 vccd1 vccd1 _2420_/Q sky130_fd_sc_hd__dfxtp_1
X_2351_ _2369_/CLK _2351_/D vssd1 vssd1 vccd1 vccd1 _2351_/Q sky130_fd_sc_hd__dfxtp_1
X_2282_ _2481_/CLK _2282_/D vssd1 vssd1 vccd1 vccd1 _2282_/Q sky130_fd_sc_hd__dfxtp_1
X_1302_ _1302_/A1 _1300_/X _1301_/X _1020_/X vssd1 vssd1 vccd1 vccd1 _1302_/X sky130_fd_sc_hd__a22o_1
XFILLER_84_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1233_ _2261_/Q _1989_/Q _1233_/S vssd1 vssd1 vccd1 vccd1 _1233_/X sky130_fd_sc_hd__mux2_1
X_1164_ _1295_/B2 _1158_/X _1163_/X _1298_/B2 vssd1 vssd1 vccd1 vccd1 _1164_/X sky130_fd_sc_hd__a22o_1
XFILLER_37_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1095_ _2179_/Q _1999_/Q _2187_/Q _2191_/Q _1287_/S0 _1013_/B vssd1 vssd1 vccd1 vccd1
+ _1095_/X sky130_fd_sc_hd__mux4_2
XFILLER_64_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1997_ _2229_/CLK _1997_/D vssd1 vssd1 vccd1 vccd1 _1997_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1920_ _2445_/Q _1980_/A0 _1920_/S vssd1 vssd1 vccd1 vccd1 _2445_/D sky130_fd_sc_hd__mux2_1
XFILLER_61_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1851_ _1931_/A _1901_/B vssd1 vssd1 vccd1 vccd1 _1855_/S sky130_fd_sc_hd__nand2_4
X_1782_ _1842_/A1 _2334_/Q _1785_/S vssd1 vssd1 vccd1 vccd1 _2334_/D sky130_fd_sc_hd__mux2_1
X_2403_ _2432_/CLK _2403_/D vssd1 vssd1 vccd1 vccd1 _2403_/Q sky130_fd_sc_hd__dfxtp_1
X_2334_ _2337_/CLK _2334_/D vssd1 vssd1 vccd1 vccd1 _2334_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2265_ _2496_/CLK _2265_/D vssd1 vssd1 vccd1 vccd1 _2265_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1216_ _2116_/Q _2120_/Q _2124_/Q _2128_/Q _1297_/S0 _1297_/S1 vssd1 vssd1 vccd1
+ vccd1 _1216_/X sky130_fd_sc_hd__mux4_1
X_2196_ _2461_/CLK _2196_/D vssd1 vssd1 vccd1 vccd1 _2196_/Q sky130_fd_sc_hd__dfxtp_1
X_1147_ _1024_/B _1145_/X _1146_/X _1143_/X vssd1 vssd1 vccd1 vccd1 _1147_/X sky130_fd_sc_hd__a31o_1
XFILLER_1_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1078_ _2082_/Q _2086_/Q _2090_/Q _2094_/Q _1303_/S0 _1304_/S1 vssd1 vssd1 vccd1
+ vccd1 _1078_/X sky130_fd_sc_hd__mux4_1
XFILLER_52_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2050_ _2094_/CLK _2050_/D vssd1 vssd1 vccd1 vccd1 _2050_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1001_ _1237_/A _1001_/B vssd1 vssd1 vccd1 vccd1 _1001_/Y sky130_fd_sc_hd__nor2_1
XFILLER_47_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1903_ _1903_/A0 _2431_/Q _1905_/S vssd1 vssd1 vccd1 vccd1 _2431_/D sky130_fd_sc_hd__mux2_1
XFILLER_30_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1834_ _2376_/Q _1969_/A0 _1835_/S vssd1 vssd1 vccd1 vccd1 _2376_/D sky130_fd_sc_hd__mux2_1
XFILLER_30_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1765_ _1765_/A0 _2321_/Q _1765_/S vssd1 vssd1 vccd1 vccd1 _2321_/D sky130_fd_sc_hd__mux2_1
X_1696_ _1726_/A _1936_/B vssd1 vssd1 vccd1 vccd1 _1700_/S sky130_fd_sc_hd__nor2_4
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2317_ _2363_/CLK _2317_/D vssd1 vssd1 vccd1 vccd1 _2317_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2248_ _2480_/CLK _2248_/D vssd1 vssd1 vccd1 vccd1 _2248_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2179_ _2241_/CLK _2179_/D vssd1 vssd1 vccd1 vccd1 _2179_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_52 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1550_ _2149_/Q _1980_/A0 _1550_/S vssd1 vssd1 vccd1 vccd1 _2149_/D sky130_fd_sc_hd__mux2_1
X_1481_ _1961_/A _1501_/A vssd1 vssd1 vccd1 vccd1 _1485_/S sky130_fd_sc_hd__nand2_4
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2102_ _2329_/CLK _2102_/D vssd1 vssd1 vccd1 vccd1 _2102_/Q sky130_fd_sc_hd__dfxtp_1
X_2033_ _2493_/CLK _2033_/D vssd1 vssd1 vccd1 vccd1 _2033_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1817_ _1822_/A0 _2362_/Q _1820_/S vssd1 vssd1 vccd1 vccd1 _2362_/D sky130_fd_sc_hd__mux2_1
X_1748_ _2307_/Q _1823_/A0 _1750_/S vssd1 vssd1 vccd1 vccd1 _2307_/D sky130_fd_sc_hd__mux2_1
X_1679_ _2252_/Q _1804_/A0 _1680_/S vssd1 vssd1 vccd1 vccd1 _2252_/D sky130_fd_sc_hd__mux2_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1602_ _1662_/A0 _2190_/Q _1605_/S vssd1 vssd1 vccd1 vccd1 _2190_/D sky130_fd_sc_hd__mux2_1
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1533_ _2135_/Q _1583_/A0 _1535_/S vssd1 vssd1 vccd1 vccd1 _2135_/D sky130_fd_sc_hd__mux2_1
X_1464_ _1464_/A _1464_/B _1464_/C vssd1 vssd1 vccd1 vccd1 _1946_/B sky130_fd_sc_hd__or3_4
Xfanout109 _1965_/A0 vssd1 vssd1 vccd1 vccd1 fanout109/X sky130_fd_sc_hd__clkbuf_4
X_1395_ _1980_/A0 _2033_/Q _1395_/S vssd1 vssd1 vccd1 vccd1 _2033_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2016_ _2363_/CLK _2016_/D vssd1 vssd1 vccd1 vccd1 _2016_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_30_clk clkbuf_2_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _2296_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_21_clk clkbuf_2_3__f_clk/X vssd1 vssd1 vccd1 vccd1 _2496_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_5_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1180_ _1180_/A _1180_/B vssd1 vssd1 vccd1 vccd1 _1180_/X sky130_fd_sc_hd__or2_1
XFILLER_76_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_12_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _2335_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_9_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1516_ _1566_/A _1916_/B vssd1 vssd1 vccd1 vccd1 _1520_/S sky130_fd_sc_hd__nor2_2
X_2496_ _2496_/CLK _2496_/D vssd1 vssd1 vccd1 vccd1 _2496_/Q sky130_fd_sc_hd__dfxtp_1
X_1447_ _2069_/Q _1800_/A0 _1447_/S vssd1 vssd1 vccd1 vccd1 _2069_/D sky130_fd_sc_hd__mux2_1
X_1378_ _1975_/A0 _2021_/Q _1378_/S vssd1 vssd1 vccd1 vccd1 _2021_/D sky130_fd_sc_hd__mux2_1
XFILLER_63_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout80 fanout85/X vssd1 vssd1 vccd1 vccd1 _1442_/B sky130_fd_sc_hd__buf_4
Xfanout91 fanout94/X vssd1 vssd1 vccd1 vccd1 _1174_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_80_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2350_ _2369_/CLK _2350_/D vssd1 vssd1 vccd1 vccd1 _2350_/Q sky130_fd_sc_hd__dfxtp_1
X_2281_ _2296_/CLK _2281_/D vssd1 vssd1 vccd1 vccd1 _2281_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1301_ _2085_/Q _2089_/Q _2093_/Q _2097_/Q _1303_/S0 _1301_/S1 vssd1 vssd1 vccd1
+ vccd1 _1301_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_1_clk clkbuf_leaf_4_clk/A vssd1 vssd1 vccd1 vccd1 _2240_/CLK sky130_fd_sc_hd__clkbuf_16
X_1232_ _2269_/Q _2273_/Q _1240_/S vssd1 vssd1 vccd1 vccd1 _1232_/X sky130_fd_sc_hd__mux2_1
X_1163_ _2388_/Q _2392_/Q _2396_/Q _2400_/Q _1253_/S0 _1253_/S1 vssd1 vssd1 vccd1
+ vccd1 _1163_/X sky130_fd_sc_hd__mux4_1
XFILLER_64_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1094_ _2227_/Q _2231_/Q _2235_/Q _2239_/Q _1287_/S0 _1013_/B vssd1 vssd1 vccd1 vccd1
+ _1094_/X sky130_fd_sc_hd__mux4_2
XFILLER_64_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1996_ _2229_/CLK _1996_/D vssd1 vssd1 vccd1 vccd1 _1996_/Q sky130_fd_sc_hd__dfxtp_1
X_2479_ _2479_/CLK _2479_/D vssd1 vssd1 vccd1 vccd1 _2479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1850_ _2389_/Q _1905_/A0 _1850_/S vssd1 vssd1 vccd1 vccd1 _2389_/D sky130_fd_sc_hd__mux2_1
X_1781_ _1821_/A _1861_/A vssd1 vssd1 vccd1 vccd1 _1785_/S sky130_fd_sc_hd__nand2_2
XFILLER_6_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2402_ _2481_/CLK _2402_/D vssd1 vssd1 vccd1 vccd1 _2402_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2333_ _2337_/CLK _2333_/D vssd1 vssd1 vccd1 vccd1 _2333_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2264_ _2496_/CLK _2264_/D vssd1 vssd1 vccd1 vccd1 _2264_/Q sky130_fd_sc_hd__dfxtp_1
X_1215_ _2132_/Q _2136_/Q _2140_/Q _2004_/Q _1297_/S0 _1297_/S1 vssd1 vssd1 vccd1
+ vccd1 _1215_/X sky130_fd_sc_hd__mux4_1
XFILLER_37_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2195_ _2461_/CLK _2195_/D vssd1 vssd1 vccd1 vccd1 _2195_/Q sky130_fd_sc_hd__dfxtp_1
X_1146_ _1258_/A _1146_/B vssd1 vssd1 vccd1 vccd1 _1146_/X sky130_fd_sc_hd__or2_1
XFILLER_1_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1077_ _2066_/Q _2070_/Q _2074_/Q _2078_/Q _1304_/S0 _1304_/S1 vssd1 vssd1 vccd1
+ vccd1 _1077_/X sky130_fd_sc_hd__mux4_1
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1979_ _1979_/A0 _2492_/Q _1980_/S vssd1 vssd1 vccd1 vccd1 _2492_/D sky130_fd_sc_hd__mux2_1
XFILLER_4_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1000_ _2242_/Q _2246_/Q _2250_/Q _2254_/Q _1245_/S0 _1409_/B vssd1 vssd1 vccd1 vccd1
+ _1001_/B sky130_fd_sc_hd__mux4_1
XFILLER_19_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1902_ _1902_/A0 _2430_/Q _1905_/S vssd1 vssd1 vccd1 vccd1 _2430_/D sky130_fd_sc_hd__mux2_1
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1833_ _2375_/Q _1973_/A0 _1835_/S vssd1 vssd1 vccd1 vccd1 _2375_/D sky130_fd_sc_hd__mux2_1
X_1764_ _1814_/A0 _2320_/Q _1765_/S vssd1 vssd1 vccd1 vccd1 _2320_/D sky130_fd_sc_hd__mux2_1
X_1695_ _2265_/Q _1845_/A1 _1695_/S vssd1 vssd1 vccd1 vccd1 _2265_/D sky130_fd_sc_hd__mux2_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2316_ _2320_/CLK _2316_/D vssd1 vssd1 vccd1 vccd1 _2316_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2247_ _2343_/CLK _2247_/D vssd1 vssd1 vccd1 vccd1 _2247_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2178_ _2241_/CLK _2178_/D vssd1 vssd1 vccd1 vccd1 _2178_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1129_ _1475_/B _1127_/X _1258_/A vssd1 vssd1 vccd1 vccd1 _1129_/X sky130_fd_sc_hd__a21o_1
XFILLER_15_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput13 _1085_/X vssd1 vssd1 vccd1 vccd1 r_val[0] sky130_fd_sc_hd__buf_4
XFILLER_76_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1480_ _2093_/Q _1505_/A0 _1480_/S vssd1 vssd1 vccd1 vccd1 _2093_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2101_ _2367_/CLK _2101_/D vssd1 vssd1 vccd1 vccd1 _2101_/Q sky130_fd_sc_hd__dfxtp_1
X_2032_ _2493_/CLK _2032_/D vssd1 vssd1 vccd1 vccd1 _2032_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1816_ _1821_/A _1976_/B vssd1 vssd1 vccd1 vccd1 _1820_/S sky130_fd_sc_hd__nand2_2
X_1747_ _2306_/Q _1762_/A0 _1750_/S vssd1 vssd1 vccd1 vccd1 _2306_/D sky130_fd_sc_hd__mux2_1
X_1678_ _2251_/Q _1983_/A1 _1680_/S vssd1 vssd1 vccd1 vccd1 _2251_/D sky130_fd_sc_hd__mux2_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1601_ _1661_/A _1921_/A vssd1 vssd1 vccd1 vccd1 _1605_/S sky130_fd_sc_hd__nand2_2
X_1532_ _2134_/Q _1582_/A0 _1535_/S vssd1 vssd1 vccd1 vccd1 _2134_/D sky130_fd_sc_hd__mux2_1
X_1463_ _1800_/A0 _2081_/Q _1463_/S vssd1 vssd1 vccd1 vccd1 _2081_/D sky130_fd_sc_hd__mux2_1
X_1394_ _1974_/A0 _2032_/Q _1395_/S vssd1 vssd1 vccd1 vccd1 _2032_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2015_ _2113_/CLK _2015_/D vssd1 vssd1 vccd1 vccd1 _2015_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1515_ _2121_/Q _1585_/A0 _1515_/S vssd1 vssd1 vccd1 vccd1 _2121_/D sky130_fd_sc_hd__mux2_1
X_2495_ _2495_/CLK _2495_/D vssd1 vssd1 vccd1 vccd1 _2495_/Q sky130_fd_sc_hd__dfxtp_1
X_1446_ _2068_/Q _1809_/A0 _1447_/S vssd1 vssd1 vccd1 vccd1 _2068_/D sky130_fd_sc_hd__mux2_1
X_1377_ _1969_/A0 _2020_/Q _1378_/S vssd1 vssd1 vccd1 vccd1 _2020_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout70 input4/X vssd1 vssd1 vccd1 vccd1 _1024_/B sky130_fd_sc_hd__buf_8
Xfanout81 fanout85/X vssd1 vssd1 vccd1 vccd1 _1253_/S1 sky130_fd_sc_hd__buf_6
Xfanout92 fanout94/X vssd1 vssd1 vccd1 vccd1 _1065_/A sky130_fd_sc_hd__buf_6
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2280_ _2481_/CLK _2280_/D vssd1 vssd1 vccd1 vccd1 _2280_/Q sky130_fd_sc_hd__dfxtp_1
X_1300_ _2069_/Q _2073_/Q _2077_/Q _2081_/Q _1304_/S0 _1301_/S1 vssd1 vssd1 vccd1
+ vccd1 _1300_/X sky130_fd_sc_hd__mux4_1
XFILLER_1_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1231_ _1048_/A _1193_/X _1207_/Y _1230_/X vssd1 vssd1 vccd1 vccd1 _1231_/X sky130_fd_sc_hd__o22a_2
XFILLER_77_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1162_ _1258_/A _1159_/X _1161_/X _1024_/B vssd1 vssd1 vccd1 vccd1 _1162_/X sky130_fd_sc_hd__o211a_1
XFILLER_64_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1093_ _1453_/C _1091_/X _1092_/X _1464_/C vssd1 vssd1 vccd1 vccd1 _1093_/X sky130_fd_sc_hd__o22a_2
XFILLER_60_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1995_ _2229_/CLK _1995_/D vssd1 vssd1 vccd1 vccd1 _1995_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2478_ _2479_/CLK _2478_/D vssd1 vssd1 vccd1 vccd1 _2478_/Q sky130_fd_sc_hd__dfxtp_1
X_1429_ _2056_/Q _1824_/A0 _1430_/S vssd1 vssd1 vccd1 vccd1 _2056_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1780_ _1800_/A0 _2333_/Q _1780_/S vssd1 vssd1 vccd1 vccd1 _2333_/D sky130_fd_sc_hd__mux2_1
X_2401_ _2433_/CLK _2401_/D vssd1 vssd1 vccd1 vccd1 _2401_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2332_ _2337_/CLK _2332_/D vssd1 vssd1 vccd1 vccd1 _2332_/Q sky130_fd_sc_hd__dfxtp_1
X_2263_ _2302_/CLK _2263_/D vssd1 vssd1 vccd1 vccd1 _2263_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2194_ _2461_/CLK _2194_/D vssd1 vssd1 vccd1 vccd1 _2194_/Q sky130_fd_sc_hd__dfxtp_1
X_1214_ _1420_/C _1210_/X _1213_/X _1209_/X vssd1 vssd1 vccd1 vccd1 _1230_/B sky130_fd_sc_hd__o211a_1
XFILLER_80_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1145_ _1220_/A _1145_/B vssd1 vssd1 vccd1 vccd1 _1145_/X sky130_fd_sc_hd__or2_1
XFILLER_25_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1076_ _1244_/A1 _1071_/X _1075_/X _1067_/X _1069_/X vssd1 vssd1 vccd1 vccd1 _1076_/X
+ sky130_fd_sc_hd__a32o_2
XFILLER_80_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1978_ _1978_/A0 _2491_/Q _1980_/S vssd1 vssd1 vccd1 vccd1 _2491_/D sky130_fd_sc_hd__mux2_1
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1901_ _1901_/A _1901_/B vssd1 vssd1 vccd1 vccd1 _1905_/S sky130_fd_sc_hd__nand2_2
XFILLER_30_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1832_ _2374_/Q _1972_/A0 _1835_/S vssd1 vssd1 vccd1 vccd1 _2374_/D sky130_fd_sc_hd__mux2_1
X_1763_ _1823_/A0 _2319_/Q _1765_/S vssd1 vssd1 vccd1 vccd1 _2319_/D sky130_fd_sc_hd__mux2_1
X_1694_ _2264_/Q _1984_/A1 _1695_/S vssd1 vssd1 vccd1 vccd1 _2264_/D sky130_fd_sc_hd__mux2_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2315_ _2363_/CLK _2315_/D vssd1 vssd1 vccd1 vccd1 _2315_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2246_ _2495_/CLK _2246_/D vssd1 vssd1 vccd1 vccd1 _2246_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2177_ _2177_/CLK _2177_/D vssd1 vssd1 vccd1 vccd1 _2177_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1128_ _2299_/Q _2011_/Q _1181_/S vssd1 vssd1 vccd1 vccd1 _1128_/X sky130_fd_sc_hd__mux2_1
XFILLER_53_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1059_ _2226_/Q _2230_/Q _2234_/Q _2238_/Q _1287_/S0 _1013_/B vssd1 vssd1 vccd1 vccd1
+ _1059_/X sky130_fd_sc_hd__mux4_2
Xoutput14 _1157_/Y vssd1 vssd1 vccd1 vccd1 r_val[1] sky130_fd_sc_hd__buf_4
XFILLER_48_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2100_ _2363_/CLK _2100_/D vssd1 vssd1 vccd1 vccd1 _2100_/Q sky130_fd_sc_hd__dfxtp_1
X_2031_ _2493_/CLK _2031_/D vssd1 vssd1 vccd1 vccd1 _2031_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1815_ _1940_/A0 _2361_/Q _1815_/S vssd1 vssd1 vccd1 vccd1 _2361_/D sky130_fd_sc_hd__mux2_1
X_1746_ _1806_/A _1906_/B vssd1 vssd1 vccd1 vccd1 _1750_/S sky130_fd_sc_hd__nor2_2
X_1677_ _2250_/Q _1982_/A1 _1680_/S vssd1 vssd1 vccd1 vccd1 _2250_/D sky130_fd_sc_hd__mux2_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2229_ _2229_/CLK _2229_/D vssd1 vssd1 vccd1 vccd1 _2229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1600_ _2189_/Q _1765_/A0 _1600_/S vssd1 vssd1 vccd1 vccd1 _2189_/D sky130_fd_sc_hd__mux2_1
X_1531_ _1641_/A _1531_/B vssd1 vssd1 vccd1 vccd1 _1535_/S sky130_fd_sc_hd__nor2_4
X_1462_ _1809_/A0 _2080_/Q _1463_/S vssd1 vssd1 vccd1 vccd1 _2080_/D sky130_fd_sc_hd__mux2_1
X_1393_ _1918_/A1 _2031_/Q _1395_/S vssd1 vssd1 vccd1 vccd1 _2031_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2014_ _2097_/CLK _2014_/D vssd1 vssd1 vccd1 vccd1 _2014_/Q sky130_fd_sc_hd__dfxtp_1
X_1729_ _2292_/Q _1739_/A0 _1730_/S vssd1 vssd1 vccd1 vccd1 _2292_/D sky130_fd_sc_hd__mux2_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1514_ _2120_/Q _1579_/A0 _1515_/S vssd1 vssd1 vccd1 vccd1 _2120_/D sky130_fd_sc_hd__mux2_1
X_2494_ _2495_/CLK _2494_/D vssd1 vssd1 vccd1 vccd1 _2494_/Q sky130_fd_sc_hd__dfxtp_1
X_1445_ _2067_/Q _1503_/A0 _1447_/S vssd1 vssd1 vccd1 vccd1 _2067_/D sky130_fd_sc_hd__mux2_1
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1376_ _1973_/A0 _2019_/Q _1378_/S vssd1 vssd1 vccd1 vccd1 _2019_/D sky130_fd_sc_hd__mux2_1
XFILLER_82_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout82 fanout85/X vssd1 vssd1 vccd1 vccd1 _1256_/S1 sky130_fd_sc_hd__buf_4
Xfanout71 _1023_/B vssd1 vssd1 vccd1 vccd1 _1244_/A1 sky130_fd_sc_hd__buf_4
Xfanout60 fanout68/X vssd1 vssd1 vccd1 vccd1 _1972_/A0 sky130_fd_sc_hd__buf_4
Xfanout93 fanout94/X vssd1 vssd1 vccd1 vccd1 _1100_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_6_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1230_ input7/X _1230_/B _1230_/C _1230_/D vssd1 vssd1 vccd1 vccd1 _1230_/X sky130_fd_sc_hd__or4_1
XFILLER_77_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1161_ _1220_/A _1161_/B vssd1 vssd1 vccd1 vccd1 _1161_/X sky130_fd_sc_hd__or2_1
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1092_ _2211_/Q _2215_/Q _2219_/Q _1995_/Q _1464_/A _1442_/B vssd1 vssd1 vccd1 vccd1
+ _1092_/X sky130_fd_sc_hd__mux4_1
XFILLER_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1994_ _2229_/CLK _1994_/D vssd1 vssd1 vccd1 vccd1 _1994_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2477_ _2477_/CLK _2477_/D vssd1 vssd1 vccd1 vccd1 _2477_/Q sky130_fd_sc_hd__dfxtp_1
X_1428_ _2055_/Q _1503_/A0 _1430_/S vssd1 vssd1 vccd1 vccd1 _2055_/D sky130_fd_sc_hd__mux2_1
XFILLER_18_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1359_ _2009_/Q _1505_/A0 _1359_/S vssd1 vssd1 vccd1 vccd1 _2009_/D sky130_fd_sc_hd__mux2_1
XFILLER_43_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2400_ _2482_/CLK _2400_/D vssd1 vssd1 vccd1 vccd1 _2400_/Q sky130_fd_sc_hd__dfxtp_1
X_2331_ _2335_/CLK _2331_/D vssd1 vssd1 vccd1 vccd1 _2331_/Q sky130_fd_sc_hd__dfxtp_1
X_2262_ _2302_/CLK _2262_/D vssd1 vssd1 vccd1 vccd1 _2262_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1213_ _1464_/C _1211_/X _1212_/X _1396_/C vssd1 vssd1 vccd1 vccd1 _1213_/X sky130_fd_sc_hd__o22a_1
XFILLER_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2193_ _2320_/CLK _2193_/D vssd1 vssd1 vccd1 vccd1 _2193_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1144_ _2403_/Q _2407_/Q _2411_/Q _2415_/Q _1256_/S0 _1256_/S1 vssd1 vssd1 vccd1
+ vccd1 _1145_/B sky130_fd_sc_hd__mux4_1
XFILLER_37_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1075_ _1065_/A _1073_/X _1074_/X vssd1 vssd1 vccd1 vccd1 _1075_/X sky130_fd_sc_hd__a21o_1
XFILLER_80_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1977_ _1977_/A0 _2490_/Q _1980_/S vssd1 vssd1 vccd1 vccd1 _2490_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1900_ _1905_/A0 _2429_/Q _1900_/S vssd1 vssd1 vccd1 vccd1 _2429_/D sky130_fd_sc_hd__mux2_1
X_1831_ _1911_/A _1886_/A vssd1 vssd1 vccd1 vccd1 _1835_/S sky130_fd_sc_hd__nor2_4
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1762_ _1762_/A0 _2318_/Q _1765_/S vssd1 vssd1 vccd1 vccd1 _2318_/D sky130_fd_sc_hd__mux2_1
X_1693_ _2263_/Q _1783_/A0 _1695_/S vssd1 vssd1 vccd1 vccd1 _2263_/D sky130_fd_sc_hd__mux2_1
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2314_ _2320_/CLK _2314_/D vssd1 vssd1 vccd1 vccd1 _2314_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2245_ _2301_/CLK _2245_/D vssd1 vssd1 vccd1 vccd1 _2245_/Q sky130_fd_sc_hd__dfxtp_1
X_2176_ _2176_/CLK _2176_/D vssd1 vssd1 vccd1 vccd1 _2176_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1127_ _2291_/Q _2295_/Q _1181_/S vssd1 vssd1 vccd1 vccd1 _1127_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1058_ _1453_/C _1056_/X _1057_/X _1464_/C vssd1 vssd1 vccd1 vccd1 _1058_/X sky130_fd_sc_hd__o22a_1
XFILLER_21_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput15 _1231_/X vssd1 vssd1 vccd1 vccd1 r_val[2] sky130_fd_sc_hd__buf_4
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_446 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2030_ _2493_/CLK _2030_/D vssd1 vssd1 vccd1 vccd1 _2030_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_42_clk clkbuf_leaf_4_clk/A vssd1 vssd1 vccd1 vccd1 _2159_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_30_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1814_ _1814_/A0 _2360_/Q _1815_/S vssd1 vssd1 vccd1 vccd1 _2360_/D sky130_fd_sc_hd__mux2_1
X_1745_ _1845_/A1 _2305_/Q _1745_/S vssd1 vssd1 vccd1 vccd1 _2305_/D sky130_fd_sc_hd__mux2_1
XFILLER_7_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1676_ _1726_/A _1916_/B vssd1 vssd1 vccd1 vccd1 _1680_/S sky130_fd_sc_hd__nor2_4
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2228_ _2229_/CLK _2228_/D vssd1 vssd1 vccd1 vccd1 _2228_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2159_ _2159_/CLK _2159_/D vssd1 vssd1 vccd1 vccd1 _2159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_446 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_33_clk clkbuf_2_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _2421_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_42_47 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_24_clk clkbuf_2_3__f_clk/X vssd1 vssd1 vccd1 vccd1 _2261_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_80_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1530_ _2133_/Q _1585_/A0 _1530_/S vssd1 vssd1 vccd1 vccd1 _2133_/D sky130_fd_sc_hd__mux2_1
X_1461_ _1778_/A0 _2079_/Q _1463_/S vssd1 vssd1 vccd1 vccd1 _2079_/D sky130_fd_sc_hd__mux2_1
X_1392_ _1977_/A0 _2030_/Q _1395_/S vssd1 vssd1 vccd1 vccd1 _2030_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2013_ _2301_/CLK _2013_/D vssd1 vssd1 vccd1 vccd1 _2013_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_15_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _2369_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1728_ _2291_/Q _1738_/A0 _1730_/S vssd1 vssd1 vccd1 vccd1 _2291_/D sky130_fd_sc_hd__mux2_1
X_1659_ _1664_/A0 _2236_/Q _1660_/S vssd1 vssd1 vccd1 vccd1 _2236_/D sky130_fd_sc_hd__mux2_1
XFILLER_85_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1513_ _2119_/Q _1583_/A0 _1515_/S vssd1 vssd1 vccd1 vccd1 _2119_/D sky130_fd_sc_hd__mux2_1
X_2493_ _2493_/CLK _2493_/D vssd1 vssd1 vccd1 vccd1 _2493_/Q sky130_fd_sc_hd__dfxtp_1
X_1444_ _2066_/Q _1822_/A0 _1447_/S vssd1 vssd1 vccd1 vccd1 _2066_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_4_clk clkbuf_leaf_4_clk/A vssd1 vssd1 vccd1 vccd1 _2461_/CLK sky130_fd_sc_hd__clkbuf_16
X_1375_ _1972_/A0 _2018_/Q _1378_/S vssd1 vssd1 vccd1 vccd1 _2018_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout83 fanout85/X vssd1 vssd1 vccd1 vccd1 _1464_/B sky130_fd_sc_hd__clkbuf_8
Xfanout61 fanout68/X vssd1 vssd1 vccd1 vccd1 _1962_/A0 sky130_fd_sc_hd__clkbuf_2
Xfanout50 _1843_/A1 vssd1 vssd1 vccd1 vccd1 _1793_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout72 input4/X vssd1 vssd1 vccd1 vccd1 _1023_/B sky130_fd_sc_hd__buf_6
XFILLER_6_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout94 input2/X vssd1 vssd1 vccd1 vccd1 fanout94/X sky130_fd_sc_hd__buf_4
XFILLER_6_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1160_ _2404_/Q _2408_/Q _2412_/Q _2416_/Q _1181_/S _0992_/A vssd1 vssd1 vccd1 vccd1
+ _1161_/B sky130_fd_sc_hd__mux4_1
XFILLER_77_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1091_ _2195_/Q _2199_/Q _2203_/Q _2207_/Q _1453_/A _1285_/S1 vssd1 vssd1 vccd1 vccd1
+ _1091_/X sky130_fd_sc_hd__mux4_1
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1993_ _2337_/CLK _1993_/D vssd1 vssd1 vccd1 vccd1 _1993_/Q sky130_fd_sc_hd__dfxtp_1
X_2476_ _2480_/CLK _2476_/D vssd1 vssd1 vccd1 vccd1 _2476_/Q sky130_fd_sc_hd__dfxtp_1
X_1427_ _2054_/Q _1762_/A0 _1430_/S vssd1 vssd1 vccd1 vccd1 _2054_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1358_ _2008_/Q _1824_/A0 _1359_/S vssd1 vssd1 vccd1 vccd1 _2008_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1289_ _1420_/C _1285_/X _1288_/X _1284_/X vssd1 vssd1 vccd1 vccd1 _1307_/B sky130_fd_sc_hd__o211a_1
XFILLER_70_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2330_ _2337_/CLK _2330_/D vssd1 vssd1 vccd1 vccd1 _2330_/Q sky130_fd_sc_hd__dfxtp_1
X_2261_ _2261_/CLK _2261_/D vssd1 vssd1 vccd1 vccd1 _2261_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1212_ _2228_/Q _2232_/Q _2236_/Q _2240_/Q _1287_/S0 _1013_/B vssd1 vssd1 vccd1 vccd1
+ _1212_/X sky130_fd_sc_hd__mux4_1
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2192_ _2320_/CLK _2192_/D vssd1 vssd1 vccd1 vccd1 _2192_/Q sky130_fd_sc_hd__dfxtp_1
X_1143_ _1298_/B2 _1140_/X _1142_/X _1295_/B2 vssd1 vssd1 vccd1 vccd1 _1143_/X sky130_fd_sc_hd__a22o_1
X_1074_ _1234_/A1 _1072_/X _1241_/B1 vssd1 vssd1 vccd1 vccd1 _1074_/X sky130_fd_sc_hd__a21o_1
XFILLER_52_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1976_ _1976_/A _1976_/B vssd1 vssd1 vccd1 vccd1 _1980_/S sky130_fd_sc_hd__nand2_2
XFILLER_60_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2459_ _2461_/CLK _2459_/D vssd1 vssd1 vccd1 vccd1 _2459_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1830_ _2373_/Q _1975_/A0 _1830_/S vssd1 vssd1 vccd1 vccd1 _2373_/D sky130_fd_sc_hd__mux2_1
X_1761_ _1821_/A _1921_/A vssd1 vssd1 vccd1 vccd1 _1765_/S sky130_fd_sc_hd__nand2_4
X_1692_ _2262_/Q _1742_/A0 _1695_/S vssd1 vssd1 vccd1 vccd1 _2262_/D sky130_fd_sc_hd__mux2_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2313_ _2363_/CLK _2313_/D vssd1 vssd1 vccd1 vccd1 _2313_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2244_ _2481_/CLK _2244_/D vssd1 vssd1 vccd1 vccd1 _2244_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2175_ _2177_/CLK _2175_/D vssd1 vssd1 vccd1 vccd1 _2175_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1126_ _2275_/Q _2279_/Q _2283_/Q _2287_/Q _1181_/S _0992_/A vssd1 vssd1 vccd1 vccd1
+ _1126_/X sky130_fd_sc_hd__mux4_1
XFILLER_38_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1057_ _2210_/Q _2214_/Q _2218_/Q _1994_/Q _1464_/A _1442_/B vssd1 vssd1 vccd1 vccd1
+ _1057_/X sky130_fd_sc_hd__mux4_1
X_1959_ _1964_/A0 _2476_/Q _1960_/S vssd1 vssd1 vccd1 vccd1 _2476_/D sky130_fd_sc_hd__mux2_1
Xoutput16 _1308_/X vssd1 vssd1 vccd1 vccd1 r_val[3] sky130_fd_sc_hd__buf_4
XFILLER_0_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clkbuf_0_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1813_ _1823_/A0 _2359_/Q _1815_/S vssd1 vssd1 vccd1 vccd1 _2359_/D sky130_fd_sc_hd__mux2_1
X_1744_ _1984_/A1 _2304_/Q _1745_/S vssd1 vssd1 vccd1 vccd1 _2304_/D sky130_fd_sc_hd__mux2_1
X_1675_ _2249_/Q _1935_/A0 _1675_/S vssd1 vssd1 vccd1 vccd1 _2249_/D sky130_fd_sc_hd__mux2_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2227_ _2240_/CLK _2227_/D vssd1 vssd1 vccd1 vccd1 _2227_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2158_ _2159_/CLK _2158_/D vssd1 vssd1 vccd1 vccd1 _2158_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1109_ _1174_/A _1107_/X _1108_/X vssd1 vssd1 vccd1 vccd1 _1109_/Y sky130_fd_sc_hd__a21oi_1
X_2089_ _2097_/CLK _2089_/D vssd1 vssd1 vccd1 vccd1 _2089_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1460_ _1777_/A0 _2078_/Q _1463_/S vssd1 vssd1 vccd1 vccd1 _2078_/D sky130_fd_sc_hd__mux2_1
X_1391_ _1901_/A _1976_/A vssd1 vssd1 vccd1 vccd1 _1395_/S sky130_fd_sc_hd__nand2_2
XFILLER_82_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2012_ _2481_/CLK _2012_/D vssd1 vssd1 vccd1 vccd1 _2012_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1727_ _2290_/Q _1732_/A0 _1730_/S vssd1 vssd1 vccd1 vccd1 _2290_/D sky130_fd_sc_hd__mux2_1
X_1658_ _1663_/A0 _2235_/Q _1660_/S vssd1 vssd1 vccd1 vccd1 _2235_/D sky130_fd_sc_hd__mux2_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1589_ _2180_/Q _1814_/A0 _1590_/S vssd1 vssd1 vccd1 vccd1 _2180_/D sky130_fd_sc_hd__mux2_1
XFILLER_58_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2492_ _2493_/CLK _2492_/D vssd1 vssd1 vccd1 vccd1 _2492_/Q sky130_fd_sc_hd__dfxtp_1
X_1512_ _2118_/Q _1582_/A0 _1515_/S vssd1 vssd1 vccd1 vccd1 _2118_/D sky130_fd_sc_hd__mux2_1
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1443_ _1486_/A _1926_/B vssd1 vssd1 vccd1 vccd1 _1447_/S sky130_fd_sc_hd__nor2_2
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1374_ _1921_/A _1901_/B vssd1 vssd1 vccd1 vccd1 _1378_/S sky130_fd_sc_hd__nand2_2
XFILLER_67_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout40 fanout44/X vssd1 vssd1 vccd1 vccd1 _1973_/A0 sky130_fd_sc_hd__buf_4
Xfanout51 _1843_/A1 vssd1 vssd1 vccd1 vccd1 _1783_/A0 sky130_fd_sc_hd__buf_4
Xfanout73 _1180_/A vssd1 vssd1 vccd1 vccd1 _1220_/A sky130_fd_sc_hd__buf_8
Xfanout62 fanout68/X vssd1 vssd1 vccd1 vccd1 _1902_/A0 sky130_fd_sc_hd__clkbuf_4
Xfanout95 _1660_/A0 vssd1 vssd1 vccd1 vccd1 _1585_/A0 sky130_fd_sc_hd__clkbuf_4
Xfanout84 fanout85/X vssd1 vssd1 vccd1 vccd1 _0992_/A sky130_fd_sc_hd__buf_4
XFILLER_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1090_ _1087_/X _1088_/X _1086_/X _1089_/X _1258_/A _1024_/B vssd1 vssd1 vccd1 vccd1
+ _1090_/X sky130_fd_sc_hd__mux4_2
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1992_ _2457_/CLK _1992_/D vssd1 vssd1 vccd1 vccd1 _1992_/Q sky130_fd_sc_hd__dfxtp_1
X_2475_ _2479_/CLK _2475_/D vssd1 vssd1 vccd1 vccd1 _2475_/Q sky130_fd_sc_hd__dfxtp_1
X_1426_ _1911_/A _1486_/A vssd1 vssd1 vccd1 vccd1 _1430_/S sky130_fd_sc_hd__nor2_4
X_1357_ _2007_/Q _1503_/A0 _1359_/S vssd1 vssd1 vccd1 vccd1 _2007_/D sky130_fd_sc_hd__mux2_1
XFILLER_28_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1288_ _1464_/C _1286_/X _1287_/X _1396_/C vssd1 vssd1 vccd1 vccd1 _1288_/X sky130_fd_sc_hd__o22a_1
XFILLER_24_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2260_ _2301_/CLK _2260_/D vssd1 vssd1 vccd1 vccd1 _2260_/Q sky130_fd_sc_hd__dfxtp_1
X_1211_ _2212_/Q _2216_/Q _2220_/Q _1996_/Q _1287_/S0 _1442_/B vssd1 vssd1 vccd1 vccd1
+ _1211_/X sky130_fd_sc_hd__mux4_1
X_2191_ _2241_/CLK _2191_/D vssd1 vssd1 vccd1 vccd1 _2191_/Q sky130_fd_sc_hd__dfxtp_1
X_1142_ _2371_/Q _2375_/Q _2379_/Q _2019_/Q _1253_/S0 _1253_/S1 vssd1 vssd1 vccd1
+ vccd1 _1142_/X sky130_fd_sc_hd__mux4_2
XFILLER_18_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1073_ _2042_/Q _2046_/Q _1277_/S vssd1 vssd1 vccd1 vccd1 _1073_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1975_ _1975_/A0 _2489_/Q _1975_/S vssd1 vssd1 vccd1 vccd1 _2489_/D sky130_fd_sc_hd__mux2_1
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2458_ _2461_/CLK _2458_/D vssd1 vssd1 vccd1 vccd1 _2458_/Q sky130_fd_sc_hd__dfxtp_1
X_1409_ _1245_/S0 _1409_/B _1409_/C vssd1 vssd1 vccd1 vccd1 _1976_/B sky130_fd_sc_hd__and3b_4
X_2389_ _2433_/CLK _2389_/D vssd1 vssd1 vccd1 vccd1 _2389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1760_ _2317_/Q _1765_/A0 _1760_/S vssd1 vssd1 vccd1 vccd1 _2317_/D sky130_fd_sc_hd__mux2_1
X_1691_ _1691_/A _1936_/B vssd1 vssd1 vccd1 vccd1 _1695_/S sky130_fd_sc_hd__nor2_2
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2312_ _2320_/CLK _2312_/D vssd1 vssd1 vccd1 vccd1 _2312_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2243_ _2301_/CLK _2243_/D vssd1 vssd1 vccd1 vccd1 _2243_/Q sky130_fd_sc_hd__dfxtp_1
X_2174_ _2177_/CLK _2174_/D vssd1 vssd1 vccd1 vccd1 _2174_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1125_ _1237_/A _1125_/B vssd1 vssd1 vccd1 vccd1 _1125_/Y sky130_fd_sc_hd__nor2_1
X_1056_ _2194_/Q _2198_/Q _2202_/Q _2206_/Q _1464_/A _1013_/B vssd1 vssd1 vccd1 vccd1
+ _1056_/X sky130_fd_sc_hd__mux4_1
XFILLER_80_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1958_ _1963_/A0 _2475_/Q _1960_/S vssd1 vssd1 vccd1 vccd1 _2475_/D sky130_fd_sc_hd__mux2_1
X_1889_ _1904_/A0 _2420_/Q _1890_/S vssd1 vssd1 vccd1 vccd1 _2420_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1812_ _1822_/A0 _2358_/Q _1815_/S vssd1 vssd1 vccd1 vccd1 _2358_/D sky130_fd_sc_hd__mux2_1
X_1743_ _1843_/A1 _2303_/Q _1745_/S vssd1 vssd1 vccd1 vccd1 _2303_/D sky130_fd_sc_hd__mux2_1
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1674_ _2248_/Q _1804_/A0 _1675_/S vssd1 vssd1 vccd1 vccd1 _2248_/D sky130_fd_sc_hd__mux2_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2226_ _2240_/CLK _2226_/D vssd1 vssd1 vccd1 vccd1 _2226_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2157_ _2449_/CLK _2157_/D vssd1 vssd1 vccd1 vccd1 _2157_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1108_ _1234_/A1 _1106_/X _1241_/B1 vssd1 vssd1 vccd1 vccd1 _1108_/X sky130_fd_sc_hd__a21o_1
X_2088_ _2097_/CLK _2088_/D vssd1 vssd1 vccd1 vccd1 _2088_/Q sky130_fd_sc_hd__dfxtp_1
X_1039_ _1033_/X _1036_/X _1037_/X vssd1 vssd1 vccd1 vccd1 _1048_/C sky130_fd_sc_hd__o21a_1
XFILLER_53_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_50 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1390_ _1935_/A0 _2029_/Q _1390_/S vssd1 vssd1 vccd1 vccd1 _2029_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2011_ _2296_/CLK _2011_/D vssd1 vssd1 vccd1 vccd1 _2011_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1726_ _1726_/A _1966_/B vssd1 vssd1 vccd1 vccd1 _1730_/S sky130_fd_sc_hd__nor2_2
X_1657_ _1662_/A0 _2234_/Q _1660_/S vssd1 vssd1 vccd1 vccd1 _2234_/D sky130_fd_sc_hd__mux2_1
X_1588_ _2179_/Q _1663_/A0 _1590_/S vssd1 vssd1 vccd1 vccd1 _2179_/D sky130_fd_sc_hd__mux2_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2209_ _2368_/CLK _2209_/D vssd1 vssd1 vccd1 vccd1 _2209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_2_0__f_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_4_clk/A sky130_fd_sc_hd__clkbuf_16
XFILLER_60_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2491_ _2493_/CLK _2491_/D vssd1 vssd1 vccd1 vccd1 _2491_/Q sky130_fd_sc_hd__dfxtp_1
X_1511_ _1911_/A _1566_/A vssd1 vssd1 vccd1 vccd1 _1515_/S sky130_fd_sc_hd__nor2_2
X_1442_ _1464_/A _1442_/B _1453_/C vssd1 vssd1 vccd1 vccd1 _1926_/B sky130_fd_sc_hd__or3_4
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1373_ _1373_/A _1385_/B vssd1 vssd1 vccd1 vccd1 _1886_/A sky130_fd_sc_hd__or2_4
XFILLER_23_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1709_ _2276_/Q _1904_/A0 _1710_/S vssd1 vssd1 vccd1 vccd1 _2276_/D sky130_fd_sc_hd__mux2_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout30 _1011_/X vssd1 vssd1 vccd1 vccd1 _1302_/A1 sky130_fd_sc_hd__buf_2
XFILLER_80_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout41 fanout44/X vssd1 vssd1 vccd1 vccd1 _1903_/A0 sky130_fd_sc_hd__clkbuf_4
Xfanout63 fanout68/X vssd1 vssd1 vccd1 vccd1 _1732_/A0 sky130_fd_sc_hd__buf_2
Xfanout74 _1274_/A vssd1 vssd1 vccd1 vccd1 _1237_/A sky130_fd_sc_hd__buf_4
Xfanout52 input9/X vssd1 vssd1 vccd1 vccd1 _1843_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout85 input2/X vssd1 vssd1 vccd1 vccd1 fanout85/X sky130_fd_sc_hd__buf_8
Xfanout96 _1660_/A0 vssd1 vssd1 vccd1 vccd1 _1980_/A0 sky130_fd_sc_hd__clkbuf_4
XFILLER_6_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1991_ _2329_/CLK _1991_/D vssd1 vssd1 vccd1 vccd1 _1991_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2474_ _2479_/CLK _2474_/D vssd1 vssd1 vccd1 vccd1 _2474_/Q sky130_fd_sc_hd__dfxtp_1
X_1425_ _2053_/Q _1505_/A0 _1425_/S vssd1 vssd1 vccd1 vccd1 _2053_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1356_ _2006_/Q _1762_/A0 _1359_/S vssd1 vssd1 vccd1 vccd1 _2006_/D sky130_fd_sc_hd__mux2_1
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1287_ _2229_/Q _2233_/Q _2237_/Q _2241_/Q _1287_/S0 _1013_/B vssd1 vssd1 vccd1 vccd1
+ _1287_/X sky130_fd_sc_hd__mux4_1
XFILLER_36_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2190_ _2240_/CLK _2190_/D vssd1 vssd1 vccd1 vccd1 _2190_/Q sky130_fd_sc_hd__dfxtp_1
X_1210_ _2180_/Q _2000_/Q _2188_/Q _2192_/Q _1285_/S0 _1285_/S1 vssd1 vssd1 vccd1
+ vccd1 _1210_/X sky130_fd_sc_hd__mux4_2
X_1141_ _2419_/Q _2023_/Q _2427_/Q _2431_/Q _1256_/S0 _1256_/S1 vssd1 vssd1 vccd1
+ vccd1 _1146_/B sky130_fd_sc_hd__mux4_1
XFILLER_65_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1072_ _2034_/Q _2038_/Q _1277_/S vssd1 vssd1 vccd1 vccd1 _1072_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1974_ _1974_/A0 _2488_/Q _1975_/S vssd1 vssd1 vccd1 vccd1 _2488_/D sky130_fd_sc_hd__mux2_1
X_2457_ _2457_/CLK _2457_/D vssd1 vssd1 vccd1 vccd1 _2457_/Q sky130_fd_sc_hd__dfxtp_1
X_1408_ _1845_/A1 _2041_/Q _1408_/S vssd1 vssd1 vccd1 vccd1 _2041_/D sky130_fd_sc_hd__mux2_1
X_2388_ _2433_/CLK _2388_/D vssd1 vssd1 vccd1 vccd1 _2388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1339_ _1998_/Q _1662_/A0 _1342_/S vssd1 vssd1 vccd1 vccd1 _1998_/D sky130_fd_sc_hd__mux2_1
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1690_ _2261_/Q _1935_/A0 _1690_/S vssd1 vssd1 vccd1 vccd1 _2261_/D sky130_fd_sc_hd__mux2_1
X_2311_ _2363_/CLK _2311_/D vssd1 vssd1 vccd1 vccd1 _2311_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2242_ _2343_/CLK _2242_/D vssd1 vssd1 vccd1 vccd1 _2242_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2173_ _2177_/CLK _2173_/D vssd1 vssd1 vccd1 vccd1 _2173_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1124_ _2243_/Q _2247_/Q _2251_/Q _2255_/Q _1245_/S0 _1174_/A vssd1 vssd1 vccd1 vccd1
+ _1125_/B sky130_fd_sc_hd__mux4_1
X_1055_ _1295_/B2 _1049_/X _1054_/X _1298_/B2 vssd1 vssd1 vccd1 vccd1 _1055_/X sky130_fd_sc_hd__a22o_1
XFILLER_53_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1957_ _1962_/A0 _2474_/Q _1960_/S vssd1 vssd1 vccd1 vccd1 _2474_/D sky130_fd_sc_hd__mux2_1
X_1888_ _1903_/A0 _2419_/Q _1890_/S vssd1 vssd1 vccd1 vccd1 _2419_/D sky130_fd_sc_hd__mux2_1
XFILLER_29_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_36_clk clkbuf_2_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _2482_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_71_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_27_clk clkbuf_2_3__f_clk/X vssd1 vssd1 vccd1 vccd1 _2343_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1811_ _1821_/A _1971_/A vssd1 vssd1 vccd1 vccd1 _1815_/S sky130_fd_sc_hd__nand2_2
X_1742_ _1742_/A0 _2302_/Q _1745_/S vssd1 vssd1 vccd1 vccd1 _2302_/D sky130_fd_sc_hd__mux2_1
XFILLER_11_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1673_ _2247_/Q _1793_/A1 _1675_/S vssd1 vssd1 vccd1 vccd1 _2247_/D sky130_fd_sc_hd__mux2_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2225_ _2302_/CLK _2225_/D vssd1 vssd1 vccd1 vccd1 _2225_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2156_ _2176_/CLK _2156_/D vssd1 vssd1 vccd1 vccd1 _2156_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2087_ _2335_/CLK _2087_/D vssd1 vssd1 vccd1 vccd1 _2087_/Q sky130_fd_sc_hd__dfxtp_1
X_1107_ _2043_/Q _2047_/Q _1233_/S vssd1 vssd1 vccd1 vccd1 _1107_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_18_clk clkbuf_2_3__f_clk/X vssd1 vssd1 vccd1 vccd1 _2497_/CLK sky130_fd_sc_hd__clkbuf_16
X_1038_ _1040_/B input6/X vssd1 vssd1 vccd1 vccd1 _1373_/A sky130_fd_sc_hd__nand2b_4
XFILLER_34_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2010_ _2301_/CLK _2010_/D vssd1 vssd1 vccd1 vccd1 _2010_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1725_ _1960_/A0 _2289_/Q _1725_/S vssd1 vssd1 vccd1 vccd1 _2289_/D sky130_fd_sc_hd__mux2_1
X_1656_ _1661_/A _1976_/B vssd1 vssd1 vccd1 vccd1 _1660_/S sky130_fd_sc_hd__nand2_2
Xclkbuf_leaf_7_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _2363_/CLK sky130_fd_sc_hd__clkbuf_16
X_1587_ _2178_/Q _1662_/A0 _1590_/S vssd1 vssd1 vccd1 vccd1 _2178_/D sky130_fd_sc_hd__mux2_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2208_ _2368_/CLK _2208_/D vssd1 vssd1 vccd1 vccd1 _2208_/Q sky130_fd_sc_hd__dfxtp_1
X_2139_ _2177_/CLK _2139_/D vssd1 vssd1 vccd1 vccd1 _2139_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2490_ _2493_/CLK _2490_/D vssd1 vssd1 vccd1 vccd1 _2490_/Q sky130_fd_sc_hd__dfxtp_1
X_1510_ _2117_/Q _1980_/A0 _1510_/S vssd1 vssd1 vccd1 vccd1 _2117_/D sky130_fd_sc_hd__mux2_1
X_1441_ _2065_/Q _1985_/A1 _1441_/S vssd1 vssd1 vccd1 vccd1 _2065_/D sky130_fd_sc_hd__mux2_1
XFILLER_4_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1372_ _1373_/A _1385_/B vssd1 vssd1 vccd1 vccd1 _1901_/B sky130_fd_sc_hd__nor2_8
XFILLER_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1708_ _2275_/Q _1963_/A0 _1710_/S vssd1 vssd1 vccd1 vccd1 _2275_/D sky130_fd_sc_hd__mux2_1
X_1639_ _1664_/A0 _2220_/Q _1640_/S vssd1 vssd1 vccd1 vccd1 _2220_/D sky130_fd_sc_hd__mux2_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout31 _1020_/A vssd1 vssd1 vccd1 vccd1 _1241_/B1 sky130_fd_sc_hd__clkbuf_8
Xfanout20 _1666_/A vssd1 vssd1 vccd1 vccd1 _1726_/A sky130_fd_sc_hd__buf_12
Xfanout53 _1662_/A0 vssd1 vssd1 vccd1 vccd1 _1582_/A0 sky130_fd_sc_hd__clkbuf_4
Xfanout42 fanout44/X vssd1 vssd1 vccd1 vccd1 _1963_/A0 sky130_fd_sc_hd__buf_4
Xfanout64 _1742_/A0 vssd1 vssd1 vccd1 vccd1 _1982_/A1 sky130_fd_sc_hd__buf_4
XFILLER_10_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout97 _1965_/A0 vssd1 vssd1 vccd1 vccd1 _1660_/A0 sky130_fd_sc_hd__buf_4
Xfanout86 _1283_/S1 vssd1 vssd1 vccd1 vccd1 _1285_/S1 sky130_fd_sc_hd__buf_6
Xfanout75 _1180_/A vssd1 vssd1 vccd1 vccd1 _1274_/A sky130_fd_sc_hd__buf_6
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1990_ _2457_/CLK _1990_/D vssd1 vssd1 vccd1 vccd1 _1990_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2473_ _2481_/CLK _2473_/D vssd1 vssd1 vccd1 vccd1 _2473_/Q sky130_fd_sc_hd__dfxtp_1
X_1424_ _2052_/Q _1824_/A0 _1425_/S vssd1 vssd1 vccd1 vccd1 _2052_/D sky130_fd_sc_hd__mux2_1
X_1355_ _1681_/B _1486_/A vssd1 vssd1 vccd1 vccd1 _1359_/S sky130_fd_sc_hd__nor2_4
XFILLER_55_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1286_ _2213_/Q _2217_/Q _2221_/Q _1997_/Q _1287_/S0 _1442_/B vssd1 vssd1 vccd1 vccd1
+ _1286_/X sky130_fd_sc_hd__mux4_1
XFILLER_24_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_447 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1140_ _2387_/Q _2391_/Q _2395_/Q _2399_/Q _1253_/S0 _1256_/S1 vssd1 vssd1 vccd1
+ vccd1 _1140_/X sky130_fd_sc_hd__mux4_1
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1071_ _1237_/A _1071_/B vssd1 vssd1 vccd1 vccd1 _1071_/X sky130_fd_sc_hd__or2_1
XFILLER_45_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1973_ _1973_/A0 _2487_/Q _1975_/S vssd1 vssd1 vccd1 vccd1 _2487_/D sky130_fd_sc_hd__mux2_1
XFILLER_60_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2456_ _2479_/CLK _2456_/D vssd1 vssd1 vccd1 vccd1 _2456_/Q sky130_fd_sc_hd__dfxtp_1
X_1407_ _1984_/A1 _2040_/Q _1408_/S vssd1 vssd1 vccd1 vccd1 _2040_/D sky130_fd_sc_hd__mux2_1
X_2387_ _2433_/CLK _2387_/D vssd1 vssd1 vccd1 vccd1 _2387_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1338_ _1646_/A _1911_/A vssd1 vssd1 vccd1 vccd1 _1342_/S sky130_fd_sc_hd__nor2_4
XFILLER_68_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1269_ _2265_/Q _2305_/Q _1270_/S vssd1 vssd1 vccd1 vccd1 _1269_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2310_ _2320_/CLK _2310_/D vssd1 vssd1 vccd1 vccd1 _2310_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2241_ _2241_/CLK _2241_/D vssd1 vssd1 vccd1 vccd1 _2241_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2172_ _2176_/CLK _2172_/D vssd1 vssd1 vccd1 vccd1 _2172_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1123_ _1174_/A _1120_/X _1122_/X vssd1 vssd1 vccd1 vccd1 _1123_/Y sky130_fd_sc_hd__a21oi_1
X_1054_ _2130_/Q _2134_/Q _2138_/Q _2002_/Q _1287_/S0 _1013_/B vssd1 vssd1 vccd1 vccd1
+ _1054_/X sky130_fd_sc_hd__mux4_1
XFILLER_65_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1956_ _1966_/A _1956_/B vssd1 vssd1 vccd1 vccd1 _1960_/S sky130_fd_sc_hd__or2_4
X_1887_ _1902_/A0 _2418_/Q _1890_/S vssd1 vssd1 vccd1 vccd1 _2418_/D sky130_fd_sc_hd__mux2_1
X_2439_ _2448_/CLK _2439_/D vssd1 vssd1 vccd1 vccd1 _2439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1810_ _1940_/A0 _2357_/Q _1810_/S vssd1 vssd1 vccd1 vccd1 _2357_/D sky130_fd_sc_hd__mux2_1
XFILLER_70_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1741_ _1861_/A _1941_/B vssd1 vssd1 vccd1 vccd1 _1745_/S sky130_fd_sc_hd__nand2_4
X_1672_ _2246_/Q _1982_/A1 _1675_/S vssd1 vssd1 vccd1 vccd1 _2246_/D sky130_fd_sc_hd__mux2_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2224_ _2302_/CLK _2224_/D vssd1 vssd1 vccd1 vccd1 _2224_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2155_ _2159_/CLK _2155_/D vssd1 vssd1 vccd1 vccd1 _2155_/Q sky130_fd_sc_hd__dfxtp_1
X_1106_ _2035_/Q _2039_/Q _1277_/S vssd1 vssd1 vccd1 vccd1 _1106_/X sky130_fd_sc_hd__mux2_1
X_2086_ _2094_/CLK _2086_/D vssd1 vssd1 vccd1 vccd1 _2086_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1037_ _1040_/B input6/X vssd1 vssd1 vccd1 vccd1 _1037_/X sky130_fd_sc_hd__and2b_4
XFILLER_53_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1939_ _1979_/A0 _2460_/Q _1940_/S vssd1 vssd1 vccd1 vccd1 _2460_/D sky130_fd_sc_hd__mux2_1
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1724_ _1904_/A0 _2288_/Q _1725_/S vssd1 vssd1 vccd1 vccd1 _2288_/D sky130_fd_sc_hd__mux2_1
XFILLER_7_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1655_ _1660_/A0 _2233_/Q _1655_/S vssd1 vssd1 vccd1 vccd1 _2233_/D sky130_fd_sc_hd__mux2_1
X_1586_ _1646_/A _1906_/B vssd1 vssd1 vccd1 vccd1 _1590_/S sky130_fd_sc_hd__nor2_2
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2207_ _2461_/CLK _2207_/D vssd1 vssd1 vccd1 vccd1 _2207_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2138_ _2232_/CLK _2138_/D vssd1 vssd1 vccd1 vccd1 _2138_/Q sky130_fd_sc_hd__dfxtp_1
X_2069_ _2337_/CLK _2069_/D vssd1 vssd1 vccd1 vccd1 _2069_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1440_ _2064_/Q _1984_/A1 _1441_/S vssd1 vssd1 vccd1 vccd1 _2064_/D sky130_fd_sc_hd__mux2_1
XFILLER_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1371_ _1505_/A0 _2017_/Q _1371_/S vssd1 vssd1 vccd1 vccd1 _2017_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1707_ _2274_/Q _1732_/A0 _1710_/S vssd1 vssd1 vccd1 vccd1 _2274_/D sky130_fd_sc_hd__mux2_1
X_1638_ _1978_/A0 _2219_/Q _1640_/S vssd1 vssd1 vccd1 vccd1 _2219_/D sky130_fd_sc_hd__mux2_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1569_ _2164_/Q _1579_/A0 _1570_/S vssd1 vssd1 vccd1 vccd1 _2164_/D sky130_fd_sc_hd__mux2_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout21 _1322_/A vssd1 vssd1 vccd1 vccd1 _1354_/A sky130_fd_sc_hd__buf_6
XFILLER_80_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout54 input8/X vssd1 vssd1 vccd1 vccd1 _1662_/A0 sky130_fd_sc_hd__clkbuf_4
Xfanout43 fanout44/X vssd1 vssd1 vccd1 vccd1 _1738_/A0 sky130_fd_sc_hd__clkbuf_2
Xfanout32 _1258_/A vssd1 vssd1 vccd1 vccd1 _1020_/A sky130_fd_sc_hd__buf_4
Xfanout65 _1742_/A0 vssd1 vssd1 vccd1 vccd1 _1842_/A1 sky130_fd_sc_hd__clkbuf_2
Xfanout76 input3/X vssd1 vssd1 vccd1 vccd1 _1180_/A sky130_fd_sc_hd__buf_6
XFILLER_22_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout98 _1960_/A0 vssd1 vssd1 vccd1 vccd1 _1975_/A0 sky130_fd_sc_hd__clkbuf_4
Xfanout87 _1283_/S1 vssd1 vssd1 vccd1 vccd1 _1304_/S1 sky130_fd_sc_hd__buf_6
XFILLER_10_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2472_ _2481_/CLK _2472_/D vssd1 vssd1 vccd1 vccd1 _2472_/Q sky130_fd_sc_hd__dfxtp_1
X_1423_ _2051_/Q _1503_/A0 _1425_/S vssd1 vssd1 vccd1 vccd1 _2051_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1354_ _1354_/A _1398_/B vssd1 vssd1 vccd1 vccd1 _1470_/B sky130_fd_sc_hd__or2_4
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1285_ _2181_/Q _2001_/Q _2189_/Q _2193_/Q _1285_/S0 _1285_/S1 vssd1 vssd1 vccd1
+ vccd1 _1285_/X sky130_fd_sc_hd__mux4_1
XFILLER_68_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1070_ _2342_/Q _2494_/Q _2422_/Q _2462_/Q _1245_/S0 _1409_/B vssd1 vssd1 vccd1 vccd1
+ _1071_/B sky130_fd_sc_hd__mux4_1
XFILLER_80_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1972_ _1972_/A0 _2486_/Q _1975_/S vssd1 vssd1 vccd1 vccd1 _2486_/D sky130_fd_sc_hd__mux2_1
XFILLER_33_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2455_ _2480_/CLK _2455_/D vssd1 vssd1 vccd1 vccd1 _2455_/Q sky130_fd_sc_hd__dfxtp_1
X_2386_ _2433_/CLK _2386_/D vssd1 vssd1 vccd1 vccd1 _2386_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1406_ _1983_/A1 _2039_/Q _1408_/S vssd1 vssd1 vccd1 vccd1 _2039_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1337_ _1366_/A _1420_/C vssd1 vssd1 vccd1 vccd1 _1911_/A sky130_fd_sc_hd__or2_4
XFILLER_68_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1268_ _1398_/A _1244_/X _1267_/Y _1354_/A _1260_/Y vssd1 vssd1 vccd1 vccd1 _1268_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_64_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1199_ _1237_/A _1199_/B vssd1 vssd1 vccd1 vccd1 _1199_/Y sky130_fd_sc_hd__nor2_1
XFILLER_36_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2240_ _2240_/CLK _2240_/D vssd1 vssd1 vccd1 vccd1 _2240_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2171_ _2177_/CLK _2171_/D vssd1 vssd1 vccd1 vccd1 _2171_/Q sky130_fd_sc_hd__dfxtp_1
X_1122_ _1234_/A1 _1121_/X _1241_/B1 vssd1 vssd1 vccd1 vccd1 _1122_/X sky130_fd_sc_hd__a21o_1
X_1053_ _1258_/A _1050_/X _1052_/X _1024_/B vssd1 vssd1 vccd1 vccd1 _1053_/X sky130_fd_sc_hd__o211a_1
XFILLER_53_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1955_ _1960_/A0 _2473_/Q _1955_/S vssd1 vssd1 vccd1 vccd1 _2473_/D sky130_fd_sc_hd__mux2_1
X_1886_ _1886_/A _1966_/B vssd1 vssd1 vccd1 vccd1 _1890_/S sky130_fd_sc_hd__or2_4
X_2438_ _2479_/CLK _2438_/D vssd1 vssd1 vccd1 vccd1 _2438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2369_ _2369_/CLK _2369_/D vssd1 vssd1 vccd1 vccd1 _2369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1740_ _1740_/A0 _2301_/Q _1740_/S vssd1 vssd1 vccd1 vccd1 _2301_/D sky130_fd_sc_hd__mux2_1
X_1671_ _1726_/A _1911_/A vssd1 vssd1 vccd1 vccd1 _1675_/S sky130_fd_sc_hd__nor2_4
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2223_ _2302_/CLK _2223_/D vssd1 vssd1 vccd1 vccd1 _2223_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2154_ _2159_/CLK _2154_/D vssd1 vssd1 vccd1 vccd1 _2154_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1105_ _2343_/Q _2495_/Q _2423_/Q _2463_/Q _1245_/S0 _1409_/B vssd1 vssd1 vccd1 vccd1
+ _1105_/X sky130_fd_sc_hd__mux4_1
XFILLER_53_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2085_ _2097_/CLK _2085_/D vssd1 vssd1 vccd1 vccd1 _2085_/Q sky130_fd_sc_hd__dfxtp_1
X_1036_ _1409_/C _1034_/X _1035_/X _1298_/B2 vssd1 vssd1 vccd1 vccd1 _1036_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1938_ _1978_/A0 _2459_/Q _1940_/S vssd1 vssd1 vccd1 vccd1 _2459_/D sky130_fd_sc_hd__mux2_1
X_1869_ _2404_/Q _1884_/A0 _1870_/S vssd1 vssd1 vccd1 vccd1 _2404_/D sky130_fd_sc_hd__mux2_1
XFILLER_1_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1723_ _1738_/A0 _2287_/Q _1725_/S vssd1 vssd1 vccd1 vccd1 _2287_/D sky130_fd_sc_hd__mux2_1
X_1654_ _1664_/A0 _2232_/Q _1655_/S vssd1 vssd1 vccd1 vccd1 _2232_/D sky130_fd_sc_hd__mux2_1
X_1585_ _1585_/A0 _2177_/Q _1585_/S vssd1 vssd1 vccd1 vccd1 _2177_/D sky130_fd_sc_hd__mux2_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2206_ _2229_/CLK _2206_/D vssd1 vssd1 vccd1 vccd1 _2206_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2137_ _2240_/CLK _2137_/D vssd1 vssd1 vccd1 vccd1 _2137_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2068_ _2337_/CLK _2068_/D vssd1 vssd1 vccd1 vccd1 _2068_/Q sky130_fd_sc_hd__dfxtp_1
X_1019_ _2434_/Q _2438_/Q _2442_/Q _2446_/Q _1464_/A _1464_/B vssd1 vssd1 vccd1 vccd1
+ _1019_/X sky130_fd_sc_hd__mux4_1
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1370_ _1824_/A0 _2016_/Q _1371_/S vssd1 vssd1 vccd1 vccd1 _2016_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1706_ _1726_/A _1946_/B vssd1 vssd1 vccd1 vccd1 _1710_/S sky130_fd_sc_hd__nor2_2
X_1637_ _1917_/A1 _2218_/Q _1640_/S vssd1 vssd1 vccd1 vccd1 _2218_/D sky130_fd_sc_hd__mux2_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1568_ _2163_/Q _1583_/A0 _1570_/S vssd1 vssd1 vccd1 vccd1 _2163_/D sky130_fd_sc_hd__mux2_1
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1499_ _1784_/A0 _2108_/Q _1500_/S vssd1 vssd1 vccd1 vccd1 _2108_/D sky130_fd_sc_hd__mux2_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout22 _1360_/B vssd1 vssd1 vccd1 vccd1 _1396_/C sky130_fd_sc_hd__buf_8
Xfanout44 input9/X vssd1 vssd1 vccd1 vccd1 fanout44/X sky130_fd_sc_hd__buf_4
Xfanout55 _1977_/A0 vssd1 vssd1 vccd1 vccd1 _1917_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout33 _0993_/Y vssd1 vssd1 vccd1 vccd1 _1258_/A sky130_fd_sc_hd__buf_8
XFILLER_10_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout77 fanout85/X vssd1 vssd1 vccd1 vccd1 _1297_/S1 sky130_fd_sc_hd__buf_6
Xfanout99 _1960_/A0 vssd1 vssd1 vccd1 vccd1 _1905_/A0 sky130_fd_sc_hd__clkbuf_4
Xfanout66 _1742_/A0 vssd1 vssd1 vccd1 vccd1 _1792_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout88 _1283_/S1 vssd1 vssd1 vccd1 vccd1 _1301_/S1 sky130_fd_sc_hd__clkbuf_4
XFILLER_13_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2471_ _2477_/CLK _2471_/D vssd1 vssd1 vccd1 vccd1 _2471_/Q sky130_fd_sc_hd__dfxtp_1
X_1422_ _2050_/Q _1762_/A0 _1425_/S vssd1 vssd1 vccd1 vccd1 _2050_/D sky130_fd_sc_hd__mux2_1
X_1353_ _1354_/A _1398_/B vssd1 vssd1 vccd1 vccd1 _1501_/A sky130_fd_sc_hd__nor2_8
XFILLER_83_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1284_ _1453_/C _1283_/X _1385_/A vssd1 vssd1 vccd1 vccd1 _1284_/X sky130_fd_sc_hd__o21ba_1
XFILLER_83_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0999_ _1409_/B _0996_/X _0998_/X vssd1 vssd1 vccd1 vccd1 _0999_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_59_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1971_ _1971_/A _1976_/A vssd1 vssd1 vccd1 vccd1 _1975_/S sky130_fd_sc_hd__nand2_2
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2454_ _2480_/CLK _2454_/D vssd1 vssd1 vccd1 vccd1 _2454_/Q sky130_fd_sc_hd__dfxtp_1
X_2385_ _2385_/CLK _2385_/D vssd1 vssd1 vccd1 vccd1 _2385_/Q sky130_fd_sc_hd__dfxtp_1
X_1405_ _1792_/A1 _2038_/Q _1408_/S vssd1 vssd1 vccd1 vccd1 _2038_/D sky130_fd_sc_hd__mux2_1
X_1336_ _1660_/A0 _1997_/Q _1336_/S vssd1 vssd1 vccd1 vccd1 _1997_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput1 ram_addr[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__clkbuf_2
XFILLER_56_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1267_ _1267_/A _1267_/B vssd1 vssd1 vccd1 vccd1 _1267_/Y sky130_fd_sc_hd__nor2_1
X_1198_ _2384_/Q _2064_/Q _2104_/Q _2144_/Q _1270_/S _1100_/A vssd1 vssd1 vccd1 vccd1
+ _1199_/B sky130_fd_sc_hd__mux4_1
XFILLER_24_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_39_clk clkbuf_leaf_4_clk/A vssd1 vssd1 vccd1 vccd1 _2449_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2170_ _2177_/CLK _2170_/D vssd1 vssd1 vccd1 vccd1 _2170_/Q sky130_fd_sc_hd__dfxtp_1
X_1121_ _2259_/Q _1987_/Q _1233_/S vssd1 vssd1 vccd1 vccd1 _1121_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1052_ _1220_/A _1052_/B vssd1 vssd1 vccd1 vccd1 _1052_/X sky130_fd_sc_hd__or2_1
XFILLER_65_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1954_ _1964_/A0 _2472_/Q _1955_/S vssd1 vssd1 vccd1 vccd1 _2472_/D sky130_fd_sc_hd__mux2_1
X_1885_ _1905_/A0 _2417_/Q _1885_/S vssd1 vssd1 vccd1 vccd1 _2417_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2437_ _2477_/CLK _2437_/D vssd1 vssd1 vccd1 vccd1 _2437_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2368_ _2368_/CLK _2368_/D vssd1 vssd1 vccd1 vccd1 _2368_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1319_ _1366_/A _1464_/C vssd1 vssd1 vccd1 vccd1 _1951_/A sky130_fd_sc_hd__nor2_8
X_2299_ _2301_/CLK _2299_/D vssd1 vssd1 vccd1 vccd1 _2299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1670_ _2245_/Q _1935_/A0 _1670_/S vssd1 vssd1 vccd1 vccd1 _2245_/D sky130_fd_sc_hd__mux2_1
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2222_ _2302_/CLK _2222_/D vssd1 vssd1 vccd1 vccd1 _2222_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2153_ _2159_/CLK _2153_/D vssd1 vssd1 vccd1 vccd1 _2153_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1104_ _1237_/A _1103_/X _1100_/Y _1102_/Y vssd1 vssd1 vccd1 vccd1 _1104_/X sky130_fd_sc_hd__a2bb2o_1
X_2084_ _2349_/CLK _2084_/D vssd1 vssd1 vccd1 vccd1 _2084_/Q sky130_fd_sc_hd__dfxtp_1
X_1035_ _2386_/Q _2390_/Q _2394_/Q _2398_/Q _1253_/S0 _1256_/S1 vssd1 vssd1 vccd1
+ vccd1 _1035_/X sky130_fd_sc_hd__mux4_1
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1937_ _1977_/A0 _2458_/Q _1940_/S vssd1 vssd1 vccd1 vccd1 _2458_/D sky130_fd_sc_hd__mux2_1
X_1868_ _2403_/Q _1903_/A0 _1870_/S vssd1 vssd1 vccd1 vccd1 _2403_/D sky130_fd_sc_hd__mux2_1
X_1799_ _1809_/A0 _2348_/Q _1800_/S vssd1 vssd1 vccd1 vccd1 _2348_/D sky130_fd_sc_hd__mux2_1
XFILLER_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1722_ _1732_/A0 _2286_/Q _1725_/S vssd1 vssd1 vccd1 vccd1 _2286_/D sky130_fd_sc_hd__mux2_1
X_1653_ _1663_/A0 _2231_/Q _1655_/S vssd1 vssd1 vccd1 vccd1 _2231_/D sky130_fd_sc_hd__mux2_1
X_1584_ _1664_/A0 _2176_/Q _1585_/S vssd1 vssd1 vccd1 vccd1 _2176_/D sky130_fd_sc_hd__mux2_1
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2205_ _2368_/CLK _2205_/D vssd1 vssd1 vccd1 vccd1 _2205_/Q sky130_fd_sc_hd__dfxtp_1
X_2136_ _2232_/CLK _2136_/D vssd1 vssd1 vccd1 vccd1 _2136_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2067_ _2335_/CLK _2067_/D vssd1 vssd1 vccd1 vccd1 _2067_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1018_ _1220_/A _1023_/B vssd1 vssd1 vccd1 vccd1 _1431_/C sky130_fd_sc_hd__or2_4
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1705_ _1740_/A0 _2273_/Q _1705_/S vssd1 vssd1 vccd1 vccd1 _2273_/D sky130_fd_sc_hd__mux2_1
X_1636_ _1646_/A _1956_/B vssd1 vssd1 vccd1 vccd1 _1640_/S sky130_fd_sc_hd__or2_4
X_1567_ _2162_/Q _1582_/A0 _1570_/S vssd1 vssd1 vccd1 vccd1 _2162_/D sky130_fd_sc_hd__mux2_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1498_ _1503_/A0 _2107_/Q _1500_/S vssd1 vssd1 vccd1 vccd1 _2107_/D sky130_fd_sc_hd__mux2_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2119_ _2159_/CLK _2119_/D vssd1 vssd1 vccd1 vccd1 _2119_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout56 input8/X vssd1 vssd1 vccd1 vccd1 _1977_/A0 sky130_fd_sc_hd__buf_4
Xfanout23 _1023_/X vssd1 vssd1 vccd1 vccd1 _1409_/C sky130_fd_sc_hd__buf_8
Xfanout34 _0992_/Y vssd1 vssd1 vccd1 vccd1 _1234_/A1 sky130_fd_sc_hd__buf_4
Xfanout45 _1808_/A0 vssd1 vssd1 vccd1 vccd1 _1823_/A0 sky130_fd_sc_hd__buf_4
Xfanout78 fanout85/X vssd1 vssd1 vccd1 vccd1 _1291_/A sky130_fd_sc_hd__clkbuf_4
Xfanout89 fanout94/X vssd1 vssd1 vccd1 vccd1 _1283_/S1 sky130_fd_sc_hd__buf_4
Xfanout67 fanout68/X vssd1 vssd1 vccd1 vccd1 _1742_/A0 sky130_fd_sc_hd__buf_4
XFILLER_10_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_77 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2470_ _2480_/CLK _2470_/D vssd1 vssd1 vccd1 vccd1 _2470_/Q sky130_fd_sc_hd__dfxtp_1
X_1421_ _1486_/A _1906_/B vssd1 vssd1 vccd1 vccd1 _1425_/S sky130_fd_sc_hd__nor2_4
X_1352_ _1360_/A _1431_/C vssd1 vssd1 vccd1 vccd1 _1681_/B sky130_fd_sc_hd__or2_4
XFILLER_68_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1283_ _2197_/Q _2201_/Q _2205_/Q _2209_/Q _1453_/A _1283_/S1 vssd1 vssd1 vccd1 vccd1
+ _1283_/X sky130_fd_sc_hd__mux4_1
XFILLER_55_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0998_ _1234_/A1 _0997_/X _1241_/B1 vssd1 vssd1 vccd1 vccd1 _0998_/X sky130_fd_sc_hd__a21o_1
X_1619_ _1814_/A0 _2204_/Q _1620_/S vssd1 vssd1 vccd1 vccd1 _2204_/D sky130_fd_sc_hd__mux2_1
XFILLER_59_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1970_ _1975_/A0 _2485_/Q _1970_/S vssd1 vssd1 vccd1 vccd1 _2485_/D sky130_fd_sc_hd__mux2_1
XFILLER_33_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2453_ _2480_/CLK _2453_/D vssd1 vssd1 vccd1 vccd1 _2453_/Q sky130_fd_sc_hd__dfxtp_1
X_1404_ _1971_/A _1941_/B vssd1 vssd1 vccd1 vccd1 _1408_/S sky130_fd_sc_hd__nand2_4
X_2384_ _2496_/CLK _2384_/D vssd1 vssd1 vccd1 vccd1 _2384_/Q sky130_fd_sc_hd__dfxtp_1
X_1335_ _1664_/A0 _1996_/Q _1336_/S vssd1 vssd1 vccd1 vccd1 _1996_/D sky130_fd_sc_hd__mux2_1
Xinput2 ram_addr[1] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__buf_2
XFILLER_56_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1266_ _1409_/C _1264_/X _1265_/X _1305_/B2 vssd1 vssd1 vccd1 vccd1 _1267_/B sky130_fd_sc_hd__a22o_1
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1197_ _1100_/A _1194_/X _1196_/X vssd1 vssd1 vccd1 vccd1 _1197_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_36_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1120_ _2267_/Q _2271_/Q _1240_/S vssd1 vssd1 vccd1 vccd1 _1120_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1051_ _2146_/Q _2150_/Q _2154_/Q _2158_/Q _1292_/S _1297_/S1 vssd1 vssd1 vccd1 vccd1
+ _1052_/B sky130_fd_sc_hd__mux4_1
XFILLER_18_163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1953_ _1963_/A0 _2471_/Q _1955_/S vssd1 vssd1 vccd1 vccd1 _2471_/D sky130_fd_sc_hd__mux2_1
X_1884_ _1884_/A0 _2416_/Q _1885_/S vssd1 vssd1 vccd1 vccd1 _2416_/D sky130_fd_sc_hd__mux2_1
X_2436_ _2482_/CLK _2436_/D vssd1 vssd1 vccd1 vccd1 _2436_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2367_ _2367_/CLK _2367_/D vssd1 vssd1 vccd1 vccd1 _2367_/Q sky130_fd_sc_hd__dfxtp_1
X_2298_ _2301_/CLK _2298_/D vssd1 vssd1 vccd1 vccd1 _2298_/Q sky130_fd_sc_hd__dfxtp_1
X_1318_ _1989_/Q _1935_/A0 _1318_/S vssd1 vssd1 vccd1 vccd1 _1989_/D sky130_fd_sc_hd__mux2_1
X_1249_ _2485_/Q _2489_/Q _2493_/Q _2033_/Q _1253_/S0 _1253_/S1 vssd1 vssd1 vccd1
+ vccd1 _1249_/X sky130_fd_sc_hd__mux4_2
XFILLER_37_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2221_ _2229_/CLK _2221_/D vssd1 vssd1 vccd1 vccd1 _2221_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2152_ _2159_/CLK _2152_/D vssd1 vssd1 vccd1 vccd1 _2152_/Q sky130_fd_sc_hd__dfxtp_1
X_1103_ _2383_/Q _2063_/Q _2103_/Q _2143_/Q _1275_/S0 _1100_/A vssd1 vssd1 vccd1 vccd1
+ _1103_/X sky130_fd_sc_hd__mux4_1
X_2083_ _2097_/CLK _2083_/D vssd1 vssd1 vccd1 vccd1 _2083_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1034_ _2418_/Q _2022_/Q _2426_/Q _2430_/Q _1256_/S0 _1253_/S1 vssd1 vssd1 vccd1
+ vccd1 _1034_/X sky130_fd_sc_hd__mux4_2
XFILLER_19_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1936_ _1966_/A _1936_/B vssd1 vssd1 vccd1 vccd1 _1940_/S sky130_fd_sc_hd__or2_4
X_1867_ _2402_/Q _1902_/A0 _1870_/S vssd1 vssd1 vccd1 vccd1 _2402_/D sky130_fd_sc_hd__mux2_1
X_1798_ _1808_/A0 _2347_/Q _1800_/S vssd1 vssd1 vccd1 vccd1 _2347_/D sky130_fd_sc_hd__mux2_1
XFILLER_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2419_ _2421_/CLK _2419_/D vssd1 vssd1 vccd1 vccd1 _2419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1721_ _1736_/A _1961_/A vssd1 vssd1 vccd1 vccd1 _1725_/S sky130_fd_sc_hd__nand2_4
X_1652_ _1662_/A0 _2230_/Q _1655_/S vssd1 vssd1 vccd1 vccd1 _2230_/D sky130_fd_sc_hd__mux2_1
X_1583_ _1583_/A0 _2175_/Q _1585_/S vssd1 vssd1 vccd1 vccd1 _2175_/D sky130_fd_sc_hd__mux2_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2204_ _2368_/CLK _2204_/D vssd1 vssd1 vccd1 vccd1 _2204_/Q sky130_fd_sc_hd__dfxtp_1
X_2135_ _2177_/CLK _2135_/D vssd1 vssd1 vccd1 vccd1 _2135_/Q sky130_fd_sc_hd__dfxtp_1
X_2066_ _2335_/CLK _2066_/D vssd1 vssd1 vccd1 vccd1 _2066_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1017_ _1274_/A _1023_/B vssd1 vssd1 vccd1 vccd1 _1017_/Y sky130_fd_sc_hd__nor2_1
XFILLER_22_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1919_ _2444_/Q _1974_/A0 _1920_/S vssd1 vssd1 vccd1 vccd1 _2444_/D sky130_fd_sc_hd__mux2_1
XFILLER_1_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1704_ _1739_/A0 _2272_/Q _1705_/S vssd1 vssd1 vccd1 vccd1 _2272_/D sky130_fd_sc_hd__mux2_1
X_1635_ _1660_/A0 _2217_/Q _1635_/S vssd1 vssd1 vccd1 vccd1 _2217_/D sky130_fd_sc_hd__mux2_1
X_1566_ _1566_/A _1966_/B vssd1 vssd1 vccd1 vccd1 _1570_/S sky130_fd_sc_hd__nor2_4
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1497_ _1777_/A0 _2106_/Q _1500_/S vssd1 vssd1 vccd1 vccd1 _2106_/D sky130_fd_sc_hd__mux2_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2118_ _2232_/CLK _2118_/D vssd1 vssd1 vccd1 vccd1 _2118_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2049_ _2049_/CLK _2049_/D vssd1 vssd1 vccd1 vccd1 _2049_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout35 _0992_/Y vssd1 vssd1 vccd1 vccd1 _1475_/B sky130_fd_sc_hd__buf_8
Xfanout24 _1475_/C vssd1 vssd1 vccd1 vccd1 _1464_/C sky130_fd_sc_hd__buf_6
Xfanout46 _1808_/A0 vssd1 vssd1 vccd1 vccd1 _1503_/A0 sky130_fd_sc_hd__buf_4
XFILLER_13_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout79 fanout85/X vssd1 vssd1 vccd1 vccd1 _1013_/B sky130_fd_sc_hd__buf_8
Xfanout68 input8/X vssd1 vssd1 vccd1 vccd1 fanout68/X sky130_fd_sc_hd__clkbuf_4
Xfanout57 _1777_/A0 vssd1 vssd1 vccd1 vccd1 _1762_/A0 sky130_fd_sc_hd__clkbuf_4
XFILLER_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1420_ _1420_/A _1442_/B _1420_/C vssd1 vssd1 vccd1 vccd1 _1906_/B sky130_fd_sc_hd__or3_4
X_1351_ _1360_/A _1431_/C vssd1 vssd1 vccd1 vccd1 _1921_/A sky130_fd_sc_hd__nor2_8
X_1282_ _1398_/A _1282_/B vssd1 vssd1 vccd1 vccd1 _1282_/Y sky130_fd_sc_hd__nor2_1
XFILLER_36_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0997_ _2258_/Q _1986_/Q _1240_/S vssd1 vssd1 vccd1 vccd1 _0997_/X sky130_fd_sc_hd__mux2_1
X_1618_ _1823_/A0 _2203_/Q _1620_/S vssd1 vssd1 vccd1 vccd1 _2203_/D sky130_fd_sc_hd__mux2_1
X_1549_ _2148_/Q _1974_/A0 _1550_/S vssd1 vssd1 vccd1 vccd1 _2148_/D sky130_fd_sc_hd__mux2_1
XFILLER_27_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2452_ _2480_/CLK _2452_/D vssd1 vssd1 vccd1 vccd1 _2452_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2383_ _2496_/CLK _2383_/D vssd1 vssd1 vccd1 vccd1 _2383_/Q sky130_fd_sc_hd__dfxtp_1
X_1403_ _2037_/Q _1845_/A1 _1403_/S vssd1 vssd1 vccd1 vccd1 _2037_/D sky130_fd_sc_hd__mux2_1
X_1334_ _1663_/A0 _1995_/Q _1336_/S vssd1 vssd1 vccd1 vccd1 _1995_/D sky130_fd_sc_hd__mux2_1
X_1265_ _2309_/Q _2313_/Q _2317_/Q _2321_/Q _1285_/S0 _1285_/S1 vssd1 vssd1 vccd1
+ vccd1 _1265_/X sky130_fd_sc_hd__mux4_2
Xinput3 ram_addr[2] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_2
X_1196_ _1234_/A1 _1195_/X _1020_/A vssd1 vssd1 vccd1 vccd1 _1196_/X sky130_fd_sc_hd__a21o_1
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1050_ _2162_/Q _2166_/Q _2170_/Q _2174_/Q _1297_/S0 _1297_/S1 vssd1 vssd1 vccd1
+ vccd1 _1050_/X sky130_fd_sc_hd__mux4_2
XFILLER_18_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1952_ _1962_/A0 _2470_/Q _1955_/S vssd1 vssd1 vccd1 vccd1 _2470_/D sky130_fd_sc_hd__mux2_1
X_1883_ _1903_/A0 _2415_/Q _1885_/S vssd1 vssd1 vccd1 vccd1 _2415_/D sky130_fd_sc_hd__mux2_1
X_2435_ _2482_/CLK _2435_/D vssd1 vssd1 vccd1 vccd1 _2435_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2366_ _2368_/CLK _2366_/D vssd1 vssd1 vccd1 vccd1 _2366_/Q sky130_fd_sc_hd__dfxtp_1
X_2297_ _2297_/CLK _2297_/D vssd1 vssd1 vccd1 vccd1 _2297_/Q sky130_fd_sc_hd__dfxtp_1
X_1317_ _1988_/Q _1739_/A0 _1318_/S vssd1 vssd1 vccd1 vccd1 _1988_/D sky130_fd_sc_hd__mux2_1
XFILLER_56_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1248_ _2469_/Q _2473_/Q _2477_/Q _2481_/Q _1475_/A _1464_/B vssd1 vssd1 vccd1 vccd1
+ _1248_/X sky130_fd_sc_hd__mux4_2
XFILLER_37_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1179_ _2276_/Q _2280_/Q _2284_/Q _2288_/Q _1181_/S _0992_/A vssd1 vssd1 vccd1 vccd1
+ _1180_/B sky130_fd_sc_hd__mux4_1
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2220_ _2229_/CLK _2220_/D vssd1 vssd1 vccd1 vccd1 _2220_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2151_ _2493_/CLK _2151_/D vssd1 vssd1 vccd1 vccd1 _2151_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1102_ _1234_/A1 _1101_/X _1241_/B1 vssd1 vssd1 vccd1 vccd1 _1102_/Y sky130_fd_sc_hd__a21oi_1
X_2082_ _2097_/CLK _2082_/D vssd1 vssd1 vccd1 vccd1 _2082_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1033_ _1020_/X _1029_/X _1031_/X _1032_/X _1295_/B2 vssd1 vssd1 vccd1 vccd1 _1033_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1935_ _1935_/A0 _2457_/Q _1935_/S vssd1 vssd1 vccd1 vccd1 _2457_/D sky130_fd_sc_hd__mux2_1
X_1866_ _1886_/A _1946_/B vssd1 vssd1 vccd1 vccd1 _1870_/S sky130_fd_sc_hd__nor2_4
X_1797_ _1822_/A0 _2346_/Q _1800_/S vssd1 vssd1 vccd1 vccd1 _2346_/D sky130_fd_sc_hd__mux2_1
X_2418_ _2433_/CLK _2418_/D vssd1 vssd1 vccd1 vccd1 _2418_/Q sky130_fd_sc_hd__dfxtp_1
X_2349_ _2349_/CLK _2349_/D vssd1 vssd1 vccd1 vccd1 _2349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1720_ _2285_/Q _1960_/A0 _1720_/S vssd1 vssd1 vccd1 vccd1 _2285_/D sky130_fd_sc_hd__mux2_1
X_1651_ _1661_/A _1971_/A vssd1 vssd1 vccd1 vccd1 _1655_/S sky130_fd_sc_hd__nand2_2
X_1582_ _1582_/A0 _2174_/Q _1585_/S vssd1 vssd1 vccd1 vccd1 _2174_/D sky130_fd_sc_hd__mux2_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2203_ _2368_/CLK _2203_/D vssd1 vssd1 vccd1 vccd1 _2203_/Q sky130_fd_sc_hd__dfxtp_1
X_2134_ _2232_/CLK _2134_/D vssd1 vssd1 vccd1 vccd1 _2134_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2065_ _2385_/CLK _2065_/D vssd1 vssd1 vccd1 vccd1 _2065_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1016_ _1453_/C _1015_/X _1385_/A vssd1 vssd1 vccd1 vccd1 _1016_/X sky130_fd_sc_hd__o21ba_1
XFILLER_22_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1918_ _2443_/Q _1918_/A1 _1920_/S vssd1 vssd1 vccd1 vccd1 _2443_/D sky130_fd_sc_hd__mux2_1
X_1849_ _2388_/Q _1904_/A0 _1850_/S vssd1 vssd1 vccd1 vccd1 _2388_/D sky130_fd_sc_hd__mux2_1
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_20_clk clkbuf_2_3__f_clk/X vssd1 vssd1 vccd1 vccd1 _2385_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_11_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _2097_/CLK sky130_fd_sc_hd__clkbuf_16
X_1703_ _1793_/A1 _2271_/Q _1705_/S vssd1 vssd1 vccd1 vccd1 _2271_/D sky130_fd_sc_hd__mux2_1
X_1634_ _1979_/A0 _2216_/Q _1635_/S vssd1 vssd1 vccd1 vccd1 _2216_/D sky130_fd_sc_hd__mux2_1
X_1565_ _1980_/A0 _2161_/Q _1565_/S vssd1 vssd1 vccd1 vccd1 _2161_/D sky130_fd_sc_hd__mux2_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1496_ _1501_/A _1976_/B vssd1 vssd1 vccd1 vccd1 _1500_/S sky130_fd_sc_hd__nand2_4
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2117_ _2448_/CLK _2117_/D vssd1 vssd1 vccd1 vccd1 _2117_/Q sky130_fd_sc_hd__dfxtp_1
X_2048_ _2049_/CLK _2048_/D vssd1 vssd1 vccd1 vccd1 _2048_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout36 _1918_/A1 vssd1 vssd1 vccd1 vccd1 _1583_/A0 sky130_fd_sc_hd__clkbuf_4
Xfanout25 _1431_/C vssd1 vssd1 vccd1 vccd1 _1420_/C sky130_fd_sc_hd__buf_6
Xfanout47 _1808_/A0 vssd1 vssd1 vccd1 vccd1 _1778_/A0 sky130_fd_sc_hd__buf_2
Xfanout69 input5/X vssd1 vssd1 vccd1 vccd1 _1040_/B sky130_fd_sc_hd__buf_8
Xfanout58 _1777_/A0 vssd1 vssd1 vccd1 vccd1 _1822_/A0 sky130_fd_sc_hd__clkbuf_4
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1350_ _1585_/A0 _2005_/Q _1350_/S vssd1 vssd1 vccd1 vccd1 _2005_/D sky130_fd_sc_hd__mux2_1
X_1281_ _1023_/B _1272_/Y _1274_/Y _1279_/Y _1280_/Y vssd1 vssd1 vccd1 vccd1 _1282_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_76_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_0_clk clkbuf_leaf_4_clk/A vssd1 vssd1 vccd1 vccd1 _2232_/CLK sky130_fd_sc_hd__clkbuf_16
X_0996_ _2266_/Q _2270_/Q _1240_/S vssd1 vssd1 vccd1 vccd1 _0996_/X sky130_fd_sc_hd__mux2_1
X_1617_ _1917_/A1 _2202_/Q _1620_/S vssd1 vssd1 vccd1 vccd1 _2202_/D sky130_fd_sc_hd__mux2_1
X_1548_ _2147_/Q _1918_/A1 _1550_/S vssd1 vssd1 vccd1 vccd1 _2147_/D sky130_fd_sc_hd__mux2_1
XFILLER_59_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1479_ _2092_/Q _1824_/A0 _1480_/S vssd1 vssd1 vccd1 vccd1 _2092_/D sky130_fd_sc_hd__mux2_1
XFILLER_54_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2451_ _2480_/CLK _2451_/D vssd1 vssd1 vccd1 vccd1 _2451_/Q sky130_fd_sc_hd__dfxtp_1
X_1402_ _2036_/Q _1984_/A1 _1403_/S vssd1 vssd1 vccd1 vccd1 _2036_/D sky130_fd_sc_hd__mux2_1
X_2382_ _2385_/CLK _2382_/D vssd1 vssd1 vccd1 vccd1 _2382_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1333_ _1917_/A1 _1994_/Q _1336_/S vssd1 vssd1 vccd1 vccd1 _1994_/D sky130_fd_sc_hd__mux2_1
X_1264_ _2357_/Q _2361_/Q _2365_/Q _2369_/Q _1453_/A _1283_/S1 vssd1 vssd1 vccd1 vccd1
+ _1264_/X sky130_fd_sc_hd__mux4_1
Xinput4 ram_addr[3] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_8
X_1195_ _2184_/Q _2224_/Q _1270_/S vssd1 vssd1 vccd1 vccd1 _1195_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_2_1__f_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_9_clk/A sky130_fd_sc_hd__clkbuf_16
XFILLER_17_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_77 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1951_ _1951_/A _1976_/A vssd1 vssd1 vccd1 vccd1 _1955_/S sky130_fd_sc_hd__nand2_4
X_1882_ _1902_/A0 _2414_/Q _1885_/S vssd1 vssd1 vccd1 vccd1 _2414_/D sky130_fd_sc_hd__mux2_1
X_2434_ _2479_/CLK _2434_/D vssd1 vssd1 vccd1 vccd1 _2434_/Q sky130_fd_sc_hd__dfxtp_1
X_2365_ _2369_/CLK _2365_/D vssd1 vssd1 vccd1 vccd1 _2365_/Q sky130_fd_sc_hd__dfxtp_1
X_1316_ _1987_/Q _1983_/A1 _1318_/S vssd1 vssd1 vccd1 vccd1 _1987_/D sky130_fd_sc_hd__mux2_1
XFILLER_84_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2296_ _2296_/CLK _2296_/D vssd1 vssd1 vccd1 vccd1 _2296_/Q sky130_fd_sc_hd__dfxtp_1
X_1247_ _2437_/Q _2441_/Q _2445_/Q _2449_/Q _1464_/A _1442_/B vssd1 vssd1 vccd1 vccd1
+ _1247_/X sky130_fd_sc_hd__mux4_1
X_1178_ _1180_/A _1177_/X _1244_/A1 vssd1 vssd1 vccd1 vccd1 _1178_/X sky130_fd_sc_hd__o21ba_1
XFILLER_52_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2150_ _2448_/CLK _2150_/D vssd1 vssd1 vccd1 vccd1 _2150_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1101_ _2183_/Q _2223_/Q _1270_/S vssd1 vssd1 vccd1 vccd1 _1101_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2081_ _2097_/CLK _2081_/D vssd1 vssd1 vccd1 vccd1 _2081_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1032_ _2370_/Q _2374_/Q _2378_/Q _2018_/Q _1253_/S0 _1253_/S1 vssd1 vssd1 vccd1
+ vccd1 _1032_/X sky130_fd_sc_hd__mux4_1
XFILLER_19_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1934_ _1964_/A0 _2456_/Q _1935_/S vssd1 vssd1 vccd1 vccd1 _2456_/D sky130_fd_sc_hd__mux2_1
X_1865_ _1975_/A0 _2401_/Q _1865_/S vssd1 vssd1 vccd1 vccd1 _2401_/D sky130_fd_sc_hd__mux2_1
X_1796_ _1806_/A _1956_/B vssd1 vssd1 vccd1 vccd1 _1800_/S sky130_fd_sc_hd__or2_2
X_2417_ _2433_/CLK _2417_/D vssd1 vssd1 vccd1 vccd1 _2417_/Q sky130_fd_sc_hd__dfxtp_1
X_2348_ _2369_/CLK _2348_/D vssd1 vssd1 vccd1 vccd1 _2348_/Q sky130_fd_sc_hd__dfxtp_1
X_2279_ _2481_/CLK _2279_/D vssd1 vssd1 vccd1 vccd1 _2279_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1650_ _1660_/A0 _2229_/Q _1650_/S vssd1 vssd1 vccd1 vccd1 _2229_/D sky130_fd_sc_hd__mux2_1
X_1581_ _1581_/A _1901_/A vssd1 vssd1 vccd1 vccd1 _1585_/S sky130_fd_sc_hd__nand2_4
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2202_ _2229_/CLK _2202_/D vssd1 vssd1 vccd1 vccd1 _2202_/Q sky130_fd_sc_hd__dfxtp_1
X_2133_ _2232_/CLK _2133_/D vssd1 vssd1 vccd1 vccd1 _2133_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2064_ _2496_/CLK _2064_/D vssd1 vssd1 vccd1 vccd1 _2064_/Q sky130_fd_sc_hd__dfxtp_1
X_1015_ _2450_/Q _2454_/Q _2458_/Q _2026_/Q _1245_/S0 _1409_/B vssd1 vssd1 vccd1 vccd1
+ _1015_/X sky130_fd_sc_hd__mux4_1
X_1917_ _2442_/Q _1917_/A1 _1920_/S vssd1 vssd1 vccd1 vccd1 _2442_/D sky130_fd_sc_hd__mux2_1
X_1848_ _2387_/Q _1903_/A0 _1850_/S vssd1 vssd1 vccd1 vccd1 _2387_/D sky130_fd_sc_hd__mux2_1
X_1779_ _1784_/A0 _2332_/Q _1780_/S vssd1 vssd1 vccd1 vccd1 _2332_/D sky130_fd_sc_hd__mux2_1
XFILLER_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1702_ _1792_/A1 _2270_/Q _1705_/S vssd1 vssd1 vccd1 vccd1 _2270_/D sky130_fd_sc_hd__mux2_1
X_1633_ _1978_/A0 _2215_/Q _1635_/S vssd1 vssd1 vccd1 vccd1 _2215_/D sky130_fd_sc_hd__mux2_1
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1564_ _1974_/A0 _2160_/Q _1565_/S vssd1 vssd1 vccd1 vccd1 _2160_/D sky130_fd_sc_hd__mux2_1
X_1495_ _2105_/Q _1985_/A1 _1495_/S vssd1 vssd1 vccd1 vccd1 _2105_/D sky130_fd_sc_hd__mux2_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2116_ _2159_/CLK _2116_/D vssd1 vssd1 vccd1 vccd1 _2116_/Q sky130_fd_sc_hd__dfxtp_1
X_2047_ _2261_/CLK _2047_/D vssd1 vssd1 vccd1 vccd1 _2047_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout37 _1978_/A0 vssd1 vssd1 vccd1 vccd1 _1918_/A1 sky130_fd_sc_hd__buf_4
Xfanout26 _1017_/Y vssd1 vssd1 vccd1 vccd1 _1295_/B2 sky130_fd_sc_hd__buf_6
Xfanout59 input8/X vssd1 vssd1 vccd1 vccd1 _1777_/A0 sky130_fd_sc_hd__buf_4
Xfanout48 input9/X vssd1 vssd1 vccd1 vccd1 _1808_/A0 sky130_fd_sc_hd__buf_4
XFILLER_1_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1280_ _1274_/A _1275_/X _1023_/B vssd1 vssd1 vccd1 vccd1 _1280_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0995_ _1040_/B input6/X vssd1 vssd1 vccd1 vccd1 _1398_/A sky130_fd_sc_hd__or2_4
XFILLER_8_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1616_ _1646_/A _1936_/B vssd1 vssd1 vccd1 vccd1 _1620_/S sky130_fd_sc_hd__or2_4
X_1547_ _2146_/Q _1977_/A0 _1550_/S vssd1 vssd1 vccd1 vccd1 _2146_/D sky130_fd_sc_hd__mux2_1
X_1478_ _2091_/Q _1503_/A0 _1480_/S vssd1 vssd1 vccd1 vccd1 _2091_/D sky130_fd_sc_hd__mux2_1
XFILLER_39_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2450_ _2480_/CLK _2450_/D vssd1 vssd1 vccd1 vccd1 _2450_/Q sky130_fd_sc_hd__dfxtp_1
X_1401_ _2035_/Q _1783_/A0 _1403_/S vssd1 vssd1 vccd1 vccd1 _2035_/D sky130_fd_sc_hd__mux2_1
X_2381_ _2482_/CLK _2381_/D vssd1 vssd1 vccd1 vccd1 _2381_/Q sky130_fd_sc_hd__dfxtp_1
X_1332_ _1961_/A _1661_/A vssd1 vssd1 vccd1 vccd1 _1336_/S sky130_fd_sc_hd__nand2_2
XFILLER_68_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1263_ _1302_/A1 _1261_/X _1262_/X _1020_/X vssd1 vssd1 vccd1 vccd1 _1267_/A sky130_fd_sc_hd__a22o_1
Xinput5 ram_addr[4] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__buf_2
XFILLER_49_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1194_ _2264_/Q _2304_/Q _1270_/S vssd1 vssd1 vccd1 vccd1 _1194_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1950_ _2469_/Q _1960_/A0 _1950_/S vssd1 vssd1 vccd1 vccd1 _2469_/D sky130_fd_sc_hd__mux2_1
X_1881_ _1961_/A _1901_/B vssd1 vssd1 vccd1 vccd1 _1885_/S sky130_fd_sc_hd__nand2_2
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2433_ _2433_/CLK _2433_/D vssd1 vssd1 vccd1 vccd1 _2433_/Q sky130_fd_sc_hd__dfxtp_1
X_2364_ _2368_/CLK _2364_/D vssd1 vssd1 vccd1 vccd1 _2364_/Q sky130_fd_sc_hd__dfxtp_1
X_1315_ _1986_/Q _1792_/A1 _1318_/S vssd1 vssd1 vccd1 vccd1 _1986_/D sky130_fd_sc_hd__mux2_1
X_2295_ _2296_/CLK _2295_/D vssd1 vssd1 vccd1 vccd1 _2295_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1246_ _1310_/A _1245_/X _1385_/A vssd1 vssd1 vccd1 vccd1 _1246_/X sky130_fd_sc_hd__o21ba_1
X_1177_ _2244_/Q _2248_/Q _2252_/Q _2256_/Q _1475_/A _1464_/B vssd1 vssd1 vccd1 vccd1
+ _1177_/X sky130_fd_sc_hd__mux4_1
XFILLER_64_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1100_ _1100_/A _1100_/B vssd1 vssd1 vccd1 vccd1 _1100_/Y sky130_fd_sc_hd__nand2_1
X_2080_ _2349_/CLK _2080_/D vssd1 vssd1 vccd1 vccd1 _2080_/Q sky130_fd_sc_hd__dfxtp_1
X_1031_ _1475_/B _1031_/B vssd1 vssd1 vccd1 vccd1 _1031_/X sky130_fd_sc_hd__or2_1
XFILLER_19_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1933_ _1963_/A0 _2455_/Q _1935_/S vssd1 vssd1 vccd1 vccd1 _2455_/D sky130_fd_sc_hd__mux2_1
X_1864_ _1969_/A0 _2400_/Q _1865_/S vssd1 vssd1 vccd1 vccd1 _2400_/D sky130_fd_sc_hd__mux2_1
X_1795_ _2345_/Q _1985_/A1 _1795_/S vssd1 vssd1 vccd1 vccd1 _2345_/D sky130_fd_sc_hd__mux2_1
X_2416_ _2416_/CLK _2416_/D vssd1 vssd1 vccd1 vccd1 _2416_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2347_ _2369_/CLK _2347_/D vssd1 vssd1 vccd1 vccd1 _2347_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2278_ _2296_/CLK _2278_/D vssd1 vssd1 vccd1 vccd1 _2278_/Q sky130_fd_sc_hd__dfxtp_1
X_1229_ _1225_/X _1228_/X _1354_/A vssd1 vssd1 vccd1 vccd1 _1230_/D sky130_fd_sc_hd__o21ba_1
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1580_ _1585_/A0 _2173_/Q _1580_/S vssd1 vssd1 vccd1 vccd1 _2173_/D sky130_fd_sc_hd__mux2_1
XFILLER_7_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2201_ _2457_/CLK _2201_/D vssd1 vssd1 vccd1 vccd1 _2201_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2132_ _2232_/CLK _2132_/D vssd1 vssd1 vccd1 vccd1 _2132_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2063_ _2385_/CLK _2063_/D vssd1 vssd1 vccd1 vccd1 _2063_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1014_ _1464_/A _1475_/B vssd1 vssd1 vccd1 vccd1 _1366_/A sky130_fd_sc_hd__nand2_8
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1916_ _1966_/A _1916_/B vssd1 vssd1 vccd1 vccd1 _1920_/S sky130_fd_sc_hd__nor2_2
XFILLER_8_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1847_ _2386_/Q _1902_/A0 _1850_/S vssd1 vssd1 vccd1 vccd1 _2386_/D sky130_fd_sc_hd__mux2_1
X_1778_ _1778_/A0 _2331_/Q _1780_/S vssd1 vssd1 vccd1 vccd1 _2331_/D sky130_fd_sc_hd__mux2_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1701_ _1736_/A _1861_/A vssd1 vssd1 vccd1 vccd1 _1705_/S sky130_fd_sc_hd__nand2_4
X_1632_ _1917_/A1 _2214_/Q _1635_/S vssd1 vssd1 vccd1 vccd1 _2214_/D sky130_fd_sc_hd__mux2_1
X_1563_ _1918_/A1 _2159_/Q _1565_/S vssd1 vssd1 vccd1 vccd1 _2159_/D sky130_fd_sc_hd__mux2_1
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1494_ _2104_/Q _1804_/A0 _1495_/S vssd1 vssd1 vccd1 vccd1 _2104_/D sky130_fd_sc_hd__mux2_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2115_ _2176_/CLK _2115_/D vssd1 vssd1 vccd1 vccd1 _2115_/Q sky130_fd_sc_hd__dfxtp_1
X_2046_ _2261_/CLK _2046_/D vssd1 vssd1 vccd1 vccd1 _2046_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout38 _1978_/A0 vssd1 vssd1 vccd1 vccd1 _1663_/A0 sky130_fd_sc_hd__clkbuf_4
Xfanout27 _1017_/Y vssd1 vssd1 vccd1 vccd1 _1305_/B2 sky130_fd_sc_hd__buf_2
Xfanout49 _1843_/A1 vssd1 vssd1 vccd1 vccd1 _1983_/A1 sky130_fd_sc_hd__buf_4
XFILLER_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0994_ _1040_/B input6/X vssd1 vssd1 vccd1 vccd1 _0994_/Y sky130_fd_sc_hd__nor2_1
X_1615_ _1940_/A0 _2201_/Q _1615_/S vssd1 vssd1 vccd1 vccd1 _2201_/D sky130_fd_sc_hd__mux2_1
X_1546_ _1566_/A _1946_/B vssd1 vssd1 vccd1 vccd1 _1550_/S sky130_fd_sc_hd__nor2_4
X_1477_ _2090_/Q _1762_/A0 _1480_/S vssd1 vssd1 vccd1 vccd1 _2090_/D sky130_fd_sc_hd__mux2_1
XFILLER_27_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2029_ _2457_/CLK _2029_/D vssd1 vssd1 vccd1 vccd1 _2029_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1400_ _2034_/Q _1792_/A1 _1403_/S vssd1 vssd1 vccd1 vccd1 _2034_/D sky130_fd_sc_hd__mux2_1
X_2380_ _2485_/CLK _2380_/D vssd1 vssd1 vccd1 vccd1 _2380_/Q sky130_fd_sc_hd__dfxtp_1
X_1331_ _1385_/A _1398_/B vssd1 vssd1 vccd1 vccd1 _1646_/A sky130_fd_sc_hd__or2_4
X_1262_ _2341_/Q _1993_/Q _2349_/Q _2353_/Q _1304_/S0 _1065_/A vssd1 vssd1 vccd1 vccd1
+ _1262_/X sky130_fd_sc_hd__mux4_1
Xinput6 ram_addr[5] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__buf_8
XFILLER_49_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1193_ _0994_/Y _1185_/X _1192_/X _1172_/X vssd1 vssd1 vccd1 vccd1 _1193_/X sky130_fd_sc_hd__a211o_1
XFILLER_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1529_ _2132_/Q _1579_/A0 _1530_/S vssd1 vssd1 vccd1 vccd1 _2132_/D sky130_fd_sc_hd__mux2_1
XFILLER_27_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1880_ _1905_/A0 _2413_/Q _1880_/S vssd1 vssd1 vccd1 vccd1 _2413_/D sky130_fd_sc_hd__mux2_1
XFILLER_41_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2432_ _2432_/CLK _2432_/D vssd1 vssd1 vccd1 vccd1 _2432_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2363_ _2363_/CLK _2363_/D vssd1 vssd1 vccd1 vccd1 _2363_/Q sky130_fd_sc_hd__dfxtp_1
X_1314_ _1641_/A _1726_/A vssd1 vssd1 vccd1 vccd1 _1318_/S sky130_fd_sc_hd__nor2_2
X_2294_ _2297_/CLK _2294_/D vssd1 vssd1 vccd1 vccd1 _2294_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1245_ _2453_/Q _2457_/Q _2461_/Q _2029_/Q _1245_/S0 _1409_/B vssd1 vssd1 vccd1 vccd1
+ _1245_/X sky130_fd_sc_hd__mux4_1
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1176_ _1234_/A1 _1175_/X _1174_/X _1241_/B1 vssd1 vssd1 vccd1 vccd1 _1176_/X sky130_fd_sc_hd__a211o_1
XFILLER_52_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1030_ _2410_/Q _2414_/Q _1181_/S vssd1 vssd1 vccd1 vccd1 _1031_/B sky130_fd_sc_hd__mux2_1
XFILLER_61_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_41_clk clkbuf_leaf_4_clk/A vssd1 vssd1 vccd1 vccd1 _2493_/CLK sky130_fd_sc_hd__clkbuf_16
X_1932_ _1962_/A0 _2454_/Q _1935_/S vssd1 vssd1 vccd1 vccd1 _2454_/D sky130_fd_sc_hd__mux2_1
X_1863_ _1973_/A0 _2399_/Q _1865_/S vssd1 vssd1 vccd1 vccd1 _2399_/D sky130_fd_sc_hd__mux2_1
X_1794_ _2344_/Q _1984_/A1 _1795_/S vssd1 vssd1 vccd1 vccd1 _2344_/D sky130_fd_sc_hd__mux2_1
X_2415_ _2416_/CLK _2415_/D vssd1 vssd1 vccd1 vccd1 _2415_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2346_ _2369_/CLK _2346_/D vssd1 vssd1 vccd1 vccd1 _2346_/Q sky130_fd_sc_hd__dfxtp_1
X_2277_ _2416_/CLK _2277_/D vssd1 vssd1 vccd1 vccd1 _2277_/Q sky130_fd_sc_hd__dfxtp_1
X_1228_ _1409_/C _1226_/X _1227_/X _1305_/B2 vssd1 vssd1 vccd1 vccd1 _1228_/X sky130_fd_sc_hd__a22o_1
X_1159_ _2420_/Q _2024_/Q _2428_/Q _2432_/Q _1256_/S0 _1256_/S1 vssd1 vssd1 vccd1
+ vccd1 _1159_/X sky130_fd_sc_hd__mux4_2
XFILLER_25_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_32_clk clkbuf_2_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _2432_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_23_clk clkbuf_2_3__f_clk/X vssd1 vssd1 vccd1 vccd1 _2049_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2200_ _2461_/CLK _2200_/D vssd1 vssd1 vccd1 vccd1 _2200_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2131_ _2177_/CLK _2131_/D vssd1 vssd1 vccd1 vccd1 _2131_/Q sky130_fd_sc_hd__dfxtp_1
X_2062_ _2385_/CLK _2062_/D vssd1 vssd1 vccd1 vccd1 _2062_/Q sky130_fd_sc_hd__dfxtp_1
X_1013_ _1464_/A _1013_/B vssd1 vssd1 vccd1 vccd1 _1360_/A sky130_fd_sc_hd__nand2_8
XFILLER_34_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1915_ _2441_/Q _1980_/A0 _1915_/S vssd1 vssd1 vccd1 vccd1 _2441_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_14_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _2349_/CLK sky130_fd_sc_hd__clkbuf_16
X_1846_ _1886_/A _1926_/B vssd1 vssd1 vccd1 vccd1 _1850_/S sky130_fd_sc_hd__nor2_2
X_1777_ _1777_/A0 _2330_/Q _1780_/S vssd1 vssd1 vccd1 vccd1 _2330_/D sky130_fd_sc_hd__mux2_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2329_ _2329_/CLK _2329_/D vssd1 vssd1 vccd1 vccd1 _2329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1700_ _2269_/Q _1740_/A0 _1700_/S vssd1 vssd1 vccd1 vccd1 _2269_/D sky130_fd_sc_hd__mux2_1
XFILLER_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1631_ _1951_/A _1661_/A vssd1 vssd1 vccd1 vccd1 _1635_/S sky130_fd_sc_hd__nand2_2
X_1562_ _1977_/A0 _2158_/Q _1565_/S vssd1 vssd1 vccd1 vccd1 _2158_/D sky130_fd_sc_hd__mux2_1
X_1493_ _2103_/Q _1783_/A0 _1495_/S vssd1 vssd1 vccd1 vccd1 _2103_/D sky130_fd_sc_hd__mux2_1
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_3_clk clkbuf_leaf_4_clk/A vssd1 vssd1 vccd1 vccd1 _2229_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2114_ _2229_/CLK _2114_/D vssd1 vssd1 vccd1 vccd1 _2114_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2045_ _2496_/CLK _2045_/D vssd1 vssd1 vccd1 vccd1 _2045_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout28 _1310_/A vssd1 vssd1 vccd1 vccd1 _1453_/C sky130_fd_sc_hd__buf_6
Xfanout17 _1691_/A vssd1 vssd1 vccd1 vccd1 _1981_/B sky130_fd_sc_hd__clkbuf_16
Xfanout39 fanout44/X vssd1 vssd1 vccd1 vccd1 _1978_/A0 sky130_fd_sc_hd__buf_4
XFILLER_10_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1829_ _2372_/Q _1969_/A0 _1830_/S vssd1 vssd1 vccd1 vccd1 _2372_/D sky130_fd_sc_hd__mux2_1
XFILLER_8_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0993_ _1274_/A vssd1 vssd1 vccd1 vccd1 _0993_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1614_ _1809_/A0 _2200_/Q _1615_/S vssd1 vssd1 vccd1 vccd1 _2200_/D sky130_fd_sc_hd__mux2_1
X_1545_ _2145_/Q _1985_/A1 _1545_/S vssd1 vssd1 vccd1 vccd1 _2145_/D sky130_fd_sc_hd__mux2_1
XFILLER_39_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1476_ _1486_/A _1956_/B vssd1 vssd1 vccd1 vccd1 _1480_/S sky130_fd_sc_hd__nor2_2
XFILLER_67_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2028_ _2479_/CLK _2028_/D vssd1 vssd1 vccd1 vccd1 _2028_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1330_ _1385_/A _1398_/B vssd1 vssd1 vccd1 vccd1 _1661_/A sky130_fd_sc_hd__nor2_8
X_1261_ _2325_/Q _2329_/Q _2333_/Q _2337_/Q _1275_/S0 _1065_/A vssd1 vssd1 vccd1 vccd1
+ _1261_/X sky130_fd_sc_hd__mux4_2
Xinput7 ram_addr[6] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__buf_6
XFILLER_49_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1192_ _1188_/X _1191_/X _1354_/A vssd1 vssd1 vccd1 vccd1 _1192_/X sky130_fd_sc_hd__o21ba_1
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1528_ _2131_/Q _1583_/A0 _1530_/S vssd1 vssd1 vccd1 vccd1 _2131_/D sky130_fd_sc_hd__mux2_1
XFILLER_19_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1459_ _1861_/A _1501_/A vssd1 vssd1 vccd1 vccd1 _1463_/S sky130_fd_sc_hd__nand2_2
XFILLER_74_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2431_ _2433_/CLK _2431_/D vssd1 vssd1 vccd1 vccd1 _2431_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2362_ _2368_/CLK _2362_/D vssd1 vssd1 vccd1 vccd1 _2362_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2293_ _2297_/CLK _2293_/D vssd1 vssd1 vccd1 vccd1 _2293_/Q sky130_fd_sc_hd__dfxtp_1
X_1313_ _1398_/A _1385_/B vssd1 vssd1 vccd1 vccd1 _1666_/A sky130_fd_sc_hd__or2_4
X_1244_ _1244_/A1 _1235_/Y _1237_/Y _1242_/Y _1243_/Y vssd1 vssd1 vccd1 vccd1 _1244_/X
+ sky130_fd_sc_hd__o32a_1
X_1175_ _2260_/Q _1988_/Q _1240_/S vssd1 vssd1 vccd1 vccd1 _1175_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_447 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1931_ _1931_/A _1976_/A vssd1 vssd1 vccd1 vccd1 _1935_/S sky130_fd_sc_hd__nand2_2
X_1862_ _1972_/A0 _2398_/Q _1865_/S vssd1 vssd1 vccd1 vccd1 _2398_/D sky130_fd_sc_hd__mux2_1
Xinput10 w_val[2] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__clkbuf_2
X_1793_ _2343_/Q _1793_/A1 _1795_/S vssd1 vssd1 vccd1 vccd1 _2343_/D sky130_fd_sc_hd__mux2_1
X_2414_ _2481_/CLK _2414_/D vssd1 vssd1 vccd1 vccd1 _2414_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2345_ _2497_/CLK _2345_/D vssd1 vssd1 vccd1 vccd1 _2345_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2276_ _2481_/CLK _2276_/D vssd1 vssd1 vccd1 vccd1 _2276_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1227_ _2052_/Q _2056_/Q _2060_/Q _2008_/Q _1303_/S0 _1304_/S1 vssd1 vssd1 vccd1
+ vccd1 _1227_/X sky130_fd_sc_hd__mux4_1
X_1158_ _2372_/Q _2376_/Q _2380_/Q _2020_/Q _1253_/S0 _1253_/S1 vssd1 vssd1 vccd1
+ vccd1 _1158_/X sky130_fd_sc_hd__mux4_1
XFILLER_37_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1089_ _2147_/Q _2151_/Q _2155_/Q _2159_/Q _1292_/S _1291_/A vssd1 vssd1 vccd1 vccd1
+ _1089_/X sky130_fd_sc_hd__mux4_1
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2130_ _2232_/CLK _2130_/D vssd1 vssd1 vccd1 vccd1 _2130_/Q sky130_fd_sc_hd__dfxtp_1
X_2061_ _2113_/CLK _2061_/D vssd1 vssd1 vccd1 vccd1 _2061_/Q sky130_fd_sc_hd__dfxtp_1
X_1012_ _1023_/B _1220_/A vssd1 vssd1 vccd1 vccd1 _1310_/A sky130_fd_sc_hd__nand2b_4
X_1914_ _2440_/Q _1974_/A0 _1915_/S vssd1 vssd1 vccd1 vccd1 _2440_/D sky130_fd_sc_hd__mux2_1
X_1845_ _2385_/Q _1845_/A1 _1845_/S vssd1 vssd1 vccd1 vccd1 _2385_/D sky130_fd_sc_hd__mux2_1
X_1776_ _1806_/A _1936_/B vssd1 vssd1 vccd1 vccd1 _1780_/S sky130_fd_sc_hd__or2_4
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2328_ _2329_/CLK _2328_/D vssd1 vssd1 vccd1 vccd1 _2328_/Q sky130_fd_sc_hd__dfxtp_1
X_2259_ _2261_/CLK _2259_/D vssd1 vssd1 vccd1 vccd1 _2259_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1630_ _2213_/Q _1660_/A0 _1630_/S vssd1 vssd1 vccd1 vccd1 _2213_/D sky130_fd_sc_hd__mux2_1
X_1561_ _1961_/A _1581_/A vssd1 vssd1 vccd1 vccd1 _1565_/S sky130_fd_sc_hd__nand2_4
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1492_ _2102_/Q _1982_/A1 _1495_/S vssd1 vssd1 vccd1 vccd1 _2102_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2113_ _2113_/CLK _2113_/D vssd1 vssd1 vccd1 vccd1 _2113_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2044_ _2496_/CLK _2044_/D vssd1 vssd1 vccd1 vccd1 _2044_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout29 _1011_/X vssd1 vssd1 vccd1 vccd1 _1298_/B2 sky130_fd_sc_hd__buf_8
XFILLER_62_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout18 _1470_/B vssd1 vssd1 vccd1 vccd1 _1486_/A sky130_fd_sc_hd__buf_12
X_1828_ _2371_/Q _1973_/A0 _1830_/S vssd1 vssd1 vccd1 vccd1 _2371_/D sky130_fd_sc_hd__mux2_1
X_1759_ _2316_/Q _1814_/A0 _1760_/S vssd1 vssd1 vccd1 vccd1 _2316_/D sky130_fd_sc_hd__mux2_1
XFILLER_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0992_ _0992_/A vssd1 vssd1 vccd1 vccd1 _0992_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1613_ _1823_/A0 _2199_/Q _1615_/S vssd1 vssd1 vccd1 vccd1 _2199_/D sky130_fd_sc_hd__mux2_1
X_1544_ _2144_/Q _1804_/A0 _1545_/S vssd1 vssd1 vccd1 vccd1 _2144_/D sky130_fd_sc_hd__mux2_1
X_1475_ _1475_/A _1475_/B _1475_/C vssd1 vssd1 vccd1 vccd1 _1956_/B sky130_fd_sc_hd__or3_4
XFILLER_39_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2027_ _2461_/CLK _2027_/D vssd1 vssd1 vccd1 vccd1 _2027_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1260_ _1037_/X _1259_/X _1251_/X vssd1 vssd1 vccd1 vccd1 _1260_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_83_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput8 w_val[0] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__clkbuf_4
X_1191_ _1409_/C _1189_/X _1190_/X _1305_/B2 vssd1 vssd1 vccd1 vccd1 _1191_/X sky130_fd_sc_hd__a22o_1
XFILLER_49_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1527_ _2130_/Q _1582_/A0 _1530_/S vssd1 vssd1 vccd1 vccd1 _2130_/D sky130_fd_sc_hd__mux2_1
X_1458_ _2077_/Q _1800_/A0 _1458_/S vssd1 vssd1 vccd1 vccd1 _2077_/D sky130_fd_sc_hd__mux2_1
X_1389_ _1969_/A0 _2028_/Q _1390_/S vssd1 vssd1 vccd1 vccd1 _2028_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2430_ _2433_/CLK _2430_/D vssd1 vssd1 vccd1 vccd1 _2430_/Q sky130_fd_sc_hd__dfxtp_1
X_2361_ _2369_/CLK _2361_/D vssd1 vssd1 vccd1 vccd1 _2361_/Q sky130_fd_sc_hd__dfxtp_1
X_2292_ _2296_/CLK _2292_/D vssd1 vssd1 vccd1 vccd1 _2292_/Q sky130_fd_sc_hd__dfxtp_1
X_1312_ _1398_/A _1385_/B vssd1 vssd1 vccd1 vccd1 _1736_/A sky130_fd_sc_hd__nor2_8
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1243_ _1180_/A _1238_/X _1024_/B vssd1 vssd1 vccd1 vccd1 _1243_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1174_ _1174_/A _1174_/B vssd1 vssd1 vccd1 vccd1 _1174_/X sky130_fd_sc_hd__and2_1
XFILLER_64_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1930_ _2453_/Q _1935_/A0 _1930_/S vssd1 vssd1 vccd1 vccd1 _2453_/D sky130_fd_sc_hd__mux2_1
X_1861_ _1861_/A _1901_/B vssd1 vssd1 vccd1 vccd1 _1865_/S sky130_fd_sc_hd__nand2_2
Xinput11 w_val[3] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__clkbuf_2
X_1792_ _2342_/Q _1792_/A1 _1795_/S vssd1 vssd1 vccd1 vccd1 _2342_/D sky130_fd_sc_hd__mux2_1
X_2413_ _2432_/CLK _2413_/D vssd1 vssd1 vccd1 vccd1 _2413_/Q sky130_fd_sc_hd__dfxtp_1
X_2344_ _2496_/CLK _2344_/D vssd1 vssd1 vccd1 vccd1 _2344_/Q sky130_fd_sc_hd__dfxtp_1
X_2275_ _2416_/CLK _2275_/D vssd1 vssd1 vccd1 vccd1 _2275_/Q sky130_fd_sc_hd__dfxtp_1
X_1226_ _2100_/Q _2016_/Q _2108_/Q _2112_/Q _1303_/S0 _1304_/S1 vssd1 vssd1 vccd1
+ vccd1 _1226_/X sky130_fd_sc_hd__mux4_1
XFILLER_25_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1157_ _1098_/X _1119_/X _1156_/X input7/X vssd1 vssd1 vccd1 vccd1 _1157_/Y sky130_fd_sc_hd__a22oi_4
X_1088_ _2115_/Q _2119_/Q _2123_/Q _2127_/Q _1297_/S0 _1297_/S1 vssd1 vssd1 vccd1
+ vccd1 _1088_/X sky130_fd_sc_hd__mux4_1
XFILLER_40_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2060_ _2113_/CLK _2060_/D vssd1 vssd1 vccd1 vccd1 _2060_/Q sky130_fd_sc_hd__dfxtp_1
X_1011_ _1244_/A1 _1237_/A vssd1 vssd1 vccd1 vccd1 _1011_/X sky130_fd_sc_hd__and2b_2
XFILLER_34_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1913_ _2439_/Q _1918_/A1 _1915_/S vssd1 vssd1 vccd1 vccd1 _2439_/D sky130_fd_sc_hd__mux2_1
X_1844_ _2384_/Q _1984_/A1 _1845_/S vssd1 vssd1 vccd1 vccd1 _2384_/D sky130_fd_sc_hd__mux2_1
X_1775_ _1985_/A1 _2329_/Q _1775_/S vssd1 vssd1 vccd1 vccd1 _2329_/D sky130_fd_sc_hd__mux2_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2327_ _2337_/CLK _2327_/D vssd1 vssd1 vccd1 vccd1 _2327_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2258_ _2261_/CLK _2258_/D vssd1 vssd1 vccd1 vccd1 _2258_/Q sky130_fd_sc_hd__dfxtp_1
X_1209_ _1453_/C _1208_/X _1385_/A vssd1 vssd1 vccd1 vccd1 _1209_/X sky130_fd_sc_hd__o21ba_1
XFILLER_25_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2189_ _2320_/CLK _2189_/D vssd1 vssd1 vccd1 vccd1 _2189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1560_ _2157_/Q _1980_/A0 _1560_/S vssd1 vssd1 vccd1 vccd1 _2157_/D sky130_fd_sc_hd__mux2_1
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1491_ _1981_/B _1916_/B vssd1 vssd1 vccd1 vccd1 _1495_/S sky130_fd_sc_hd__nor2_4
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2112_ _2363_/CLK _2112_/D vssd1 vssd1 vccd1 vccd1 _2112_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2043_ _2261_/CLK _2043_/D vssd1 vssd1 vccd1 vccd1 _2043_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout19 _1531_/B vssd1 vssd1 vccd1 vccd1 _1566_/A sky130_fd_sc_hd__buf_12
XFILLER_50_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1827_ _2370_/Q _1972_/A0 _1830_/S vssd1 vssd1 vccd1 vccd1 _2370_/D sky130_fd_sc_hd__mux2_1
X_1758_ _2315_/Q _1823_/A0 _1760_/S vssd1 vssd1 vccd1 vccd1 _2315_/D sky130_fd_sc_hd__mux2_1
X_1689_ _2260_/Q _1739_/A0 _1690_/S vssd1 vssd1 vccd1 vccd1 _2260_/D sky130_fd_sc_hd__mux2_1
XFILLER_38_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0991_ input7/X vssd1 vssd1 vccd1 vccd1 _1048_/A sky130_fd_sc_hd__inv_2
X_1612_ _1917_/A1 _2198_/Q _1615_/S vssd1 vssd1 vccd1 vccd1 _2198_/D sky130_fd_sc_hd__mux2_1
XFILLER_5_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1543_ _2143_/Q _1783_/A0 _1545_/S vssd1 vssd1 vccd1 vccd1 _2143_/D sky130_fd_sc_hd__mux2_1
XFILLER_5_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1474_ _2089_/Q _1800_/A0 _1474_/S vssd1 vssd1 vccd1 vccd1 _2089_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2026_ _2457_/CLK _2026_/D vssd1 vssd1 vccd1 vccd1 _2026_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1190_ _2308_/Q _2312_/Q _2316_/Q _2320_/Q _1285_/S0 _1285_/S1 vssd1 vssd1 vccd1
+ vccd1 _1190_/X sky130_fd_sc_hd__mux4_2
XFILLER_76_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput9 w_val[1] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__buf_2
XFILLER_32_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1526_ _1566_/A _1926_/B vssd1 vssd1 vccd1 vccd1 _1530_/S sky130_fd_sc_hd__nor2_4
X_1457_ _2076_/Q _1809_/A0 _1458_/S vssd1 vssd1 vccd1 vccd1 _2076_/D sky130_fd_sc_hd__mux2_1
X_1388_ _1963_/A0 _2027_/Q _1390_/S vssd1 vssd1 vccd1 vccd1 _2027_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2009_ _2113_/CLK _2009_/D vssd1 vssd1 vccd1 vccd1 _2009_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2360_ _2368_/CLK _2360_/D vssd1 vssd1 vccd1 vccd1 _2360_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2291_ _2296_/CLK _2291_/D vssd1 vssd1 vccd1 vccd1 _2291_/Q sky130_fd_sc_hd__dfxtp_1
X_1311_ input7/X _1329_/B vssd1 vssd1 vccd1 vccd1 _1385_/B sky130_fd_sc_hd__nand2_8
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1242_ _1174_/A _1240_/X _1241_/X vssd1 vssd1 vccd1 vccd1 _1242_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_49_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1173_ _2268_/Q _2272_/Q _1240_/S vssd1 vssd1 vccd1 vccd1 _1174_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_44_clk clkbuf_leaf_4_clk/A vssd1 vssd1 vccd1 vccd1 _2177_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_20_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1509_ _2116_/Q _1974_/A0 _1510_/S vssd1 vssd1 vccd1 vccd1 _2116_/D sky130_fd_sc_hd__mux2_1
X_2489_ _2493_/CLK _2489_/D vssd1 vssd1 vccd1 vccd1 _2489_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_35_clk clkbuf_2_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _2485_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_51_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_26_clk clkbuf_2_3__f_clk/X vssd1 vssd1 vccd1 vccd1 _2301_/CLK sky130_fd_sc_hd__clkbuf_16
X_1860_ _1975_/A0 _2397_/Q _1860_/S vssd1 vssd1 vccd1 vccd1 _2397_/D sky130_fd_sc_hd__mux2_1
Xinput12 wen vssd1 vssd1 vccd1 vccd1 _1329_/B sky130_fd_sc_hd__buf_4
X_1791_ _1981_/B _1946_/B vssd1 vssd1 vccd1 vccd1 _1795_/S sky130_fd_sc_hd__nor2_2
XFILLER_6_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2412_ _2416_/CLK _2412_/D vssd1 vssd1 vccd1 vccd1 _2412_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2343_ _2343_/CLK _2343_/D vssd1 vssd1 vccd1 vccd1 _2343_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2274_ _2296_/CLK _2274_/D vssd1 vssd1 vccd1 vccd1 _2274_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1225_ _1302_/A1 _1223_/X _1224_/X _1020_/X vssd1 vssd1 vccd1 vccd1 _1225_/X sky130_fd_sc_hd__a22o_1
XFILLER_37_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1156_ _1398_/A _1132_/X _1155_/Y _1354_/A _1148_/Y vssd1 vssd1 vccd1 vccd1 _1156_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1087_ _2131_/Q _2135_/Q _2139_/Q _2003_/Q _1297_/S0 _1297_/S1 vssd1 vssd1 vccd1
+ vccd1 _1087_/X sky130_fd_sc_hd__mux4_2
Xclkbuf_leaf_17_clk clkbuf_2_3__f_clk/X vssd1 vssd1 vccd1 vccd1 _2495_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_33_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1989_ _2297_/CLK _1989_/D vssd1 vssd1 vccd1 vccd1 _1989_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1010_ _1040_/B input6/X vssd1 vssd1 vccd1 vccd1 _1385_/A sky130_fd_sc_hd__nand2_8
XFILLER_19_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1912_ _2438_/Q _1917_/A1 _1915_/S vssd1 vssd1 vccd1 vccd1 _2438_/D sky130_fd_sc_hd__mux2_1
X_1843_ _2383_/Q _1843_/A1 _1845_/S vssd1 vssd1 vccd1 vccd1 _2383_/D sky130_fd_sc_hd__mux2_1
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1774_ _1944_/A0 _2328_/Q _1775_/S vssd1 vssd1 vccd1 vccd1 _2328_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_6_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _2320_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_69_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2326_ _2337_/CLK _2326_/D vssd1 vssd1 vccd1 vccd1 _2326_/Q sky130_fd_sc_hd__dfxtp_1
X_2257_ _2343_/CLK _2257_/D vssd1 vssd1 vccd1 vccd1 _2257_/Q sky130_fd_sc_hd__dfxtp_1
X_1208_ _2196_/Q _2200_/Q _2204_/Q _2208_/Q _1453_/A _1283_/S1 vssd1 vssd1 vccd1 vccd1
+ _1208_/X sky130_fd_sc_hd__mux4_1
XFILLER_72_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2188_ _2320_/CLK _2188_/D vssd1 vssd1 vccd1 vccd1 _2188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1139_ _1420_/C _1135_/X _1138_/X _1134_/X vssd1 vssd1 vccd1 vccd1 _1139_/X sky130_fd_sc_hd__o211a_1
XFILLER_21_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1490_ _2101_/Q _1505_/A0 _1490_/S vssd1 vssd1 vccd1 vccd1 _2101_/D sky130_fd_sc_hd__mux2_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2111_ _2113_/CLK _2111_/D vssd1 vssd1 vccd1 vccd1 _2111_/Q sky130_fd_sc_hd__dfxtp_1
X_2042_ _2261_/CLK _2042_/D vssd1 vssd1 vccd1 vccd1 _2042_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1826_ _1886_/A _1906_/B vssd1 vssd1 vccd1 vccd1 _1830_/S sky130_fd_sc_hd__nor2_2
X_1757_ _2314_/Q _1762_/A0 _1760_/S vssd1 vssd1 vccd1 vccd1 _2314_/D sky130_fd_sc_hd__mux2_1
X_1688_ _2259_/Q _1793_/A1 _1690_/S vssd1 vssd1 vccd1 vccd1 _2259_/D sky130_fd_sc_hd__mux2_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2309_ _2363_/CLK _2309_/D vssd1 vssd1 vccd1 vccd1 _2309_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1611_ _1931_/A _1661_/A vssd1 vssd1 vccd1 vccd1 _1615_/S sky130_fd_sc_hd__nand2_2
X_1542_ _2142_/Q _1842_/A1 _1545_/S vssd1 vssd1 vccd1 vccd1 _2142_/D sky130_fd_sc_hd__mux2_1
X_1473_ _2088_/Q _1784_/A0 _1474_/S vssd1 vssd1 vccd1 vccd1 _2088_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2025_ _2433_/CLK _2025_/D vssd1 vssd1 vccd1 vccd1 _2025_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1809_ _1809_/A0 _2356_/Q _1810_/S vssd1 vssd1 vccd1 vccd1 _2356_/D sky130_fd_sc_hd__mux2_1
XFILLER_77_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1525_ _2129_/Q _1585_/A0 _1525_/S vssd1 vssd1 vccd1 vccd1 _2129_/D sky130_fd_sc_hd__mux2_1
X_1456_ _2075_/Q _1778_/A0 _1458_/S vssd1 vssd1 vccd1 vccd1 _2075_/D sky130_fd_sc_hd__mux2_1
X_1387_ _1972_/A0 _2026_/Q _1390_/S vssd1 vssd1 vccd1 vccd1 _2026_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2008_ _2113_/CLK _2008_/D vssd1 vssd1 vccd1 vccd1 _2008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1310_ _1310_/A _1366_/A vssd1 vssd1 vccd1 vccd1 _1641_/A sky130_fd_sc_hd__or2_4
X_2290_ _2301_/CLK _2290_/D vssd1 vssd1 vccd1 vccd1 _2290_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1241_ _1475_/B _1239_/X _1241_/B1 vssd1 vssd1 vccd1 vccd1 _1241_/X sky130_fd_sc_hd__a21o_1
XFILLER_2_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1172_ _1040_/B _1162_/X _1164_/X _1171_/X input6/X vssd1 vssd1 vccd1 vccd1 _1172_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_49_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1508_ _2115_/Q _1918_/A1 _1510_/S vssd1 vssd1 vccd1 vccd1 _2115_/D sky130_fd_sc_hd__mux2_1
X_2488_ _2493_/CLK _2488_/D vssd1 vssd1 vccd1 vccd1 _2488_/Q sky130_fd_sc_hd__dfxtp_1
X_1439_ _2063_/Q _1783_/A0 _1441_/S vssd1 vssd1 vccd1 vccd1 _2063_/D sky130_fd_sc_hd__mux2_1
XFILLER_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1790_ _2341_/Q _1985_/A1 _1790_/S vssd1 vssd1 vccd1 vccd1 _2341_/D sky130_fd_sc_hd__mux2_1
X_2411_ _2432_/CLK _2411_/D vssd1 vssd1 vccd1 vccd1 _2411_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2342_ _2497_/CLK _2342_/D vssd1 vssd1 vccd1 vccd1 _2342_/Q sky130_fd_sc_hd__dfxtp_1
X_2273_ _2297_/CLK _2273_/D vssd1 vssd1 vccd1 vccd1 _2273_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1224_ _2084_/Q _2088_/Q _2092_/Q _2096_/Q _1303_/S0 _1301_/S1 vssd1 vssd1 vccd1
+ vccd1 _1224_/X sky130_fd_sc_hd__mux4_1
XFILLER_80_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1155_ _1155_/A _1155_/B vssd1 vssd1 vccd1 vccd1 _1155_/Y sky130_fd_sc_hd__nor2_1
X_1086_ _2163_/Q _2167_/Q _2171_/Q _2175_/Q _1297_/S0 _1297_/S1 vssd1 vssd1 vccd1
+ vccd1 _1086_/X sky130_fd_sc_hd__mux4_1
XFILLER_25_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1988_ _2301_/CLK _1988_/D vssd1 vssd1 vccd1 vccd1 _1988_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_2__f_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_2__f_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_16_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1911_ _1911_/A _1966_/A vssd1 vssd1 vccd1 vccd1 _1915_/S sky130_fd_sc_hd__nor2_2
X_1842_ _2382_/Q _1842_/A1 _1845_/S vssd1 vssd1 vccd1 vccd1 _2382_/D sky130_fd_sc_hd__mux2_1
XFILLER_8_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1773_ _1783_/A0 _2327_/Q _1775_/S vssd1 vssd1 vccd1 vccd1 _2327_/D sky130_fd_sc_hd__mux2_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2325_ _2385_/CLK _2325_/D vssd1 vssd1 vccd1 vccd1 _2325_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2256_ _2480_/CLK _2256_/D vssd1 vssd1 vccd1 vccd1 _2256_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1207_ _1398_/A _1207_/B vssd1 vssd1 vccd1 vccd1 _1207_/Y sky130_fd_sc_hd__nor2_1
XFILLER_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2187_ _2241_/CLK _2187_/D vssd1 vssd1 vccd1 vccd1 _2187_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1138_ _1464_/C _1136_/X _1137_/X _1396_/C vssd1 vssd1 vccd1 vccd1 _1138_/X sky130_fd_sc_hd__o22a_1
XFILLER_40_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1069_ _1237_/A _1068_/X _1244_/A1 vssd1 vssd1 vccd1 vccd1 _1069_/X sky130_fd_sc_hd__o21ba_1
XFILLER_80_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2110_ _2367_/CLK _2110_/D vssd1 vssd1 vccd1 vccd1 _2110_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2041_ _2049_/CLK _2041_/D vssd1 vssd1 vccd1 vccd1 _2041_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1825_ _1940_/A0 _2369_/Q _1825_/S vssd1 vssd1 vccd1 vccd1 _2369_/D sky130_fd_sc_hd__mux2_1
X_1756_ _1806_/A _1916_/B vssd1 vssd1 vccd1 vccd1 _1760_/S sky130_fd_sc_hd__nor2_4
X_1687_ _2258_/Q _1792_/A1 _1690_/S vssd1 vssd1 vccd1 vccd1 _2258_/D sky130_fd_sc_hd__mux2_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2308_ _2320_/CLK _2308_/D vssd1 vssd1 vccd1 vccd1 _2308_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2239_ _2240_/CLK _2239_/D vssd1 vssd1 vccd1 vccd1 _2239_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1610_ _2197_/Q _1765_/A0 _1610_/S vssd1 vssd1 vccd1 vccd1 _2197_/D sky130_fd_sc_hd__mux2_1
XFILLER_5_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1541_ _1681_/B _1981_/B vssd1 vssd1 vccd1 vccd1 _1545_/S sky130_fd_sc_hd__nor2_2
X_1472_ _2087_/Q _1778_/A0 _1474_/S vssd1 vssd1 vccd1 vccd1 _2087_/D sky130_fd_sc_hd__mux2_1
XFILLER_5_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_76 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2024_ _2421_/CLK _2024_/D vssd1 vssd1 vccd1 vccd1 _2024_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1808_ _1808_/A0 _2355_/Q _1810_/S vssd1 vssd1 vccd1 vccd1 _2355_/D sky130_fd_sc_hd__mux2_1
XFILLER_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1739_ _1739_/A0 _2300_/Q _1740_/S vssd1 vssd1 vccd1 vccd1 _2300_/D sky130_fd_sc_hd__mux2_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1524_ _2128_/Q _1579_/A0 _1525_/S vssd1 vssd1 vccd1 vccd1 _2128_/D sky130_fd_sc_hd__mux2_1
X_1455_ _2074_/Q _1822_/A0 _1458_/S vssd1 vssd1 vccd1 vccd1 _2074_/D sky130_fd_sc_hd__mux2_1
X_1386_ _1861_/A _1976_/A vssd1 vssd1 vccd1 vccd1 _1390_/S sky130_fd_sc_hd__nand2_2
XFILLER_67_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2007_ _2094_/CLK _2007_/D vssd1 vssd1 vccd1 vccd1 _2007_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1240_ _2301_/Q _2013_/Q _1240_/S vssd1 vssd1 vccd1 vccd1 _1240_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1171_ _1167_/X _1170_/X _1040_/B vssd1 vssd1 vccd1 vccd1 _1171_/X sky130_fd_sc_hd__a21bo_1
XFILLER_52_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2487_ _2493_/CLK _2487_/D vssd1 vssd1 vccd1 vccd1 _2487_/Q sky130_fd_sc_hd__dfxtp_1
X_1507_ _2114_/Q _1977_/A0 _1510_/S vssd1 vssd1 vccd1 vccd1 _2114_/D sky130_fd_sc_hd__mux2_1
X_1438_ _2062_/Q _1982_/A1 _1441_/S vssd1 vssd1 vccd1 vccd1 _2062_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1369_ _1503_/A0 _2015_/Q _1371_/S vssd1 vssd1 vccd1 vccd1 _2015_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2410_ _2481_/CLK _2410_/D vssd1 vssd1 vccd1 vccd1 _2410_/Q sky130_fd_sc_hd__dfxtp_1
X_2341_ _2497_/CLK _2341_/D vssd1 vssd1 vccd1 vccd1 _2341_/Q sky130_fd_sc_hd__dfxtp_1
X_2272_ _2301_/CLK _2272_/D vssd1 vssd1 vccd1 vccd1 _2272_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1223_ _2068_/Q _2072_/Q _2076_/Q _2080_/Q _1304_/S0 _1301_/S1 vssd1 vssd1 vccd1
+ vccd1 _1223_/X sky130_fd_sc_hd__mux4_1
XFILLER_84_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1154_ _1409_/C _1152_/X _1153_/X _1305_/B2 vssd1 vssd1 vccd1 vccd1 _1155_/B sky130_fd_sc_hd__a22o_1
XFILLER_80_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1085_ _1009_/Y _1048_/X _1084_/X input7/X vssd1 vssd1 vccd1 vccd1 _1085_/X sky130_fd_sc_hd__o22a_2
XFILLER_33_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1987_ _2297_/CLK _1987_/D vssd1 vssd1 vccd1 vccd1 _1987_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_451 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1910_ _2437_/Q _1975_/A0 _1910_/S vssd1 vssd1 vccd1 vccd1 _2437_/D sky130_fd_sc_hd__mux2_1
XFILLER_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1841_ _1981_/B _1906_/B vssd1 vssd1 vccd1 vccd1 _1845_/S sky130_fd_sc_hd__nor2_4
XFILLER_30_443 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1772_ _1842_/A1 _2326_/Q _1775_/S vssd1 vssd1 vccd1 vccd1 _2326_/D sky130_fd_sc_hd__mux2_1
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2324_ _2329_/CLK _2324_/D vssd1 vssd1 vccd1 vccd1 _2324_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2255_ _2480_/CLK _2255_/D vssd1 vssd1 vccd1 vccd1 _2255_/Q sky130_fd_sc_hd__dfxtp_1
X_2186_ _2241_/CLK _2186_/D vssd1 vssd1 vccd1 vccd1 _2186_/Q sky130_fd_sc_hd__dfxtp_1
X_1206_ _1023_/B _1197_/Y _1199_/Y _1204_/Y _1205_/Y vssd1 vssd1 vccd1 vccd1 _1207_/B
+ sky130_fd_sc_hd__o32a_2
X_1137_ _2483_/Q _2487_/Q _2491_/Q _2031_/Q _1253_/S0 _1253_/S1 vssd1 vssd1 vccd1
+ vccd1 _1137_/X sky130_fd_sc_hd__mux4_2
XFILLER_65_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1068_ _2382_/Q _2062_/Q _2102_/Q _2142_/Q _1275_/S0 _1065_/A vssd1 vssd1 vccd1 vccd1
+ _1068_/X sky130_fd_sc_hd__mux4_1
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2040_ _2049_/CLK _2040_/D vssd1 vssd1 vccd1 vccd1 _2040_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1824_ _1824_/A0 _2368_/Q _1825_/S vssd1 vssd1 vccd1 vccd1 _2368_/D sky130_fd_sc_hd__mux2_1
X_1755_ _2313_/Q _1765_/A0 _1755_/S vssd1 vssd1 vccd1 vccd1 _2313_/D sky130_fd_sc_hd__mux2_1
X_1686_ _1726_/A _1926_/B vssd1 vssd1 vccd1 vccd1 _1690_/S sky130_fd_sc_hd__nor2_2
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2307_ _2320_/CLK _2307_/D vssd1 vssd1 vccd1 vccd1 _2307_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2238_ _2240_/CLK _2238_/D vssd1 vssd1 vccd1 vccd1 _2238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2169_ _2176_/CLK _2169_/D vssd1 vssd1 vccd1 vccd1 _2169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1540_ _2141_/Q _1585_/A0 _1540_/S vssd1 vssd1 vccd1 vccd1 _2141_/D sky130_fd_sc_hd__mux2_1
X_1471_ _2086_/Q _1777_/A0 _1474_/S vssd1 vssd1 vccd1 vccd1 _2086_/D sky130_fd_sc_hd__mux2_1
XFILLER_5_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2023_ _2421_/CLK _2023_/D vssd1 vssd1 vccd1 vccd1 _2023_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1807_ _1822_/A0 _2354_/Q _1810_/S vssd1 vssd1 vccd1 vccd1 _2354_/D sky130_fd_sc_hd__mux2_1
X_1738_ _1738_/A0 _2299_/Q _1740_/S vssd1 vssd1 vccd1 vccd1 _2299_/D sky130_fd_sc_hd__mux2_1
X_1669_ _2244_/Q _1804_/A0 _1670_/S vssd1 vssd1 vccd1 vccd1 _2244_/D sky130_fd_sc_hd__mux2_1
XFILLER_49_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1523_ _2127_/Q _1583_/A0 _1525_/S vssd1 vssd1 vccd1 vccd1 _2127_/D sky130_fd_sc_hd__mux2_1
X_1454_ _1486_/A _1936_/B vssd1 vssd1 vccd1 vccd1 _1458_/S sky130_fd_sc_hd__nor2_2
X_1385_ _1385_/A _1385_/B vssd1 vssd1 vccd1 vccd1 _1966_/A sky130_fd_sc_hd__or2_4
XFILLER_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2006_ _2094_/CLK _2006_/D vssd1 vssd1 vccd1 vccd1 _2006_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_38_clk clkbuf_2_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _2479_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1170_ _1396_/C _1168_/X _1169_/X _1420_/C vssd1 vssd1 vccd1 vccd1 _1170_/X sky130_fd_sc_hd__o22a_1
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_29_clk clkbuf_2_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _2481_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_64_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2486_ _2493_/CLK _2486_/D vssd1 vssd1 vccd1 vccd1 _2486_/Q sky130_fd_sc_hd__dfxtp_1
X_1506_ _1566_/A _1906_/B vssd1 vssd1 vccd1 vccd1 _1510_/S sky130_fd_sc_hd__nor2_2
X_1437_ _1911_/A _1981_/B vssd1 vssd1 vccd1 vccd1 _1441_/S sky130_fd_sc_hd__nor2_4
X_1368_ _1762_/A0 _2014_/Q _1371_/S vssd1 vssd1 vccd1 vccd1 _2014_/D sky130_fd_sc_hd__mux2_1
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1299_ _1295_/X _1298_/X _1037_/X vssd1 vssd1 vccd1 vccd1 _1307_/C sky130_fd_sc_hd__o21a_1
XFILLER_23_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2340_ _2495_/CLK _2340_/D vssd1 vssd1 vccd1 vccd1 _2340_/Q sky130_fd_sc_hd__dfxtp_1
X_2271_ _2297_/CLK _2271_/D vssd1 vssd1 vccd1 vccd1 _2271_/Q sky130_fd_sc_hd__dfxtp_1
X_1222_ _1217_/X _1221_/X _1037_/X vssd1 vssd1 vccd1 vccd1 _1230_/C sky130_fd_sc_hd__o21a_1
XFILLER_77_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1153_ _2307_/Q _2311_/Q _2315_/Q _2319_/Q _1285_/S0 _1285_/S1 vssd1 vssd1 vccd1
+ vccd1 _1153_/X sky130_fd_sc_hd__mux4_2
XFILLER_80_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1084_ _0994_/Y _1076_/X _1083_/X _1063_/X vssd1 vssd1 vccd1 vccd1 _1084_/X sky130_fd_sc_hd__a211o_1
XFILLER_33_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1986_ _2261_/CLK _1986_/D vssd1 vssd1 vccd1 vccd1 _1986_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_9_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _2113_/CLK sky130_fd_sc_hd__clkbuf_16
X_2469_ _2481_/CLK _2469_/D vssd1 vssd1 vccd1 vccd1 _2469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1840_ _2381_/Q _1975_/A0 _1840_/S vssd1 vssd1 vccd1 vccd1 _2381_/D sky130_fd_sc_hd__mux2_1
XFILLER_30_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1771_ _1931_/A _1821_/A vssd1 vssd1 vccd1 vccd1 _1775_/S sky130_fd_sc_hd__nand2_4
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2323_ _2385_/CLK _2323_/D vssd1 vssd1 vccd1 vccd1 _2323_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2254_ _2457_/CLK _2254_/D vssd1 vssd1 vccd1 vccd1 _2254_/Q sky130_fd_sc_hd__dfxtp_1
X_2185_ _2302_/CLK _2185_/D vssd1 vssd1 vccd1 vccd1 _2185_/Q sky130_fd_sc_hd__dfxtp_1
X_1205_ _1237_/A _1200_/X _1023_/B vssd1 vssd1 vccd1 vccd1 _1205_/Y sky130_fd_sc_hd__o21ai_1
X_1136_ _2467_/Q _2471_/Q _2475_/Q _2479_/Q _1475_/A _1464_/B vssd1 vssd1 vccd1 vccd1
+ _1136_/X sky130_fd_sc_hd__mux4_1
XFILLER_53_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1067_ _1234_/A1 _1066_/X _1065_/X _1241_/B1 vssd1 vssd1 vccd1 vccd1 _1067_/X sky130_fd_sc_hd__a211o_1
X_1969_ _1969_/A0 _2484_/Q _1970_/S vssd1 vssd1 vccd1 vccd1 _2484_/D sky130_fd_sc_hd__mux2_1
XFILLER_4_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1823_ _1823_/A0 _2367_/Q _1825_/S vssd1 vssd1 vccd1 vccd1 _2367_/D sky130_fd_sc_hd__mux2_1
X_1754_ _2312_/Q _1814_/A0 _1755_/S vssd1 vssd1 vccd1 vccd1 _2312_/D sky130_fd_sc_hd__mux2_1
X_1685_ _2257_/Q _1935_/A0 _1685_/S vssd1 vssd1 vccd1 vccd1 _2257_/D sky130_fd_sc_hd__mux2_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2306_ _2368_/CLK _2306_/D vssd1 vssd1 vccd1 vccd1 _2306_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2237_ _2241_/CLK _2237_/D vssd1 vssd1 vccd1 vccd1 _2237_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2168_ _2176_/CLK _2168_/D vssd1 vssd1 vccd1 vccd1 _2168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1119_ _1398_/A _1111_/X _1118_/Y _1354_/A _1048_/A vssd1 vssd1 vccd1 vccd1 _1119_/X
+ sky130_fd_sc_hd__o221a_2
X_2099_ _2367_/CLK _2099_/D vssd1 vssd1 vccd1 vccd1 _2099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_447 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1470_ _1981_/A _1470_/B vssd1 vssd1 vccd1 vccd1 _1474_/S sky130_fd_sc_hd__nor2_4
XFILLER_79_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2022_ _2432_/CLK _2022_/D vssd1 vssd1 vccd1 vccd1 _2022_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1806_ _1806_/A _1966_/B vssd1 vssd1 vccd1 vccd1 _1810_/S sky130_fd_sc_hd__or2_4
X_1737_ _1792_/A1 _2298_/Q _1740_/S vssd1 vssd1 vccd1 vccd1 _2298_/D sky130_fd_sc_hd__mux2_1
X_1668_ _2243_/Q _1793_/A1 _1670_/S vssd1 vssd1 vccd1 vccd1 _2243_/D sky130_fd_sc_hd__mux2_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1599_ _2188_/Q _1814_/A0 _1600_/S vssd1 vssd1 vccd1 vccd1 _2188_/D sky130_fd_sc_hd__mux2_1
XFILLER_85_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1522_ _2126_/Q _1662_/A0 _1525_/S vssd1 vssd1 vccd1 vccd1 _2126_/D sky130_fd_sc_hd__mux2_1
X_1453_ _1453_/A _1475_/B _1453_/C vssd1 vssd1 vccd1 vccd1 _1936_/B sky130_fd_sc_hd__or3_4
X_1384_ _1385_/A _1385_/B vssd1 vssd1 vccd1 vccd1 _1976_/A sky130_fd_sc_hd__nor2_8
X_2005_ _2240_/CLK _2005_/D vssd1 vssd1 vccd1 vccd1 _2005_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1505_ _1505_/A0 _2113_/Q _1505_/S vssd1 vssd1 vccd1 vccd1 _2113_/D sky130_fd_sc_hd__mux2_1
X_2485_ _2485_/CLK _2485_/D vssd1 vssd1 vccd1 vccd1 _2485_/Q sky130_fd_sc_hd__dfxtp_1
X_1436_ _2061_/Q _1505_/A0 _1436_/S vssd1 vssd1 vccd1 vccd1 _2061_/D sky130_fd_sc_hd__mux2_1
X_1367_ _1501_/A _1971_/A vssd1 vssd1 vccd1 vccd1 _1371_/S sky130_fd_sc_hd__nand2_4
XFILLER_28_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1298_ _1409_/C _1296_/X _1297_/X _1298_/B2 vssd1 vssd1 vccd1 vccd1 _1298_/X sky130_fd_sc_hd__a22o_1
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2270_ _2343_/CLK _2270_/D vssd1 vssd1 vccd1 vccd1 _2270_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1221_ _1258_/A _1218_/X _1220_/X _1024_/B vssd1 vssd1 vccd1 vccd1 _1221_/X sky130_fd_sc_hd__o211a_1
XFILLER_77_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1152_ _2355_/Q _2359_/Q _2363_/Q _2367_/Q _1285_/S0 _1285_/S1 vssd1 vssd1 vccd1
+ vccd1 _1152_/X sky130_fd_sc_hd__mux4_1
XFILLER_18_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1083_ _1079_/X _1082_/X _1354_/A vssd1 vssd1 vccd1 vccd1 _1083_/X sky130_fd_sc_hd__o21ba_1
XFILLER_60_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1985_ _2497_/Q _1985_/A1 _1985_/S vssd1 vssd1 vccd1 vccd1 _2497_/D sky130_fd_sc_hd__mux2_1
X_2468_ _2480_/CLK _2468_/D vssd1 vssd1 vccd1 vccd1 _2468_/Q sky130_fd_sc_hd__dfxtp_1
X_1419_ _2049_/Q _1845_/A1 _1419_/S vssd1 vssd1 vccd1 vccd1 _2049_/D sky130_fd_sc_hd__mux2_1
X_2399_ _2485_/CLK _2399_/D vssd1 vssd1 vccd1 vccd1 _2399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1770_ _2325_/Q _1985_/A1 _1770_/S vssd1 vssd1 vccd1 vccd1 _2325_/D sky130_fd_sc_hd__mux2_1
XFILLER_8_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2322_ _2329_/CLK _2322_/D vssd1 vssd1 vccd1 vccd1 _2322_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2253_ _2343_/CLK _2253_/D vssd1 vssd1 vccd1 vccd1 _2253_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1204_ _1100_/A _1202_/X _1203_/X vssd1 vssd1 vccd1 vccd1 _1204_/Y sky130_fd_sc_hd__a21oi_1
X_2184_ _2302_/CLK _2184_/D vssd1 vssd1 vccd1 vccd1 _2184_/Q sky130_fd_sc_hd__dfxtp_1
X_1135_ _2435_/Q _2439_/Q _2443_/Q _2447_/Q _1292_/S _1253_/S1 vssd1 vssd1 vccd1 vccd1
+ _1135_/X sky130_fd_sc_hd__mux4_1
XFILLER_65_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1066_ _2182_/Q _2222_/Q _1277_/S vssd1 vssd1 vccd1 vccd1 _1066_/X sky130_fd_sc_hd__mux2_1
X_1968_ _1973_/A0 _2483_/Q _1970_/S vssd1 vssd1 vccd1 vccd1 _2483_/D sky130_fd_sc_hd__mux2_1
X_1899_ _1904_/A0 _2428_/Q _1900_/S vssd1 vssd1 vccd1 vccd1 _2428_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1822_ _1822_/A0 _2366_/Q _1825_/S vssd1 vssd1 vccd1 vccd1 _2366_/D sky130_fd_sc_hd__mux2_1
XFILLER_30_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1753_ _2311_/Q _1823_/A0 _1755_/S vssd1 vssd1 vccd1 vccd1 _2311_/D sky130_fd_sc_hd__mux2_1
X_1684_ _2256_/Q _1804_/A0 _1685_/S vssd1 vssd1 vccd1 vccd1 _2256_/D sky130_fd_sc_hd__mux2_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2305_ _2496_/CLK _2305_/D vssd1 vssd1 vccd1 vccd1 _2305_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2236_ _2240_/CLK _2236_/D vssd1 vssd1 vccd1 vccd1 _2236_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2167_ _2176_/CLK _2167_/D vssd1 vssd1 vccd1 vccd1 _2167_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2098_ _2367_/CLK _2098_/D vssd1 vssd1 vccd1 vccd1 _2098_/Q sky130_fd_sc_hd__dfxtp_1
X_1118_ _1118_/A _1118_/B vssd1 vssd1 vccd1 vccd1 _1118_/Y sky130_fd_sc_hd__nor2_1
XFILLER_80_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1049_ _2114_/Q _2118_/Q _2122_/Q _2126_/Q _1287_/S0 _1013_/B vssd1 vssd1 vccd1 vccd1
+ _1049_/X sky130_fd_sc_hd__mux4_1
XFILLER_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2021_ _2482_/CLK _2021_/D vssd1 vssd1 vccd1 vccd1 _2021_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1805_ _1940_/A0 _2353_/Q _1805_/S vssd1 vssd1 vccd1 vccd1 _2353_/D sky130_fd_sc_hd__mux2_1
X_1736_ _1736_/A _1976_/B vssd1 vssd1 vccd1 vccd1 _1740_/S sky130_fd_sc_hd__nand2_2
XFILLER_49_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1667_ _2242_/Q _1982_/A1 _1670_/S vssd1 vssd1 vccd1 vccd1 _2242_/D sky130_fd_sc_hd__mux2_1
X_1598_ _2187_/Q _1663_/A0 _1600_/S vssd1 vssd1 vccd1 vccd1 _2187_/D sky130_fd_sc_hd__mux2_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2219_ _2229_/CLK _2219_/D vssd1 vssd1 vccd1 vccd1 _2219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1521_ _1566_/A _1681_/B vssd1 vssd1 vccd1 vccd1 _1525_/S sky130_fd_sc_hd__nor2_2
X_1452_ _2073_/Q _1800_/A0 _1452_/S vssd1 vssd1 vccd1 vccd1 _2073_/D sky130_fd_sc_hd__mux2_1
X_1383_ _1975_/A0 _2025_/Q _1383_/S vssd1 vssd1 vccd1 vccd1 _2025_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2004_ _2232_/CLK _2004_/D vssd1 vssd1 vccd1 vccd1 _2004_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1719_ _2284_/Q _1904_/A0 _1720_/S vssd1 vssd1 vccd1 vccd1 _2284_/D sky130_fd_sc_hd__mux2_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1504_ _1784_/A0 _2112_/Q _1505_/S vssd1 vssd1 vccd1 vccd1 _2112_/D sky130_fd_sc_hd__mux2_1
X_2484_ _2485_/CLK _2484_/D vssd1 vssd1 vccd1 vccd1 _2484_/Q sky130_fd_sc_hd__dfxtp_1
X_1435_ _2060_/Q _1824_/A0 _1436_/S vssd1 vssd1 vccd1 vccd1 _2060_/D sky130_fd_sc_hd__mux2_1
X_1366_ _1366_/A _1396_/C vssd1 vssd1 vccd1 vccd1 _1971_/A sky130_fd_sc_hd__nor2_8
X_1297_ _2133_/Q _2137_/Q _2141_/Q _2005_/Q _1297_/S0 _1297_/S1 vssd1 vssd1 vccd1
+ vccd1 _1297_/X sky130_fd_sc_hd__mux4_1
XFILLER_36_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1220_ _1220_/A _1220_/B vssd1 vssd1 vccd1 vccd1 _1220_/X sky130_fd_sc_hd__or2_1
X_1151_ _1302_/A1 _1149_/X _1150_/X _1020_/X vssd1 vssd1 vccd1 vccd1 _1155_/A sky130_fd_sc_hd__a22o_1
X_1082_ _1409_/C _1080_/X _1081_/X _1295_/B2 vssd1 vssd1 vccd1 vccd1 _1082_/X sky130_fd_sc_hd__a22o_1
XFILLER_18_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1984_ _2496_/Q _1984_/A1 _1985_/S vssd1 vssd1 vccd1 vccd1 _2496_/D sky130_fd_sc_hd__mux2_1
XFILLER_9_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2467_ _2477_/CLK _2467_/D vssd1 vssd1 vccd1 vccd1 _2467_/Q sky130_fd_sc_hd__dfxtp_1
X_1418_ _2048_/Q _1984_/A1 _1419_/S vssd1 vssd1 vccd1 vccd1 _2048_/D sky130_fd_sc_hd__mux2_1
X_2398_ _2482_/CLK _2398_/D vssd1 vssd1 vccd1 vccd1 _2398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1349_ _1579_/A0 _2004_/Q _1350_/S vssd1 vssd1 vccd1 vccd1 _2004_/D sky130_fd_sc_hd__mux2_1
XFILLER_71_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2321_ _2363_/CLK _2321_/D vssd1 vssd1 vccd1 vccd1 _2321_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2252_ _2480_/CLK _2252_/D vssd1 vssd1 vccd1 vccd1 _2252_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1203_ _1234_/A1 _1201_/X _1020_/A vssd1 vssd1 vccd1 vccd1 _1203_/X sky130_fd_sc_hd__a21o_1
X_2183_ _2302_/CLK _2183_/D vssd1 vssd1 vccd1 vccd1 _2183_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1134_ _1453_/C _1133_/X _1385_/A vssd1 vssd1 vccd1 vccd1 _1134_/X sky130_fd_sc_hd__o21ba_1
XFILLER_53_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1065_ _1065_/A _1065_/B vssd1 vssd1 vccd1 vccd1 _1065_/X sky130_fd_sc_hd__and2_1
XFILLER_18_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1967_ _1972_/A0 _2482_/Q _1970_/S vssd1 vssd1 vccd1 vccd1 _2482_/D sky130_fd_sc_hd__mux2_1
X_1898_ _1903_/A0 _2427_/Q _1900_/S vssd1 vssd1 vccd1 vccd1 _2427_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1821_ _1821_/A _1901_/A vssd1 vssd1 vccd1 vccd1 _1825_/S sky130_fd_sc_hd__nand2_2
Xclkbuf_leaf_10_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _2094_/CLK sky130_fd_sc_hd__clkbuf_16
X_1752_ _2310_/Q _1762_/A0 _1755_/S vssd1 vssd1 vccd1 vccd1 _2310_/D sky130_fd_sc_hd__mux2_1
XFILLER_7_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1683_ _2255_/Q _1983_/A1 _1685_/S vssd1 vssd1 vccd1 vccd1 _2255_/D sky130_fd_sc_hd__mux2_1
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2304_ _2496_/CLK _2304_/D vssd1 vssd1 vccd1 vccd1 _2304_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2235_ _2240_/CLK _2235_/D vssd1 vssd1 vccd1 vccd1 _2235_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2166_ _2177_/CLK _2166_/D vssd1 vssd1 vccd1 vccd1 _2166_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1117_ _1409_/C _1115_/X _1116_/X _1295_/B2 vssd1 vssd1 vccd1 vccd1 _1118_/B sky130_fd_sc_hd__a22o_1
XFILLER_80_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2097_ _2097_/CLK _2097_/D vssd1 vssd1 vccd1 vccd1 _2097_/Q sky130_fd_sc_hd__dfxtp_1
X_1048_ _1048_/A _1048_/B _1048_/C _1048_/D vssd1 vssd1 vccd1 vccd1 _1048_/X sky130_fd_sc_hd__or4_1
XFILLER_0_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2020_ _2485_/CLK _2020_/D vssd1 vssd1 vccd1 vccd1 _2020_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1804_ _1804_/A0 _2352_/Q _1805_/S vssd1 vssd1 vccd1 vccd1 _2352_/D sky130_fd_sc_hd__mux2_1
X_1735_ _1960_/A0 _2297_/Q _1735_/S vssd1 vssd1 vccd1 vccd1 _2297_/D sky130_fd_sc_hd__mux2_1
X_1666_ _1666_/A _1906_/B vssd1 vssd1 vccd1 vccd1 _1670_/S sky130_fd_sc_hd__nor2_4
X_1597_ _2186_/Q _1662_/A0 _1600_/S vssd1 vssd1 vccd1 vccd1 _2186_/D sky130_fd_sc_hd__mux2_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2218_ _2229_/CLK _2218_/D vssd1 vssd1 vccd1 vccd1 _2218_/Q sky130_fd_sc_hd__dfxtp_1
X_2149_ _2159_/CLK _2149_/D vssd1 vssd1 vccd1 vccd1 _2149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1520_ _2125_/Q _1585_/A0 _1520_/S vssd1 vssd1 vccd1 vccd1 _2125_/D sky130_fd_sc_hd__mux2_1
X_1451_ _2072_/Q _1809_/A0 _1452_/S vssd1 vssd1 vccd1 vccd1 _2072_/D sky130_fd_sc_hd__mux2_1
X_1382_ _1904_/A0 _2024_/Q _1383_/S vssd1 vssd1 vccd1 vccd1 _2024_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2003_ _2177_/CLK _2003_/D vssd1 vssd1 vccd1 vccd1 _2003_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1718_ _2283_/Q _1738_/A0 _1720_/S vssd1 vssd1 vccd1 vccd1 _2283_/D sky130_fd_sc_hd__mux2_1
X_1649_ _1664_/A0 _2228_/Q _1650_/S vssd1 vssd1 vccd1 vccd1 _2228_/D sky130_fd_sc_hd__mux2_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1503_ _1503_/A0 _2111_/Q _1505_/S vssd1 vssd1 vccd1 vccd1 _2111_/D sky130_fd_sc_hd__mux2_1
X_2483_ _2485_/CLK _2483_/D vssd1 vssd1 vccd1 vccd1 _2483_/Q sky130_fd_sc_hd__dfxtp_1
X_1434_ _2059_/Q _1503_/A0 _1436_/S vssd1 vssd1 vccd1 vccd1 _2059_/D sky130_fd_sc_hd__mux2_1
X_1365_ _1935_/A0 _2013_/Q _1365_/S vssd1 vssd1 vccd1 vccd1 _2013_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1296_ _2165_/Q _2169_/Q _2173_/Q _2177_/Q _1297_/S0 _1297_/S1 vssd1 vssd1 vccd1
+ vccd1 _1296_/X sky130_fd_sc_hd__mux4_2
XFILLER_55_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1150_ _2339_/Q _1991_/Q _2347_/Q _2351_/Q _1245_/S0 _1409_/B vssd1 vssd1 vccd1 vccd1
+ _1150_/X sky130_fd_sc_hd__mux4_1
XFILLER_65_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1081_ _2050_/Q _2054_/Q _2058_/Q _2006_/Q _1303_/S0 _1304_/S1 vssd1 vssd1 vccd1
+ vccd1 _1081_/X sky130_fd_sc_hd__mux4_1
XFILLER_18_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1983_ _2495_/Q _1983_/A1 _1985_/S vssd1 vssd1 vccd1 vccd1 _2495_/D sky130_fd_sc_hd__mux2_1
X_2466_ _2479_/CLK _2466_/D vssd1 vssd1 vccd1 vccd1 _2466_/Q sky130_fd_sc_hd__dfxtp_1
X_1417_ _2047_/Q _1793_/A1 _1419_/S vssd1 vssd1 vccd1 vccd1 _2047_/D sky130_fd_sc_hd__mux2_1
X_2397_ _2485_/CLK _2397_/D vssd1 vssd1 vccd1 vccd1 _2397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1348_ _1583_/A0 _2003_/Q _1350_/S vssd1 vssd1 vccd1 vccd1 _2003_/D sky130_fd_sc_hd__mux2_1
XFILLER_56_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1279_ _1100_/A _1277_/X _1278_/X vssd1 vssd1 vccd1 vccd1 _1279_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_83_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout140 _1304_/S0 vssd1 vssd1 vccd1 vccd1 _1303_/S0 sky130_fd_sc_hd__buf_8
XFILLER_47_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2320_ _2320_/CLK _2320_/D vssd1 vssd1 vccd1 vccd1 _2320_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2251_ _2480_/CLK _2251_/D vssd1 vssd1 vccd1 vccd1 _2251_/Q sky130_fd_sc_hd__dfxtp_1
X_1202_ _2044_/Q _2048_/Q _1277_/S vssd1 vssd1 vccd1 vccd1 _1202_/X sky130_fd_sc_hd__mux2_1
X_2182_ _2302_/CLK _2182_/D vssd1 vssd1 vccd1 vccd1 _2182_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1133_ _2451_/Q _2455_/Q _2459_/Q _2027_/Q _1475_/A _1464_/B vssd1 vssd1 vccd1 vccd1
+ _1133_/X sky130_fd_sc_hd__mux4_1
XFILLER_65_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1064_ _2262_/Q _2302_/Q _1277_/S vssd1 vssd1 vccd1 vccd1 _1065_/B sky130_fd_sc_hd__mux2_1
XFILLER_80_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1966_ _1966_/A _1966_/B vssd1 vssd1 vccd1 vccd1 _1970_/S sky130_fd_sc_hd__or2_4
X_1897_ _1902_/A0 _2426_/Q _1900_/S vssd1 vssd1 vccd1 vccd1 _2426_/D sky130_fd_sc_hd__mux2_1
X_2449_ _2449_/CLK _2449_/D vssd1 vssd1 vccd1 vccd1 _2449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1820_ _1940_/A0 _2365_/Q _1820_/S vssd1 vssd1 vccd1 vccd1 _2365_/D sky130_fd_sc_hd__mux2_1
X_1751_ _1806_/A _1911_/A vssd1 vssd1 vccd1 vccd1 _1755_/S sky130_fd_sc_hd__nor2_4
XFILLER_7_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1682_ _2254_/Q _1982_/A1 _1685_/S vssd1 vssd1 vccd1 vccd1 _2254_/D sky130_fd_sc_hd__mux2_1
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2303_ _2385_/CLK _2303_/D vssd1 vssd1 vccd1 vccd1 _2303_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2234_ _2240_/CLK _2234_/D vssd1 vssd1 vccd1 vccd1 _2234_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2165_ _2176_/CLK _2165_/D vssd1 vssd1 vccd1 vccd1 _2165_/Q sky130_fd_sc_hd__dfxtp_1
X_1116_ _2051_/Q _2055_/Q _2059_/Q _2007_/Q _1303_/S0 _1304_/S1 vssd1 vssd1 vccd1
+ vccd1 _1116_/X sky130_fd_sc_hd__mux4_2
XFILLER_38_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2096_ _2097_/CLK _2096_/D vssd1 vssd1 vccd1 vccd1 _2096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1047_ _1043_/X _1046_/X _1354_/A vssd1 vssd1 vccd1 vccd1 _1048_/D sky130_fd_sc_hd__o21ba_1
XFILLER_80_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1949_ _2468_/Q _1964_/A0 _1950_/S vssd1 vssd1 vccd1 vccd1 _2468_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1803_ _1983_/A1 _2351_/Q _1805_/S vssd1 vssd1 vccd1 vccd1 _2351_/D sky130_fd_sc_hd__mux2_1
X_1734_ _1904_/A0 _2296_/Q _1735_/S vssd1 vssd1 vccd1 vccd1 _2296_/D sky130_fd_sc_hd__mux2_1
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1665_ _1965_/A0 _2241_/Q _1665_/S vssd1 vssd1 vccd1 vccd1 _2241_/D sky130_fd_sc_hd__mux2_1
X_1596_ _1646_/A _1916_/B vssd1 vssd1 vccd1 vccd1 _1600_/S sky130_fd_sc_hd__nor2_4
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2217_ _2229_/CLK _2217_/D vssd1 vssd1 vccd1 vccd1 _2217_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2148_ _2159_/CLK _2148_/D vssd1 vssd1 vccd1 vccd1 _2148_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2079_ _2335_/CLK _2079_/D vssd1 vssd1 vccd1 vccd1 _2079_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1450_ _2071_/Q _1778_/A0 _1452_/S vssd1 vssd1 vccd1 vccd1 _2071_/D sky130_fd_sc_hd__mux2_1
X_1381_ _1973_/A0 _2023_/Q _1383_/S vssd1 vssd1 vccd1 vccd1 _2023_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2002_ _2232_/CLK _2002_/D vssd1 vssd1 vccd1 vccd1 _2002_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1717_ _2282_/Q _1732_/A0 _1720_/S vssd1 vssd1 vccd1 vccd1 _2282_/D sky130_fd_sc_hd__mux2_1
X_1648_ _1663_/A0 _2227_/Q _1650_/S vssd1 vssd1 vccd1 vccd1 _2227_/D sky130_fd_sc_hd__mux2_1
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1579_ _1579_/A0 _2172_/Q _1580_/S vssd1 vssd1 vccd1 vccd1 _2172_/D sky130_fd_sc_hd__mux2_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2482_ _2482_/CLK _2482_/D vssd1 vssd1 vccd1 vccd1 _2482_/Q sky130_fd_sc_hd__dfxtp_1
X_1502_ _1777_/A0 _2110_/Q _1505_/S vssd1 vssd1 vccd1 vccd1 _2110_/D sky130_fd_sc_hd__mux2_1
X_1433_ _2058_/Q _1762_/A0 _1436_/S vssd1 vssd1 vccd1 vccd1 _2058_/D sky130_fd_sc_hd__mux2_1
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1364_ _1739_/A0 _2012_/Q _1365_/S vssd1 vssd1 vccd1 vccd1 _2012_/D sky130_fd_sc_hd__mux2_1
X_1295_ _1020_/X _1291_/X _1293_/X _1294_/X _1295_/B2 vssd1 vssd1 vccd1 vccd1 _1295_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_63_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1080_ _2098_/Q _2014_/Q _2106_/Q _2110_/Q _1303_/S0 _1304_/S1 vssd1 vssd1 vccd1
+ vccd1 _1080_/X sky130_fd_sc_hd__mux4_1
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1982_ _2494_/Q _1982_/A1 _1985_/S vssd1 vssd1 vccd1 vccd1 _2494_/D sky130_fd_sc_hd__mux2_1
XFILLER_13_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2465_ _2497_/CLK _2465_/D vssd1 vssd1 vccd1 vccd1 _2465_/Q sky130_fd_sc_hd__dfxtp_1
X_2396_ _2482_/CLK _2396_/D vssd1 vssd1 vccd1 vccd1 _2396_/Q sky130_fd_sc_hd__dfxtp_1
X_1416_ _2046_/Q _1792_/A1 _1419_/S vssd1 vssd1 vccd1 vccd1 _2046_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1347_ _1582_/A0 _2002_/Q _1350_/S vssd1 vssd1 vccd1 vccd1 _2002_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1278_ _0992_/Y _1276_/X _1020_/A vssd1 vssd1 vccd1 vccd1 _1278_/X sky130_fd_sc_hd__a21o_1
XFILLER_36_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout130 _1420_/A vssd1 vssd1 vccd1 vccd1 _1464_/A sky130_fd_sc_hd__buf_12
Xfanout141 fanout148/X vssd1 vssd1 vccd1 vccd1 _1304_/S0 sky130_fd_sc_hd__buf_6
XFILLER_59_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2250_ _2457_/CLK _2250_/D vssd1 vssd1 vccd1 vccd1 _2250_/Q sky130_fd_sc_hd__dfxtp_1
X_1201_ _2036_/Q _2040_/Q _1277_/S vssd1 vssd1 vccd1 vccd1 _1201_/X sky130_fd_sc_hd__mux2_1
X_2181_ _2368_/CLK _2181_/D vssd1 vssd1 vccd1 vccd1 _2181_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1132_ _1244_/A1 _1123_/Y _1125_/Y _1130_/Y _1131_/Y vssd1 vssd1 vccd1 vccd1 _1132_/X
+ sky130_fd_sc_hd__o32a_1
X_1063_ _1040_/B _1053_/X _1055_/X _1062_/X input6/X vssd1 vssd1 vccd1 vccd1 _1063_/X
+ sky130_fd_sc_hd__o311a_2
XFILLER_18_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1965_ _1965_/A0 _2481_/Q _1965_/S vssd1 vssd1 vccd1 vccd1 _2481_/D sky130_fd_sc_hd__mux2_1
X_1896_ _1901_/B _1976_/B vssd1 vssd1 vccd1 vccd1 _1900_/S sky130_fd_sc_hd__nand2_2
X_2448_ _2448_/CLK _2448_/D vssd1 vssd1 vccd1 vccd1 _2448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2379_ _2485_/CLK _2379_/D vssd1 vssd1 vccd1 vccd1 _2379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1750_ _2309_/Q _1765_/A0 _1750_/S vssd1 vssd1 vccd1 vccd1 _2309_/D sky130_fd_sc_hd__mux2_1
XFILLER_7_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1681_ _1726_/A _1681_/B vssd1 vssd1 vccd1 vccd1 _1685_/S sky130_fd_sc_hd__nor2_4
X_2302_ _2302_/CLK _2302_/D vssd1 vssd1 vccd1 vccd1 _2302_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2233_ _2241_/CLK _2233_/D vssd1 vssd1 vccd1 vccd1 _2233_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2164_ _2176_/CLK _2164_/D vssd1 vssd1 vccd1 vccd1 _2164_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1115_ _2099_/Q _2015_/Q _2107_/Q _2111_/Q _1303_/S0 _1304_/S1 vssd1 vssd1 vccd1
+ vccd1 _1115_/X sky130_fd_sc_hd__mux4_1
X_2095_ _2097_/CLK _2095_/D vssd1 vssd1 vccd1 vccd1 _2095_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1046_ _1409_/C _1044_/X _1045_/X _1295_/B2 vssd1 vssd1 vccd1 vccd1 _1046_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1948_ _2467_/Q _1963_/A0 _1950_/S vssd1 vssd1 vccd1 vccd1 _2467_/D sky130_fd_sc_hd__mux2_1
X_1879_ _1884_/A0 _2412_/Q _1880_/S vssd1 vssd1 vccd1 vccd1 _2412_/D sky130_fd_sc_hd__mux2_1
XFILLER_76_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_451 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_3__f_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_3__f_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_75_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1802_ _1822_/A0 _2350_/Q _1805_/S vssd1 vssd1 vccd1 vccd1 _2350_/D sky130_fd_sc_hd__mux2_1
X_1733_ _1738_/A0 _2295_/Q _1735_/S vssd1 vssd1 vccd1 vccd1 _2295_/D sky130_fd_sc_hd__mux2_1
X_1664_ _1664_/A0 _2240_/Q _1665_/S vssd1 vssd1 vccd1 vccd1 _2240_/D sky130_fd_sc_hd__mux2_1
X_1595_ _2185_/Q _1845_/A1 _1595_/S vssd1 vssd1 vccd1 vccd1 _2185_/D sky130_fd_sc_hd__mux2_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2216_ _2229_/CLK _2216_/D vssd1 vssd1 vccd1 vccd1 _2216_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2147_ _2493_/CLK _2147_/D vssd1 vssd1 vccd1 vccd1 _2147_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2078_ _2335_/CLK _2078_/D vssd1 vssd1 vccd1 vccd1 _2078_/Q sky130_fd_sc_hd__dfxtp_1
X_1029_ _1464_/B _1029_/B vssd1 vssd1 vccd1 vccd1 _1029_/X sky130_fd_sc_hd__or2_1
XFILLER_30_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1380_ _1902_/A0 _2022_/Q _1383_/S vssd1 vssd1 vccd1 vccd1 _2022_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2001_ _2320_/CLK _2001_/D vssd1 vssd1 vccd1 vccd1 _2001_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1716_ _1726_/A _1956_/B vssd1 vssd1 vccd1 vccd1 _1720_/S sky130_fd_sc_hd__nor2_2
X_1647_ _1662_/A0 _2226_/Q _1650_/S vssd1 vssd1 vccd1 vccd1 _2226_/D sky130_fd_sc_hd__mux2_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1578_ _1583_/A0 _2171_/Q _1580_/S vssd1 vssd1 vccd1 vccd1 _2171_/D sky130_fd_sc_hd__mux2_1
XFILLER_58_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2481_ _2481_/CLK _2481_/D vssd1 vssd1 vccd1 vccd1 _2481_/Q sky130_fd_sc_hd__dfxtp_1
X_1501_ _1501_/A _1901_/A vssd1 vssd1 vccd1 vccd1 _1505_/S sky130_fd_sc_hd__nand2_4
X_1432_ _1486_/A _1916_/B vssd1 vssd1 vccd1 vccd1 _1436_/S sky130_fd_sc_hd__nor2_4
XFILLER_68_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1363_ _1963_/A0 _2011_/Q _1365_/S vssd1 vssd1 vccd1 vccd1 _2011_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1294_ _2117_/Q _2121_/Q _2125_/Q _2129_/Q _1297_/S0 _1291_/A vssd1 vssd1 vccd1 vccd1
+ _1294_/X sky130_fd_sc_hd__mux4_1
XFILLER_55_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1981_ _1981_/A _1981_/B vssd1 vssd1 vccd1 vccd1 _1985_/S sky130_fd_sc_hd__nor2_2
Xclkbuf_leaf_40_clk clkbuf_leaf_4_clk/A vssd1 vssd1 vccd1 vccd1 _2448_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2464_ _2497_/CLK _2464_/D vssd1 vssd1 vccd1 vccd1 _2464_/Q sky130_fd_sc_hd__dfxtp_1
X_2395_ _2485_/CLK _2395_/D vssd1 vssd1 vccd1 vccd1 _2395_/Q sky130_fd_sc_hd__dfxtp_1
X_1415_ _1901_/A _1941_/B vssd1 vssd1 vccd1 vccd1 _1419_/S sky130_fd_sc_hd__and2_2
X_1346_ _1861_/A _1581_/A vssd1 vssd1 vccd1 vccd1 _1350_/S sky130_fd_sc_hd__nand2_2
XFILLER_68_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1277_ _2045_/Q _2049_/Q _1277_/S vssd1 vssd1 vccd1 vccd1 _1277_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_31_clk clkbuf_2_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _2416_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_3_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout131 _1420_/A vssd1 vssd1 vccd1 vccd1 _1287_/S0 sky130_fd_sc_hd__buf_8
Xfanout120 _1884_/A0 vssd1 vssd1 vccd1 vccd1 _1964_/A0 sky130_fd_sc_hd__clkbuf_2
XFILLER_47_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout142 _1233_/S vssd1 vssd1 vccd1 vccd1 _1240_/S sky130_fd_sc_hd__buf_6
XFILLER_47_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_22_clk clkbuf_2_3__f_clk/X vssd1 vssd1 vccd1 vccd1 _2302_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_42_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2180_ _2320_/CLK _2180_/D vssd1 vssd1 vccd1 vccd1 _2180_/Q sky130_fd_sc_hd__dfxtp_1
X_1200_ _2344_/Q _2496_/Q _2424_/Q _2464_/Q _1275_/S0 _1100_/A vssd1 vssd1 vccd1 vccd1
+ _1200_/X sky130_fd_sc_hd__mux4_1
X_1131_ _1220_/A _1126_/X _1024_/B vssd1 vssd1 vccd1 vccd1 _1131_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_65_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1062_ _1058_/X _1061_/X _1040_/B vssd1 vssd1 vccd1 vccd1 _1062_/X sky130_fd_sc_hd__a21bo_1
XFILLER_33_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1964_ _1964_/A0 _2480_/Q _1965_/S vssd1 vssd1 vccd1 vccd1 _2480_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_13_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _2337_/CLK sky130_fd_sc_hd__clkbuf_16
X_1895_ _2425_/Q _1985_/A1 _1895_/S vssd1 vssd1 vccd1 vccd1 _2425_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2447_ _2448_/CLK _2447_/D vssd1 vssd1 vccd1 vccd1 _2447_/Q sky130_fd_sc_hd__dfxtp_1
X_2378_ _2482_/CLK _2378_/D vssd1 vssd1 vccd1 vccd1 _2378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1329_ input7/X _1329_/B vssd1 vssd1 vccd1 vccd1 _1398_/B sky130_fd_sc_hd__nand2b_4
XFILLER_12_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1680_ _2253_/Q _1935_/A0 _1680_/S vssd1 vssd1 vccd1 vccd1 _2253_/D sky130_fd_sc_hd__mux2_1
XFILLER_7_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2301_ _2301_/CLK _2301_/D vssd1 vssd1 vccd1 vccd1 _2301_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2232_ _2232_/CLK _2232_/D vssd1 vssd1 vccd1 vccd1 _2232_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_2_clk clkbuf_leaf_4_clk/A vssd1 vssd1 vccd1 vccd1 _2241_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2163_ _2176_/CLK _2163_/D vssd1 vssd1 vccd1 vccd1 _2163_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1114_ _1298_/B2 _1112_/X _1113_/X _1020_/X vssd1 vssd1 vccd1 vccd1 _1118_/A sky130_fd_sc_hd__a22o_1
X_2094_ _2094_/CLK _2094_/D vssd1 vssd1 vccd1 vccd1 _2094_/Q sky130_fd_sc_hd__dfxtp_1
X_1045_ _2306_/Q _2310_/Q _2314_/Q _2318_/Q _1285_/S0 _1285_/S1 vssd1 vssd1 vccd1
+ vccd1 _1045_/X sky130_fd_sc_hd__mux4_2
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1947_ _2466_/Q _1962_/A0 _1950_/S vssd1 vssd1 vccd1 vccd1 _2466_/D sky130_fd_sc_hd__mux2_1
X_1878_ _1903_/A0 _2411_/Q _1880_/S vssd1 vssd1 vccd1 vccd1 _2411_/D sky130_fd_sc_hd__mux2_1
XFILLER_76_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1801_ _1821_/A _1961_/A vssd1 vssd1 vccd1 vccd1 _1805_/S sky130_fd_sc_hd__nand2_2
X_1732_ _1732_/A0 _2294_/Q _1735_/S vssd1 vssd1 vccd1 vccd1 _2294_/D sky130_fd_sc_hd__mux2_1
XFILLER_7_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1663_ _1663_/A0 _2239_/Q _1665_/S vssd1 vssd1 vccd1 vccd1 _2239_/D sky130_fd_sc_hd__mux2_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1594_ _2184_/Q _1739_/A0 _1595_/S vssd1 vssd1 vccd1 vccd1 _2184_/D sky130_fd_sc_hd__mux2_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2215_ _2479_/CLK _2215_/D vssd1 vssd1 vccd1 vccd1 _2215_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2146_ _2493_/CLK _2146_/D vssd1 vssd1 vccd1 vccd1 _2146_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2077_ _2097_/CLK _2077_/D vssd1 vssd1 vccd1 vccd1 _2077_/Q sky130_fd_sc_hd__dfxtp_1
X_1028_ _2402_/Q _2406_/Q _1181_/S vssd1 vssd1 vccd1 vccd1 _1029_/B sky130_fd_sc_hd__mux2_1
XFILLER_30_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2000_ _2320_/CLK _2000_/D vssd1 vssd1 vccd1 vccd1 _2000_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1715_ _2281_/Q _1960_/A0 _1715_/S vssd1 vssd1 vccd1 vccd1 _2281_/D sky130_fd_sc_hd__mux2_1
X_1646_ _1646_/A _1966_/B vssd1 vssd1 vccd1 vccd1 _1650_/S sky130_fd_sc_hd__or2_4
X_1577_ _1582_/A0 _2170_/Q _1580_/S vssd1 vssd1 vccd1 vccd1 _2170_/D sky130_fd_sc_hd__mux2_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2129_ _2232_/CLK _2129_/D vssd1 vssd1 vccd1 vccd1 _2129_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2480_ _2480_/CLK _2480_/D vssd1 vssd1 vccd1 vccd1 _2480_/Q sky130_fd_sc_hd__dfxtp_1
X_1500_ _1505_/A0 _2109_/Q _1500_/S vssd1 vssd1 vccd1 vccd1 _2109_/D sky130_fd_sc_hd__mux2_1
X_1431_ _1475_/A _1475_/B _1431_/C vssd1 vssd1 vccd1 vccd1 _1916_/B sky130_fd_sc_hd__or3_4
X_1362_ _1732_/A0 _2010_/Q _1365_/S vssd1 vssd1 vccd1 vccd1 _2010_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1293_ _1475_/B _1293_/B vssd1 vssd1 vccd1 vccd1 _1293_/X sky130_fd_sc_hd__or2_1
XFILLER_83_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1629_ _2212_/Q _1979_/A0 _1630_/S vssd1 vssd1 vccd1 vccd1 _2212_/D sky130_fd_sc_hd__mux2_1
XFILLER_59_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1980_ _1980_/A0 _2493_/Q _1980_/S vssd1 vssd1 vccd1 vccd1 _2493_/D sky130_fd_sc_hd__mux2_1
XFILLER_33_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2463_ _2495_/CLK _2463_/D vssd1 vssd1 vccd1 vccd1 _2463_/Q sky130_fd_sc_hd__dfxtp_1
X_2394_ _2477_/CLK _2394_/D vssd1 vssd1 vccd1 vccd1 _2394_/Q sky130_fd_sc_hd__dfxtp_1
X_1414_ _1845_/A1 _2045_/Q _1414_/S vssd1 vssd1 vccd1 vccd1 _2045_/D sky130_fd_sc_hd__mux2_1
X_1345_ _1373_/A _1398_/B vssd1 vssd1 vccd1 vccd1 _1531_/B sky130_fd_sc_hd__or2_4
XFILLER_28_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1276_ _2037_/Q _2041_/Q _1277_/S vssd1 vssd1 vccd1 vccd1 _1276_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout121 _1884_/A0 vssd1 vssd1 vccd1 vccd1 _1904_/A0 sky130_fd_sc_hd__buf_4
XFILLER_59_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout110 input11/X vssd1 vssd1 vccd1 vccd1 _1965_/A0 sky130_fd_sc_hd__buf_4
Xfanout132 _1182_/S vssd1 vssd1 vccd1 vccd1 _1420_/A sky130_fd_sc_hd__buf_6
Xfanout143 _1233_/S vssd1 vssd1 vccd1 vccd1 _1245_/S0 sky130_fd_sc_hd__buf_6
XFILLER_59_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1130_ _0992_/A _1128_/X _1129_/X vssd1 vssd1 vccd1 vccd1 _1130_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_80_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1061_ _1396_/C _1059_/X _1060_/X _1420_/C vssd1 vssd1 vccd1 vccd1 _1061_/X sky130_fd_sc_hd__o22a_1
XFILLER_73_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1963_ _1963_/A0 _2479_/Q _1965_/S vssd1 vssd1 vccd1 vccd1 _2479_/D sky130_fd_sc_hd__mux2_1
X_1894_ _2424_/Q _1944_/A0 _1895_/S vssd1 vssd1 vccd1 vccd1 _2424_/D sky130_fd_sc_hd__mux2_1
X_2446_ _2449_/CLK _2446_/D vssd1 vssd1 vccd1 vccd1 _2446_/Q sky130_fd_sc_hd__dfxtp_1
X_2377_ _2485_/CLK _2377_/D vssd1 vssd1 vccd1 vccd1 _2377_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1328_ _1360_/A _1475_/C vssd1 vssd1 vccd1 vccd1 _1961_/A sky130_fd_sc_hd__nor2_8
XFILLER_83_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1259_ _1257_/X _1258_/X _1254_/X vssd1 vssd1 vccd1 vccd1 _1259_/X sky130_fd_sc_hd__a21o_1
XFILLER_56_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2300_ _2480_/CLK _2300_/D vssd1 vssd1 vccd1 vccd1 _2300_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2231_ _2240_/CLK _2231_/D vssd1 vssd1 vccd1 vccd1 _2231_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2162_ _2177_/CLK _2162_/D vssd1 vssd1 vccd1 vccd1 _2162_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1113_ _2083_/Q _2087_/Q _2091_/Q _2095_/Q _1304_/S0 _1301_/S1 vssd1 vssd1 vccd1
+ vccd1 _1113_/X sky130_fd_sc_hd__mux4_1
X_2093_ _2097_/CLK _2093_/D vssd1 vssd1 vccd1 vccd1 _2093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1044_ _2354_/Q _2358_/Q _2362_/Q _2366_/Q _1285_/S0 _1285_/S1 vssd1 vssd1 vccd1
+ vccd1 _1044_/X sky130_fd_sc_hd__mux4_1
XFILLER_65_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1946_ _1966_/A _1946_/B vssd1 vssd1 vccd1 vccd1 _1950_/S sky130_fd_sc_hd__nor2_2
X_1877_ _1902_/A0 _2410_/Q _1880_/S vssd1 vssd1 vccd1 vccd1 _2410_/D sky130_fd_sc_hd__mux2_1
X_2429_ _2433_/CLK _2429_/D vssd1 vssd1 vccd1 vccd1 _2429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1800_ _1800_/A0 _2349_/Q _1800_/S vssd1 vssd1 vccd1 vccd1 _2349_/D sky130_fd_sc_hd__mux2_1
X_1731_ _1736_/A _1971_/A vssd1 vssd1 vccd1 vccd1 _1735_/S sky130_fd_sc_hd__nand2_2
X_1662_ _1662_/A0 _2238_/Q _1665_/S vssd1 vssd1 vccd1 vccd1 _2238_/D sky130_fd_sc_hd__mux2_1
X_1593_ _2183_/Q _1783_/A0 _1595_/S vssd1 vssd1 vccd1 vccd1 _2183_/D sky130_fd_sc_hd__mux2_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2214_ _2479_/CLK _2214_/D vssd1 vssd1 vccd1 vccd1 _2214_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2145_ _2385_/CLK _2145_/D vssd1 vssd1 vccd1 vccd1 _2145_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2076_ _2349_/CLK _2076_/D vssd1 vssd1 vccd1 vccd1 _2076_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1027_ _1420_/C _1019_/X _1026_/X _1016_/X vssd1 vssd1 vccd1 vccd1 _1048_/B sky130_fd_sc_hd__o211a_1
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1929_ _2452_/Q _1964_/A0 _1930_/S vssd1 vssd1 vccd1 vccd1 _2452_/D sky130_fd_sc_hd__mux2_1
XFILLER_30_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1714_ _2280_/Q _1904_/A0 _1715_/S vssd1 vssd1 vccd1 vccd1 _2280_/D sky130_fd_sc_hd__mux2_1
X_1645_ _2225_/Q _1845_/A1 _1645_/S vssd1 vssd1 vccd1 vccd1 _2225_/D sky130_fd_sc_hd__mux2_1
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1576_ _1581_/A _1976_/B vssd1 vssd1 vccd1 vccd1 _1580_/S sky130_fd_sc_hd__nand2_4
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2128_ _2232_/CLK _2128_/D vssd1 vssd1 vccd1 vccd1 _2128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2059_ _2113_/CLK _2059_/D vssd1 vssd1 vccd1 vccd1 _2059_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1430_ _2057_/Q _1505_/A0 _1430_/S vssd1 vssd1 vccd1 vccd1 _2057_/D sky130_fd_sc_hd__mux2_1
X_1361_ _1736_/A _1901_/A vssd1 vssd1 vccd1 vccd1 _1365_/S sky130_fd_sc_hd__nand2_2
X_1292_ _2157_/Q _2161_/Q _1292_/S vssd1 vssd1 vccd1 vccd1 _1293_/B sky130_fd_sc_hd__mux2_1
XFILLER_55_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1628_ _2211_/Q _1663_/A0 _1630_/S vssd1 vssd1 vccd1 vccd1 _2211_/D sky130_fd_sc_hd__mux2_1
X_1559_ _2156_/Q _1974_/A0 _1560_/S vssd1 vssd1 vccd1 vccd1 _2156_/D sky130_fd_sc_hd__mux2_1
XTAP_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_47 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2462_ _2497_/CLK _2462_/D vssd1 vssd1 vccd1 vccd1 _2462_/Q sky130_fd_sc_hd__dfxtp_1
X_2393_ _2433_/CLK _2393_/D vssd1 vssd1 vccd1 vccd1 _2393_/Q sky130_fd_sc_hd__dfxtp_1
X_1413_ _1984_/A1 _2044_/Q _1414_/S vssd1 vssd1 vccd1 vccd1 _2044_/D sky130_fd_sc_hd__mux2_1
XFILLER_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1344_ _1373_/A _1398_/B vssd1 vssd1 vccd1 vccd1 _1581_/A sky130_fd_sc_hd__nor2_8
X_1275_ _2345_/Q _2497_/Q _2425_/Q _2465_/Q _1275_/S0 _1065_/A vssd1 vssd1 vccd1 vccd1
+ _1275_/X sky130_fd_sc_hd__mux4_1
XFILLER_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout100 _1965_/A0 vssd1 vssd1 vccd1 vccd1 _1960_/A0 sky130_fd_sc_hd__buf_4
Xfanout111 _1664_/A0 vssd1 vssd1 vccd1 vccd1 _1579_/A0 sky130_fd_sc_hd__clkbuf_4
Xfanout122 fanout127/X vssd1 vssd1 vccd1 vccd1 _1884_/A0 sky130_fd_sc_hd__clkbuf_4
Xfanout133 _1182_/S vssd1 vssd1 vccd1 vccd1 _1253_/S0 sky130_fd_sc_hd__buf_8
XFILLER_59_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout144 _1233_/S vssd1 vssd1 vccd1 vccd1 _1277_/S sky130_fd_sc_hd__buf_6
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1060_ _2178_/Q _1998_/Q _2186_/Q _2190_/Q _1287_/S0 _1013_/B vssd1 vssd1 vccd1 vccd1
+ _1060_/X sky130_fd_sc_hd__mux4_2
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1962_ _1962_/A0 _2478_/Q _1965_/S vssd1 vssd1 vccd1 vccd1 _2478_/D sky130_fd_sc_hd__mux2_1
X_1893_ _2423_/Q _1983_/A1 _1895_/S vssd1 vssd1 vccd1 vccd1 _2423_/D sky130_fd_sc_hd__mux2_1
X_2445_ _2449_/CLK _2445_/D vssd1 vssd1 vccd1 vccd1 _2445_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2376_ _2485_/CLK _2376_/D vssd1 vssd1 vccd1 vccd1 _2376_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1327_ _1800_/A0 _1993_/Q _1327_/S vssd1 vssd1 vccd1 vccd1 _1993_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1258_ _1258_/A _1258_/B vssd1 vssd1 vccd1 vccd1 _1258_/X sky130_fd_sc_hd__or2_1
XFILLER_83_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1189_ _2356_/Q _2360_/Q _2364_/Q _2368_/Q _1285_/S0 _1285_/S1 vssd1 vssd1 vccd1
+ vccd1 _1189_/X sky130_fd_sc_hd__mux4_1
XFILLER_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2230_ _2240_/CLK _2230_/D vssd1 vssd1 vccd1 vccd1 _2230_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2161_ _2448_/CLK _2161_/D vssd1 vssd1 vccd1 vccd1 _2161_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1112_ _2067_/Q _2071_/Q _2075_/Q _2079_/Q _1304_/S0 _1301_/S1 vssd1 vssd1 vccd1
+ vccd1 _1112_/X sky130_fd_sc_hd__mux4_2
X_2092_ _2367_/CLK _2092_/D vssd1 vssd1 vccd1 vccd1 _2092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1043_ _1298_/B2 _1041_/X _1042_/X _1020_/X vssd1 vssd1 vccd1 vccd1 _1043_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1945_ _1985_/A1 _2465_/Q _1945_/S vssd1 vssd1 vccd1 vccd1 _2465_/D sky130_fd_sc_hd__mux2_1
XFILLER_9_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1876_ _1886_/A _1956_/B vssd1 vssd1 vccd1 vccd1 _1880_/S sky130_fd_sc_hd__or2_4
X_2428_ _2432_/CLK _2428_/D vssd1 vssd1 vccd1 vccd1 _2428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2359_ _2367_/CLK _2359_/D vssd1 vssd1 vccd1 vccd1 _2359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1730_ _2293_/Q _1740_/A0 _1730_/S vssd1 vssd1 vccd1 vccd1 _2293_/D sky130_fd_sc_hd__mux2_1
XFILLER_7_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1661_ _1661_/A _1901_/A vssd1 vssd1 vccd1 vccd1 _1665_/S sky130_fd_sc_hd__nand2_4
X_1592_ _2182_/Q _1742_/A0 _1595_/S vssd1 vssd1 vccd1 vccd1 _2182_/D sky130_fd_sc_hd__mux2_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2213_ _2229_/CLK _2213_/D vssd1 vssd1 vccd1 vccd1 _2213_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_443 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2144_ _2496_/CLK _2144_/D vssd1 vssd1 vccd1 vccd1 _2144_/Q sky130_fd_sc_hd__dfxtp_1
X_2075_ _2335_/CLK _2075_/D vssd1 vssd1 vccd1 vccd1 _2075_/Q sky130_fd_sc_hd__dfxtp_1
X_1026_ _1464_/C _1022_/X _1396_/C _1025_/X vssd1 vssd1 vccd1 vccd1 _1026_/X sky130_fd_sc_hd__o22a_1
XFILLER_22_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1928_ _2451_/Q _1963_/A0 _1930_/S vssd1 vssd1 vccd1 vccd1 _2451_/D sky130_fd_sc_hd__mux2_1
X_1859_ _1969_/A0 _2396_/Q _1860_/S vssd1 vssd1 vccd1 vccd1 _2396_/D sky130_fd_sc_hd__mux2_1
XFILLER_1_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1713_ _2279_/Q _1963_/A0 _1715_/S vssd1 vssd1 vccd1 vccd1 _2279_/D sky130_fd_sc_hd__mux2_1
XFILLER_6_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1644_ _2224_/Q _1739_/A0 _1645_/S vssd1 vssd1 vccd1 vccd1 _2224_/D sky130_fd_sc_hd__mux2_1
X_1575_ _1585_/A0 _2169_/Q _1575_/S vssd1 vssd1 vccd1 vccd1 _2169_/D sky130_fd_sc_hd__mux2_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2127_ _2176_/CLK _2127_/D vssd1 vssd1 vccd1 vccd1 _2127_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2058_ _2094_/CLK _2058_/D vssd1 vssd1 vccd1 vccd1 _2058_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1009_ _1398_/A _1009_/B vssd1 vssd1 vccd1 vccd1 _1009_/Y sky130_fd_sc_hd__nor2_1
XFILLER_22_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1360_ _1360_/A _1360_/B vssd1 vssd1 vccd1 vccd1 _1901_/A sky130_fd_sc_hd__nor2_8
X_1291_ _1291_/A _1291_/B vssd1 vssd1 vccd1 vccd1 _1291_/X sky130_fd_sc_hd__or2_1
XFILLER_63_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_43_clk clkbuf_leaf_4_clk/A vssd1 vssd1 vccd1 vccd1 _2176_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1627_ _2210_/Q _1917_/A1 _1630_/S vssd1 vssd1 vccd1 vccd1 _2210_/D sky130_fd_sc_hd__mux2_1
X_1558_ _2155_/Q _1918_/A1 _1560_/S vssd1 vssd1 vccd1 vccd1 _2155_/D sky130_fd_sc_hd__mux2_1
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1489_ _2100_/Q _1784_/A0 _1490_/S vssd1 vssd1 vccd1 vccd1 _2100_/D sky130_fd_sc_hd__mux2_1
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_34_clk clkbuf_2_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _2433_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_22_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_25_clk clkbuf_2_3__f_clk/X vssd1 vssd1 vccd1 vccd1 _2297_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_41_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2461_ _2461_/CLK _2461_/D vssd1 vssd1 vccd1 vccd1 _2461_/Q sky130_fd_sc_hd__dfxtp_1
X_1412_ _1793_/A1 _2043_/Q _1414_/S vssd1 vssd1 vccd1 vccd1 _2043_/D sky130_fd_sc_hd__mux2_1
X_2392_ _2433_/CLK _2392_/D vssd1 vssd1 vccd1 vccd1 _2392_/Q sky130_fd_sc_hd__dfxtp_1
X_1343_ _1453_/C _1360_/A vssd1 vssd1 vccd1 vccd1 _1861_/A sky130_fd_sc_hd__nor2_8
X_1274_ _1274_/A _1274_/B vssd1 vssd1 vccd1 vccd1 _1274_/Y sky130_fd_sc_hd__nor2_1
XFILLER_76_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_16_clk clkbuf_2_3__f_clk/X vssd1 vssd1 vccd1 vccd1 _2457_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_51_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout112 fanout127/X vssd1 vssd1 vccd1 vccd1 _1664_/A0 sky130_fd_sc_hd__clkbuf_4
Xfanout101 fanout109/X vssd1 vssd1 vccd1 vccd1 _1765_/A0 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout145 _1275_/S0 vssd1 vssd1 vccd1 vccd1 _1270_/S sky130_fd_sc_hd__clkbuf_4
Xfanout134 _1182_/S vssd1 vssd1 vccd1 vccd1 _1256_/S0 sky130_fd_sc_hd__buf_4
Xfanout123 _1944_/A0 vssd1 vssd1 vccd1 vccd1 _1804_/A0 sky130_fd_sc_hd__buf_4
XFILLER_74_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1961_ _1961_/A _1976_/A vssd1 vssd1 vccd1 vccd1 _1965_/S sky130_fd_sc_hd__nand2_2
X_1892_ _2422_/Q _1982_/A1 _1895_/S vssd1 vssd1 vccd1 vccd1 _2422_/D sky130_fd_sc_hd__mux2_1
X_2444_ _2448_/CLK _2444_/D vssd1 vssd1 vccd1 vccd1 _2444_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_5_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _2368_/CLK sky130_fd_sc_hd__clkbuf_16
X_2375_ _2485_/CLK _2375_/D vssd1 vssd1 vccd1 vccd1 _2375_/Q sky130_fd_sc_hd__dfxtp_1
X_1326_ _1804_/A0 _1992_/Q _1327_/S vssd1 vssd1 vccd1 vccd1 _1992_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1257_ _1180_/A _1256_/X input4/X vssd1 vssd1 vccd1 vccd1 _1257_/X sky130_fd_sc_hd__o21a_1
X_1188_ _1302_/A1 _1186_/X _1187_/X _1020_/X vssd1 vssd1 vccd1 vccd1 _1188_/X sky130_fd_sc_hd__a22o_1
XFILLER_71_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2160_ _2176_/CLK _2160_/D vssd1 vssd1 vccd1 vccd1 _2160_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2091_ _2097_/CLK _2091_/D vssd1 vssd1 vccd1 vccd1 _2091_/Q sky130_fd_sc_hd__dfxtp_1
X_1111_ _1244_/A1 _1104_/X _1109_/Y _1110_/Y vssd1 vssd1 vccd1 vccd1 _1111_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1042_ _2338_/Q _1990_/Q _2346_/Q _2350_/Q _1285_/S0 _1409_/B vssd1 vssd1 vccd1 vccd1
+ _1042_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1944_ _1944_/A0 _2464_/Q _1945_/S vssd1 vssd1 vccd1 vccd1 _2464_/D sky130_fd_sc_hd__mux2_1
X_1875_ _1905_/A0 _2409_/Q _1875_/S vssd1 vssd1 vccd1 vccd1 _2409_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2427_ _2433_/CLK _2427_/D vssd1 vssd1 vccd1 vccd1 _2427_/Q sky130_fd_sc_hd__dfxtp_1
X_2358_ _2368_/CLK _2358_/D vssd1 vssd1 vccd1 vccd1 _2358_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2289_ _2416_/CLK _2289_/D vssd1 vssd1 vccd1 vccd1 _2289_/Q sky130_fd_sc_hd__dfxtp_1
X_1309_ _1310_/A _1366_/A vssd1 vssd1 vccd1 vccd1 _1931_/A sky130_fd_sc_hd__nor2_8
XFILLER_84_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1660_ _1660_/A0 _2237_/Q _1660_/S vssd1 vssd1 vccd1 vccd1 _2237_/D sky130_fd_sc_hd__mux2_1
X_1591_ _1981_/B _1926_/B vssd1 vssd1 vccd1 vccd1 _1595_/S sky130_fd_sc_hd__nor2_2
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2212_ _2229_/CLK _2212_/D vssd1 vssd1 vccd1 vccd1 _2212_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2143_ _2385_/CLK _2143_/D vssd1 vssd1 vccd1 vccd1 _2143_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2074_ _2335_/CLK _2074_/D vssd1 vssd1 vccd1 vccd1 _2074_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1025_ _2482_/Q _2486_/Q _2490_/Q _2030_/Q _1292_/S _1253_/S1 vssd1 vssd1 vccd1 vccd1
+ _1025_/X sky130_fd_sc_hd__mux4_2
XFILLER_22_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1927_ _2450_/Q _1962_/A0 _1930_/S vssd1 vssd1 vccd1 vccd1 _2450_/D sky130_fd_sc_hd__mux2_1
X_1858_ _1973_/A0 _2395_/Q _1860_/S vssd1 vssd1 vccd1 vccd1 _2395_/D sky130_fd_sc_hd__mux2_1
XFILLER_30_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1789_ _2340_/Q _1804_/A0 _1790_/S vssd1 vssd1 vccd1 vccd1 _2340_/D sky130_fd_sc_hd__mux2_1
XFILLER_1_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1712_ _2278_/Q _1732_/A0 _1715_/S vssd1 vssd1 vccd1 vccd1 _2278_/D sky130_fd_sc_hd__mux2_1
XFILLER_61_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1643_ _2223_/Q _1783_/A0 _1645_/S vssd1 vssd1 vccd1 vccd1 _2223_/D sky130_fd_sc_hd__mux2_1
XANTENNA_1 _1503_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1574_ _1579_/A0 _2168_/Q _1575_/S vssd1 vssd1 vccd1 vccd1 _2168_/D sky130_fd_sc_hd__mux2_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2126_ _2232_/CLK _2126_/D vssd1 vssd1 vccd1 vccd1 _2126_/Q sky130_fd_sc_hd__dfxtp_1
X_2057_ _2094_/CLK _2057_/D vssd1 vssd1 vccd1 vccd1 _2057_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1008_ _1244_/A1 _0999_/Y _1001_/Y _1006_/Y _1007_/Y vssd1 vssd1 vccd1 vccd1 _1009_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_1_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1290_ _2149_/Q _2153_/Q _1292_/S vssd1 vssd1 vccd1 vccd1 _1291_/B sky130_fd_sc_hd__mux2_1
XFILLER_36_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1626_ _1646_/A _1946_/B vssd1 vssd1 vccd1 vccd1 _1630_/S sky130_fd_sc_hd__nor2_4
X_1557_ _2154_/Q _1977_/A0 _1560_/S vssd1 vssd1 vccd1 vccd1 _2154_/D sky130_fd_sc_hd__mux2_1
XFILLER_59_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1488_ _2099_/Q _1503_/A0 _1490_/S vssd1 vssd1 vccd1 vccd1 _2099_/D sky130_fd_sc_hd__mux2_1
XTAP_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2109_ _2113_/CLK _2109_/D vssd1 vssd1 vccd1 vccd1 _2109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2460_ _2461_/CLK _2460_/D vssd1 vssd1 vccd1 vccd1 _2460_/Q sky130_fd_sc_hd__dfxtp_1
X_1411_ _1792_/A1 _2042_/Q _1414_/S vssd1 vssd1 vccd1 vccd1 _2042_/D sky130_fd_sc_hd__mux2_1
X_2391_ _2433_/CLK _2391_/D vssd1 vssd1 vccd1 vccd1 _2391_/Q sky130_fd_sc_hd__dfxtp_1
X_1342_ _2001_/Q _1765_/A0 _1342_/S vssd1 vssd1 vccd1 vccd1 _2001_/D sky130_fd_sc_hd__mux2_1
X_1273_ _2385_/Q _2065_/Q _2105_/Q _2145_/Q _1275_/S0 _1065_/A vssd1 vssd1 vccd1 vccd1
+ _1274_/B sky130_fd_sc_hd__mux4_1
XFILLER_76_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout113 _1979_/A0 vssd1 vssd1 vccd1 vccd1 _1974_/A0 sky130_fd_sc_hd__buf_4
X_1609_ _2196_/Q _1809_/A0 _1610_/S vssd1 vssd1 vccd1 vccd1 _2196_/D sky130_fd_sc_hd__mux2_1
Xfanout102 fanout109/X vssd1 vssd1 vccd1 vccd1 _1940_/A0 sky130_fd_sc_hd__buf_2
Xfanout135 _1475_/A vssd1 vssd1 vccd1 vccd1 _1181_/S sky130_fd_sc_hd__buf_6
Xfanout124 _1739_/A0 vssd1 vssd1 vccd1 vccd1 _1984_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout146 _1233_/S vssd1 vssd1 vccd1 vccd1 _1275_/S0 sky130_fd_sc_hd__buf_8
XFILLER_74_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1960_ _1960_/A0 _2477_/Q _1960_/S vssd1 vssd1 vccd1 vccd1 _2477_/D sky130_fd_sc_hd__mux2_1
X_1891_ _1981_/B _1956_/B vssd1 vssd1 vccd1 vccd1 _1895_/S sky130_fd_sc_hd__nor2_2
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2443_ _2448_/CLK _2443_/D vssd1 vssd1 vccd1 vccd1 _2443_/Q sky130_fd_sc_hd__dfxtp_1
X_2374_ _2482_/CLK _2374_/D vssd1 vssd1 vccd1 vccd1 _2374_/Q sky130_fd_sc_hd__dfxtp_1
X_1325_ _1983_/A1 _1991_/Q _1327_/S vssd1 vssd1 vccd1 vccd1 _1991_/D sky130_fd_sc_hd__mux2_1
XFILLER_56_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1256_ _2405_/Q _2409_/Q _2413_/Q _2417_/Q _1256_/S0 _1256_/S1 vssd1 vssd1 vccd1
+ vccd1 _1256_/X sky130_fd_sc_hd__mux4_1
XFILLER_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1187_ _2340_/Q _1992_/Q _2348_/Q _2352_/Q _1245_/S0 _1409_/B vssd1 vssd1 vccd1 vccd1
+ _1187_/X sky130_fd_sc_hd__mux4_1
XFILLER_64_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1110_ _1237_/A _1105_/X _1244_/A1 vssd1 vssd1 vccd1 vccd1 _1110_/Y sky130_fd_sc_hd__o21ai_1
X_2090_ _2097_/CLK _2090_/D vssd1 vssd1 vccd1 vccd1 _2090_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1041_ _2322_/Q _2326_/Q _2330_/Q _2334_/Q _1275_/S0 _1065_/A vssd1 vssd1 vccd1 vccd1
+ _1041_/X sky130_fd_sc_hd__mux4_2
XFILLER_61_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1943_ _1983_/A1 _2463_/Q _1945_/S vssd1 vssd1 vccd1 vccd1 _2463_/D sky130_fd_sc_hd__mux2_1
X_1874_ _1884_/A0 _2408_/Q _1875_/S vssd1 vssd1 vccd1 vccd1 _2408_/D sky130_fd_sc_hd__mux2_1
X_2426_ _2433_/CLK _2426_/D vssd1 vssd1 vccd1 vccd1 _2426_/Q sky130_fd_sc_hd__dfxtp_1
X_2357_ _2369_/CLK _2357_/D vssd1 vssd1 vccd1 vccd1 _2357_/Q sky130_fd_sc_hd__dfxtp_1
X_2288_ _2481_/CLK _2288_/D vssd1 vssd1 vccd1 vccd1 _2288_/Q sky130_fd_sc_hd__dfxtp_1
X_1308_ input7/X _1268_/X _1282_/Y _1307_/X vssd1 vssd1 vccd1 vccd1 _1308_/X sky130_fd_sc_hd__o2bb2a_2
XFILLER_69_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1239_ _2293_/Q _2297_/Q _1240_/S vssd1 vssd1 vccd1 vccd1 _1239_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1590_ _2181_/Q _1765_/A0 _1590_/S vssd1 vssd1 vccd1 vccd1 _2181_/D sky130_fd_sc_hd__mux2_1
XFILLER_50_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2211_ _2479_/CLK _2211_/D vssd1 vssd1 vccd1 vccd1 _2211_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2142_ _2329_/CLK _2142_/D vssd1 vssd1 vccd1 vccd1 _2142_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2073_ _2335_/CLK _2073_/D vssd1 vssd1 vccd1 vccd1 _2073_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1024_ _1220_/A _1024_/B vssd1 vssd1 vccd1 vccd1 _1360_/B sky130_fd_sc_hd__nand2_4
XFILLER_53_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1926_ _1966_/A _1926_/B vssd1 vssd1 vccd1 vccd1 _1930_/S sky130_fd_sc_hd__nor2_2
X_1857_ _1972_/A0 _2394_/Q _1860_/S vssd1 vssd1 vccd1 vccd1 _2394_/D sky130_fd_sc_hd__mux2_1
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1788_ _2339_/Q _1983_/A1 _1790_/S vssd1 vssd1 vccd1 vccd1 _2339_/D sky130_fd_sc_hd__mux2_1
X_2409_ _2432_/CLK _2409_/D vssd1 vssd1 vccd1 vccd1 _2409_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1711_ _1726_/A _1981_/A vssd1 vssd1 vccd1 vccd1 _1715_/S sky130_fd_sc_hd__nor2_4
X_1642_ _2222_/Q _1742_/A0 _1645_/S vssd1 vssd1 vccd1 vccd1 _2222_/D sky130_fd_sc_hd__mux2_1
XANTENNA_2 _1220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1573_ _1583_/A0 _2167_/Q _1575_/S vssd1 vssd1 vccd1 vccd1 _2167_/D sky130_fd_sc_hd__mux2_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2125_ _2232_/CLK _2125_/D vssd1 vssd1 vccd1 vccd1 _2125_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2056_ _2113_/CLK _2056_/D vssd1 vssd1 vccd1 vccd1 _2056_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1007_ _1220_/A _1002_/X _1024_/B vssd1 vssd1 vccd1 vccd1 _1007_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_34_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1909_ _2436_/Q _1969_/A0 _1910_/S vssd1 vssd1 vccd1 vccd1 _2436_/D sky130_fd_sc_hd__mux2_1
XFILLER_1_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1625_ _1940_/A0 _2209_/Q _1625_/S vssd1 vssd1 vccd1 vccd1 _2209_/D sky130_fd_sc_hd__mux2_1
X_1556_ _1566_/A _1956_/B vssd1 vssd1 vccd1 vccd1 _1560_/S sky130_fd_sc_hd__nor2_4
XTAP_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1487_ _2098_/Q _1777_/A0 _1490_/S vssd1 vssd1 vccd1 vccd1 _2098_/D sky130_fd_sc_hd__mux2_1
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2108_ _2113_/CLK _2108_/D vssd1 vssd1 vccd1 vccd1 _2108_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2039_ _2261_/CLK _2039_/D vssd1 vssd1 vccd1 vccd1 _2039_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_451 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1410_ _1941_/B _1976_/B vssd1 vssd1 vccd1 vccd1 _1414_/S sky130_fd_sc_hd__nand2_2
X_2390_ _2477_/CLK _2390_/D vssd1 vssd1 vccd1 vccd1 _2390_/Q sky130_fd_sc_hd__dfxtp_1
X_1341_ _2000_/Q _1814_/A0 _1342_/S vssd1 vssd1 vccd1 vccd1 _2000_/D sky130_fd_sc_hd__mux2_1
X_1272_ _1100_/A _1269_/X _1271_/X vssd1 vssd1 vccd1 vccd1 _1272_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_24_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1608_ _2195_/Q _1823_/A0 _1610_/S vssd1 vssd1 vccd1 vccd1 _2195_/D sky130_fd_sc_hd__mux2_1
Xfanout103 fanout109/X vssd1 vssd1 vccd1 vccd1 _1505_/A0 sky130_fd_sc_hd__clkbuf_4
X_1539_ _2140_/Q _1579_/A0 _1540_/S vssd1 vssd1 vccd1 vccd1 _2140_/D sky130_fd_sc_hd__mux2_1
Xfanout136 _1182_/S vssd1 vssd1 vccd1 vccd1 _1475_/A sky130_fd_sc_hd__buf_6
Xfanout114 fanout127/X vssd1 vssd1 vccd1 vccd1 _1979_/A0 sky130_fd_sc_hd__clkbuf_4
Xfanout147 fanout148/X vssd1 vssd1 vccd1 vccd1 _1233_/S sky130_fd_sc_hd__buf_6
Xfanout125 _1944_/A0 vssd1 vssd1 vccd1 vccd1 _1739_/A0 sky130_fd_sc_hd__buf_4
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_451 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1890_ _1905_/A0 _2421_/Q _1890_/S vssd1 vssd1 vccd1 vccd1 _2421_/D sky130_fd_sc_hd__mux2_1
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2442_ _2479_/CLK _2442_/D vssd1 vssd1 vccd1 vccd1 _2442_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2373_ _2482_/CLK _2373_/D vssd1 vssd1 vccd1 vccd1 _2373_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1324_ _1822_/A0 _1990_/Q _1327_/S vssd1 vssd1 vccd1 vccd1 _1990_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1255_ _2421_/Q _2025_/Q _2429_/Q _2433_/Q _1256_/S0 _1256_/S1 vssd1 vssd1 vccd1
+ vccd1 _1258_/B sky130_fd_sc_hd__mux4_1
XFILLER_64_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1186_ _2324_/Q _2328_/Q _2332_/Q _2336_/Q _1275_/S0 _1065_/A vssd1 vssd1 vccd1 vccd1
+ _1186_/X sky130_fd_sc_hd__mux4_2
XFILLER_52_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_443 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1040_ input6/X _1040_/B vssd1 vssd1 vccd1 vccd1 _1322_/A sky130_fd_sc_hd__nand2b_4
XFILLER_34_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1942_ _1982_/A1 _2462_/Q _1945_/S vssd1 vssd1 vccd1 vccd1 _2462_/D sky130_fd_sc_hd__mux2_1
X_1873_ _1903_/A0 _2407_/Q _1875_/S vssd1 vssd1 vccd1 vccd1 _2407_/D sky130_fd_sc_hd__mux2_1
X_2425_ _2497_/CLK _2425_/D vssd1 vssd1 vccd1 vccd1 _2425_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2356_ _2368_/CLK _2356_/D vssd1 vssd1 vccd1 vccd1 _2356_/Q sky130_fd_sc_hd__dfxtp_1
X_2287_ _2481_/CLK _2287_/D vssd1 vssd1 vccd1 vccd1 _2287_/Q sky130_fd_sc_hd__dfxtp_1
X_1307_ input7/X _1307_/B _1307_/C _1307_/D vssd1 vssd1 vccd1 vccd1 _1307_/X sky130_fd_sc_hd__or4_1
XFILLER_56_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1238_ _2277_/Q _2281_/Q _2285_/Q _2289_/Q _1181_/S _0992_/A vssd1 vssd1 vccd1 vccd1
+ _1238_/X sky130_fd_sc_hd__mux4_1
XFILLER_56_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1169_ _2436_/Q _2440_/Q _2444_/Q _2448_/Q _1292_/S _1291_/A vssd1 vssd1 vccd1 vccd1
+ _1169_/X sky130_fd_sc_hd__mux4_1
XFILLER_52_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2210_ _2449_/CLK _2210_/D vssd1 vssd1 vccd1 vccd1 _2210_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2141_ _2177_/CLK _2141_/D vssd1 vssd1 vccd1 vccd1 _2141_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2072_ _2349_/CLK _2072_/D vssd1 vssd1 vccd1 vccd1 _2072_/Q sky130_fd_sc_hd__dfxtp_1
X_1023_ _1274_/A _1023_/B vssd1 vssd1 vccd1 vccd1 _1023_/X sky130_fd_sc_hd__and2_2
XFILLER_81_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1925_ _1980_/A0 _2449_/Q _1925_/S vssd1 vssd1 vccd1 vccd1 _2449_/D sky130_fd_sc_hd__mux2_1
X_1856_ _1886_/A _1936_/B vssd1 vssd1 vccd1 vccd1 _1860_/S sky130_fd_sc_hd__or2_4
X_1787_ _2338_/Q _1982_/A1 _1790_/S vssd1 vssd1 vccd1 vccd1 _2338_/D sky130_fd_sc_hd__mux2_1
XFILLER_39_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2408_ _2416_/CLK _2408_/D vssd1 vssd1 vccd1 vccd1 _2408_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2339_ _2495_/CLK _2339_/D vssd1 vssd1 vccd1 vccd1 _2339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1710_ _2277_/Q _1960_/A0 _1710_/S vssd1 vssd1 vccd1 vccd1 _2277_/D sky130_fd_sc_hd__mux2_1
X_1641_ _1641_/A _1981_/B vssd1 vssd1 vccd1 vccd1 _1645_/S sky130_fd_sc_hd__nor2_2
XFILLER_6_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1572_ _1582_/A0 _2166_/Q _1575_/S vssd1 vssd1 vccd1 vccd1 _2166_/D sky130_fd_sc_hd__mux2_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2124_ _2232_/CLK _2124_/D vssd1 vssd1 vccd1 vccd1 _2124_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2055_ _2094_/CLK _2055_/D vssd1 vssd1 vccd1 vccd1 _2055_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1006_ _1174_/A _1004_/X _1005_/X vssd1 vssd1 vccd1 vccd1 _1006_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_22_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1908_ _2435_/Q _1973_/A0 _1910_/S vssd1 vssd1 vccd1 vccd1 _2435_/D sky130_fd_sc_hd__mux2_1
X_1839_ _2380_/Q _1969_/A0 _1840_/S vssd1 vssd1 vccd1 vccd1 _2380_/D sky130_fd_sc_hd__mux2_1
XFILLER_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_37_clk clkbuf_2_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _2477_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_28_clk clkbuf_2_2__f_clk/X vssd1 vssd1 vccd1 vccd1 _2480_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_56_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1624_ _1809_/A0 _2208_/Q _1625_/S vssd1 vssd1 vccd1 vccd1 _2208_/D sky130_fd_sc_hd__mux2_1
X_1555_ _2153_/Q _1980_/A0 _1555_/S vssd1 vssd1 vccd1 vccd1 _2153_/D sky130_fd_sc_hd__mux2_1
X_1486_ _1486_/A _1966_/B vssd1 vssd1 vccd1 vccd1 _1490_/S sky130_fd_sc_hd__nor2_2
XTAP_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2107_ _2113_/CLK _2107_/D vssd1 vssd1 vccd1 vccd1 _2107_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_19_clk clkbuf_2_3__f_clk/X vssd1 vssd1 vccd1 vccd1 _2329_/CLK sky130_fd_sc_hd__clkbuf_16
X_2038_ _2049_/CLK _2038_/D vssd1 vssd1 vccd1 vccd1 _2038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1340_ _1999_/Q _1663_/A0 _1342_/S vssd1 vssd1 vccd1 vccd1 _1999_/D sky130_fd_sc_hd__mux2_1
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1271_ _0992_/Y _1270_/X _1020_/A vssd1 vssd1 vccd1 vccd1 _1271_/X sky130_fd_sc_hd__a21o_1
XFILLER_51_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_8_clk clkbuf_leaf_9_clk/A vssd1 vssd1 vccd1 vccd1 _2367_/CLK sky130_fd_sc_hd__clkbuf_16
X_1607_ _2194_/Q _1917_/A1 _1610_/S vssd1 vssd1 vccd1 vccd1 _2194_/D sky130_fd_sc_hd__mux2_1
Xfanout104 fanout109/X vssd1 vssd1 vccd1 vccd1 _1800_/A0 sky130_fd_sc_hd__clkbuf_4
Xfanout137 fanout148/X vssd1 vssd1 vccd1 vccd1 _1182_/S sky130_fd_sc_hd__buf_6
X_1538_ _2139_/Q _1918_/A1 _1540_/S vssd1 vssd1 vccd1 vccd1 _2139_/D sky130_fd_sc_hd__mux2_1
Xfanout115 _1824_/A0 vssd1 vssd1 vccd1 vccd1 _1814_/A0 sky130_fd_sc_hd__clkbuf_4
Xfanout126 fanout127/X vssd1 vssd1 vccd1 vccd1 _1944_/A0 sky130_fd_sc_hd__clkbuf_4
Xfanout148 input1/X vssd1 vssd1 vccd1 vccd1 fanout148/X sky130_fd_sc_hd__buf_6
X_1469_ _2085_/Q _1800_/A0 _1469_/S vssd1 vssd1 vccd1 vccd1 _2085_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2441_ _2449_/CLK _2441_/D vssd1 vssd1 vccd1 vccd1 _2441_/Q sky130_fd_sc_hd__dfxtp_1
X_2372_ _2485_/CLK _2372_/D vssd1 vssd1 vccd1 vccd1 _2372_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1323_ _1951_/A _1821_/A vssd1 vssd1 vccd1 vccd1 _1327_/S sky130_fd_sc_hd__nand2_2
X_1254_ _1298_/B2 _1252_/X _1253_/X _1295_/B2 vssd1 vssd1 vccd1 vccd1 _1254_/X sky130_fd_sc_hd__a22o_1
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1185_ _1244_/A1 _1180_/X _1184_/X _1176_/X _1178_/X vssd1 vssd1 vccd1 vccd1 _1185_/X
+ sky130_fd_sc_hd__a32o_2
XFILLER_52_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1941_ _1961_/A _1941_/B vssd1 vssd1 vccd1 vccd1 _1945_/S sky130_fd_sc_hd__nand2_2
X_1872_ _1902_/A0 _2406_/Q _1875_/S vssd1 vssd1 vccd1 vccd1 _2406_/D sky130_fd_sc_hd__mux2_1
XFILLER_69_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2424_ _2497_/CLK _2424_/D vssd1 vssd1 vccd1 vccd1 _2424_/Q sky130_fd_sc_hd__dfxtp_1
X_2355_ _2369_/CLK _2355_/D vssd1 vssd1 vccd1 vccd1 _2355_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1306_ _1302_/X _1305_/X _1354_/A vssd1 vssd1 vccd1 vccd1 _1307_/D sky130_fd_sc_hd__o21ba_1
X_2286_ _2296_/CLK _2286_/D vssd1 vssd1 vccd1 vccd1 _2286_/Q sky130_fd_sc_hd__dfxtp_1
X_1237_ _1237_/A _1237_/B vssd1 vssd1 vccd1 vccd1 _1237_/Y sky130_fd_sc_hd__nor2_1
X_1168_ _2484_/Q _2488_/Q _2492_/Q _2032_/Q _1292_/S _1291_/A vssd1 vssd1 vccd1 vccd1
+ _1168_/X sky130_fd_sc_hd__mux4_2
XFILLER_25_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1099_ _2263_/Q _2303_/Q _1277_/S vssd1 vssd1 vccd1 vccd1 _1100_/B sky130_fd_sc_hd__mux2_1
XFILLER_12_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2140_ _2232_/CLK _2140_/D vssd1 vssd1 vccd1 vccd1 _2140_/Q sky130_fd_sc_hd__dfxtp_1
X_2071_ _2335_/CLK _2071_/D vssd1 vssd1 vccd1 vccd1 _2071_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1022_ _2466_/Q _2470_/Q _2474_/Q _2478_/Q _1475_/A _1464_/B vssd1 vssd1 vccd1 vccd1
+ _1022_/X sky130_fd_sc_hd__mux4_1
XFILLER_61_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1924_ _1974_/A0 _2448_/Q _1925_/S vssd1 vssd1 vccd1 vccd1 _2448_/D sky130_fd_sc_hd__mux2_1
X_1855_ _1905_/A0 _2393_/Q _1855_/S vssd1 vssd1 vccd1 vccd1 _2393_/D sky130_fd_sc_hd__mux2_1
X_1786_ _1806_/A _1946_/B vssd1 vssd1 vccd1 vccd1 _1790_/S sky130_fd_sc_hd__nor2_2
X_2407_ _2432_/CLK _2407_/D vssd1 vssd1 vccd1 vccd1 _2407_/Q sky130_fd_sc_hd__dfxtp_1
X_2338_ _2495_/CLK _2338_/D vssd1 vssd1 vccd1 vccd1 _2338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2269_ _2297_/CLK _2269_/D vssd1 vssd1 vccd1 vccd1 _2269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1640_ _1660_/A0 _2221_/Q _1640_/S vssd1 vssd1 vccd1 vccd1 _2221_/D sky130_fd_sc_hd__mux2_1
X_1571_ _1581_/A _1971_/A vssd1 vssd1 vccd1 vccd1 _1575_/S sky130_fd_sc_hd__nand2_4
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2123_ _2176_/CLK _2123_/D vssd1 vssd1 vccd1 vccd1 _2123_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2054_ _2094_/CLK _2054_/D vssd1 vssd1 vccd1 vccd1 _2054_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1005_ _1475_/B _1003_/X _1241_/B1 vssd1 vssd1 vccd1 vccd1 _1005_/X sky130_fd_sc_hd__a21o_1
XFILLER_22_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1907_ _2434_/Q _1972_/A0 _1910_/S vssd1 vssd1 vccd1 vccd1 _2434_/D sky130_fd_sc_hd__mux2_1
X_1838_ _2379_/Q _1973_/A0 _1840_/S vssd1 vssd1 vccd1 vccd1 _2379_/D sky130_fd_sc_hd__mux2_1
X_1769_ _2324_/Q _1804_/A0 _1770_/S vssd1 vssd1 vccd1 vccd1 _2324_/D sky130_fd_sc_hd__mux2_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1623_ _1808_/A0 _2207_/Q _1625_/S vssd1 vssd1 vccd1 vccd1 _2207_/D sky130_fd_sc_hd__mux2_1
X_1554_ _2152_/Q _1974_/A0 _1555_/S vssd1 vssd1 vccd1 vccd1 _2152_/D sky130_fd_sc_hd__mux2_1
X_1485_ _1505_/A0 _2097_/Q _1485_/S vssd1 vssd1 vccd1 vccd1 _2097_/D sky130_fd_sc_hd__mux2_1
.ends

