// This is the unpowered netlist.
module wrapped_tms1x00 (oram_csb,
    ram_csb,
    ram_web,
    wb_clk_i,
    wb_rst_i,
    wbs_we_i,
    io_in,
    io_oeb,
    io_out,
    oram_addr,
    oram_value,
    ram_adrb,
    ram_wmask,
    wbs_adr_i);
 output oram_csb;
 output ram_csb;
 output ram_web;
 input wb_clk_i;
 input wb_rst_i;
 input wbs_we_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 output [8:0] oram_addr;
 input [31:0] oram_value;
 output [8:0] ram_adrb;
 output [3:0] ram_wmask;
 input [31:0] wbs_adr_i;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire net120;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net121;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net122;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net125;
 wire net123;
 wire net124;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net105;
 wire net106;
 wire net107;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net119;
 wire net126;
 wire net127;
 wire net128;
 wire clknet_leaf_0_wb_clk_i;
 wire \tms1x00.A[0] ;
 wire \tms1x00.A[1] ;
 wire \tms1x00.A[2] ;
 wire \tms1x00.A[3] ;
 wire \tms1x00.CL ;
 wire \tms1x00.K_latch[0] ;
 wire \tms1x00.K_latch[1] ;
 wire \tms1x00.K_latch[2] ;
 wire \tms1x00.K_latch[3] ;
 wire \tms1x00.N[0] ;
 wire \tms1x00.N[1] ;
 wire \tms1x00.N[2] ;
 wire \tms1x00.N[3] ;
 wire \tms1x00.PA[0] ;
 wire \tms1x00.PA[1] ;
 wire \tms1x00.PA[2] ;
 wire \tms1x00.PA[3] ;
 wire \tms1x00.PB[0] ;
 wire \tms1x00.PB[1] ;
 wire \tms1x00.PB[2] ;
 wire \tms1x00.PB[3] ;
 wire \tms1x00.PC[0] ;
 wire \tms1x00.PC[1] ;
 wire \tms1x00.PC[2] ;
 wire \tms1x00.PC[3] ;
 wire \tms1x00.PC[4] ;
 wire \tms1x00.PC[5] ;
 wire \tms1x00.P[0] ;
 wire \tms1x00.P[1] ;
 wire \tms1x00.P[2] ;
 wire \tms1x00.P[3] ;
 wire \tms1x00.RAM[0][0] ;
 wire \tms1x00.RAM[0][1] ;
 wire \tms1x00.RAM[0][2] ;
 wire \tms1x00.RAM[0][3] ;
 wire \tms1x00.RAM[100][0] ;
 wire \tms1x00.RAM[100][1] ;
 wire \tms1x00.RAM[100][2] ;
 wire \tms1x00.RAM[100][3] ;
 wire \tms1x00.RAM[101][0] ;
 wire \tms1x00.RAM[101][1] ;
 wire \tms1x00.RAM[101][2] ;
 wire \tms1x00.RAM[101][3] ;
 wire \tms1x00.RAM[102][0] ;
 wire \tms1x00.RAM[102][1] ;
 wire \tms1x00.RAM[102][2] ;
 wire \tms1x00.RAM[102][3] ;
 wire \tms1x00.RAM[103][0] ;
 wire \tms1x00.RAM[103][1] ;
 wire \tms1x00.RAM[103][2] ;
 wire \tms1x00.RAM[103][3] ;
 wire \tms1x00.RAM[104][0] ;
 wire \tms1x00.RAM[104][1] ;
 wire \tms1x00.RAM[104][2] ;
 wire \tms1x00.RAM[104][3] ;
 wire \tms1x00.RAM[105][0] ;
 wire \tms1x00.RAM[105][1] ;
 wire \tms1x00.RAM[105][2] ;
 wire \tms1x00.RAM[105][3] ;
 wire \tms1x00.RAM[106][0] ;
 wire \tms1x00.RAM[106][1] ;
 wire \tms1x00.RAM[106][2] ;
 wire \tms1x00.RAM[106][3] ;
 wire \tms1x00.RAM[107][0] ;
 wire \tms1x00.RAM[107][1] ;
 wire \tms1x00.RAM[107][2] ;
 wire \tms1x00.RAM[107][3] ;
 wire \tms1x00.RAM[108][0] ;
 wire \tms1x00.RAM[108][1] ;
 wire \tms1x00.RAM[108][2] ;
 wire \tms1x00.RAM[108][3] ;
 wire \tms1x00.RAM[109][0] ;
 wire \tms1x00.RAM[109][1] ;
 wire \tms1x00.RAM[109][2] ;
 wire \tms1x00.RAM[109][3] ;
 wire \tms1x00.RAM[10][0] ;
 wire \tms1x00.RAM[10][1] ;
 wire \tms1x00.RAM[10][2] ;
 wire \tms1x00.RAM[10][3] ;
 wire \tms1x00.RAM[110][0] ;
 wire \tms1x00.RAM[110][1] ;
 wire \tms1x00.RAM[110][2] ;
 wire \tms1x00.RAM[110][3] ;
 wire \tms1x00.RAM[111][0] ;
 wire \tms1x00.RAM[111][1] ;
 wire \tms1x00.RAM[111][2] ;
 wire \tms1x00.RAM[111][3] ;
 wire \tms1x00.RAM[112][0] ;
 wire \tms1x00.RAM[112][1] ;
 wire \tms1x00.RAM[112][2] ;
 wire \tms1x00.RAM[112][3] ;
 wire \tms1x00.RAM[113][0] ;
 wire \tms1x00.RAM[113][1] ;
 wire \tms1x00.RAM[113][2] ;
 wire \tms1x00.RAM[113][3] ;
 wire \tms1x00.RAM[114][0] ;
 wire \tms1x00.RAM[114][1] ;
 wire \tms1x00.RAM[114][2] ;
 wire \tms1x00.RAM[114][3] ;
 wire \tms1x00.RAM[115][0] ;
 wire \tms1x00.RAM[115][1] ;
 wire \tms1x00.RAM[115][2] ;
 wire \tms1x00.RAM[115][3] ;
 wire \tms1x00.RAM[116][0] ;
 wire \tms1x00.RAM[116][1] ;
 wire \tms1x00.RAM[116][2] ;
 wire \tms1x00.RAM[116][3] ;
 wire \tms1x00.RAM[117][0] ;
 wire \tms1x00.RAM[117][1] ;
 wire \tms1x00.RAM[117][2] ;
 wire \tms1x00.RAM[117][3] ;
 wire \tms1x00.RAM[118][0] ;
 wire \tms1x00.RAM[118][1] ;
 wire \tms1x00.RAM[118][2] ;
 wire \tms1x00.RAM[118][3] ;
 wire \tms1x00.RAM[119][0] ;
 wire \tms1x00.RAM[119][1] ;
 wire \tms1x00.RAM[119][2] ;
 wire \tms1x00.RAM[119][3] ;
 wire \tms1x00.RAM[11][0] ;
 wire \tms1x00.RAM[11][1] ;
 wire \tms1x00.RAM[11][2] ;
 wire \tms1x00.RAM[11][3] ;
 wire \tms1x00.RAM[120][0] ;
 wire \tms1x00.RAM[120][1] ;
 wire \tms1x00.RAM[120][2] ;
 wire \tms1x00.RAM[120][3] ;
 wire \tms1x00.RAM[121][0] ;
 wire \tms1x00.RAM[121][1] ;
 wire \tms1x00.RAM[121][2] ;
 wire \tms1x00.RAM[121][3] ;
 wire \tms1x00.RAM[122][0] ;
 wire \tms1x00.RAM[122][1] ;
 wire \tms1x00.RAM[122][2] ;
 wire \tms1x00.RAM[122][3] ;
 wire \tms1x00.RAM[123][0] ;
 wire \tms1x00.RAM[123][1] ;
 wire \tms1x00.RAM[123][2] ;
 wire \tms1x00.RAM[123][3] ;
 wire \tms1x00.RAM[124][0] ;
 wire \tms1x00.RAM[124][1] ;
 wire \tms1x00.RAM[124][2] ;
 wire \tms1x00.RAM[124][3] ;
 wire \tms1x00.RAM[125][0] ;
 wire \tms1x00.RAM[125][1] ;
 wire \tms1x00.RAM[125][2] ;
 wire \tms1x00.RAM[125][3] ;
 wire \tms1x00.RAM[126][0] ;
 wire \tms1x00.RAM[126][1] ;
 wire \tms1x00.RAM[126][2] ;
 wire \tms1x00.RAM[126][3] ;
 wire \tms1x00.RAM[127][0] ;
 wire \tms1x00.RAM[127][1] ;
 wire \tms1x00.RAM[127][2] ;
 wire \tms1x00.RAM[127][3] ;
 wire \tms1x00.RAM[12][0] ;
 wire \tms1x00.RAM[12][1] ;
 wire \tms1x00.RAM[12][2] ;
 wire \tms1x00.RAM[12][3] ;
 wire \tms1x00.RAM[13][0] ;
 wire \tms1x00.RAM[13][1] ;
 wire \tms1x00.RAM[13][2] ;
 wire \tms1x00.RAM[13][3] ;
 wire \tms1x00.RAM[14][0] ;
 wire \tms1x00.RAM[14][1] ;
 wire \tms1x00.RAM[14][2] ;
 wire \tms1x00.RAM[14][3] ;
 wire \tms1x00.RAM[15][0] ;
 wire \tms1x00.RAM[15][1] ;
 wire \tms1x00.RAM[15][2] ;
 wire \tms1x00.RAM[15][3] ;
 wire \tms1x00.RAM[16][0] ;
 wire \tms1x00.RAM[16][1] ;
 wire \tms1x00.RAM[16][2] ;
 wire \tms1x00.RAM[16][3] ;
 wire \tms1x00.RAM[17][0] ;
 wire \tms1x00.RAM[17][1] ;
 wire \tms1x00.RAM[17][2] ;
 wire \tms1x00.RAM[17][3] ;
 wire \tms1x00.RAM[18][0] ;
 wire \tms1x00.RAM[18][1] ;
 wire \tms1x00.RAM[18][2] ;
 wire \tms1x00.RAM[18][3] ;
 wire \tms1x00.RAM[19][0] ;
 wire \tms1x00.RAM[19][1] ;
 wire \tms1x00.RAM[19][2] ;
 wire \tms1x00.RAM[19][3] ;
 wire \tms1x00.RAM[1][0] ;
 wire \tms1x00.RAM[1][1] ;
 wire \tms1x00.RAM[1][2] ;
 wire \tms1x00.RAM[1][3] ;
 wire \tms1x00.RAM[20][0] ;
 wire \tms1x00.RAM[20][1] ;
 wire \tms1x00.RAM[20][2] ;
 wire \tms1x00.RAM[20][3] ;
 wire \tms1x00.RAM[21][0] ;
 wire \tms1x00.RAM[21][1] ;
 wire \tms1x00.RAM[21][2] ;
 wire \tms1x00.RAM[21][3] ;
 wire \tms1x00.RAM[22][0] ;
 wire \tms1x00.RAM[22][1] ;
 wire \tms1x00.RAM[22][2] ;
 wire \tms1x00.RAM[22][3] ;
 wire \tms1x00.RAM[23][0] ;
 wire \tms1x00.RAM[23][1] ;
 wire \tms1x00.RAM[23][2] ;
 wire \tms1x00.RAM[23][3] ;
 wire \tms1x00.RAM[24][0] ;
 wire \tms1x00.RAM[24][1] ;
 wire \tms1x00.RAM[24][2] ;
 wire \tms1x00.RAM[24][3] ;
 wire \tms1x00.RAM[25][0] ;
 wire \tms1x00.RAM[25][1] ;
 wire \tms1x00.RAM[25][2] ;
 wire \tms1x00.RAM[25][3] ;
 wire \tms1x00.RAM[26][0] ;
 wire \tms1x00.RAM[26][1] ;
 wire \tms1x00.RAM[26][2] ;
 wire \tms1x00.RAM[26][3] ;
 wire \tms1x00.RAM[27][0] ;
 wire \tms1x00.RAM[27][1] ;
 wire \tms1x00.RAM[27][2] ;
 wire \tms1x00.RAM[27][3] ;
 wire \tms1x00.RAM[28][0] ;
 wire \tms1x00.RAM[28][1] ;
 wire \tms1x00.RAM[28][2] ;
 wire \tms1x00.RAM[28][3] ;
 wire \tms1x00.RAM[29][0] ;
 wire \tms1x00.RAM[29][1] ;
 wire \tms1x00.RAM[29][2] ;
 wire \tms1x00.RAM[29][3] ;
 wire \tms1x00.RAM[2][0] ;
 wire \tms1x00.RAM[2][1] ;
 wire \tms1x00.RAM[2][2] ;
 wire \tms1x00.RAM[2][3] ;
 wire \tms1x00.RAM[30][0] ;
 wire \tms1x00.RAM[30][1] ;
 wire \tms1x00.RAM[30][2] ;
 wire \tms1x00.RAM[30][3] ;
 wire \tms1x00.RAM[31][0] ;
 wire \tms1x00.RAM[31][1] ;
 wire \tms1x00.RAM[31][2] ;
 wire \tms1x00.RAM[31][3] ;
 wire \tms1x00.RAM[32][0] ;
 wire \tms1x00.RAM[32][1] ;
 wire \tms1x00.RAM[32][2] ;
 wire \tms1x00.RAM[32][3] ;
 wire \tms1x00.RAM[33][0] ;
 wire \tms1x00.RAM[33][1] ;
 wire \tms1x00.RAM[33][2] ;
 wire \tms1x00.RAM[33][3] ;
 wire \tms1x00.RAM[34][0] ;
 wire \tms1x00.RAM[34][1] ;
 wire \tms1x00.RAM[34][2] ;
 wire \tms1x00.RAM[34][3] ;
 wire \tms1x00.RAM[35][0] ;
 wire \tms1x00.RAM[35][1] ;
 wire \tms1x00.RAM[35][2] ;
 wire \tms1x00.RAM[35][3] ;
 wire \tms1x00.RAM[36][0] ;
 wire \tms1x00.RAM[36][1] ;
 wire \tms1x00.RAM[36][2] ;
 wire \tms1x00.RAM[36][3] ;
 wire \tms1x00.RAM[37][0] ;
 wire \tms1x00.RAM[37][1] ;
 wire \tms1x00.RAM[37][2] ;
 wire \tms1x00.RAM[37][3] ;
 wire \tms1x00.RAM[38][0] ;
 wire \tms1x00.RAM[38][1] ;
 wire \tms1x00.RAM[38][2] ;
 wire \tms1x00.RAM[38][3] ;
 wire \tms1x00.RAM[39][0] ;
 wire \tms1x00.RAM[39][1] ;
 wire \tms1x00.RAM[39][2] ;
 wire \tms1x00.RAM[39][3] ;
 wire \tms1x00.RAM[3][0] ;
 wire \tms1x00.RAM[3][1] ;
 wire \tms1x00.RAM[3][2] ;
 wire \tms1x00.RAM[3][3] ;
 wire \tms1x00.RAM[40][0] ;
 wire \tms1x00.RAM[40][1] ;
 wire \tms1x00.RAM[40][2] ;
 wire \tms1x00.RAM[40][3] ;
 wire \tms1x00.RAM[41][0] ;
 wire \tms1x00.RAM[41][1] ;
 wire \tms1x00.RAM[41][2] ;
 wire \tms1x00.RAM[41][3] ;
 wire \tms1x00.RAM[42][0] ;
 wire \tms1x00.RAM[42][1] ;
 wire \tms1x00.RAM[42][2] ;
 wire \tms1x00.RAM[42][3] ;
 wire \tms1x00.RAM[43][0] ;
 wire \tms1x00.RAM[43][1] ;
 wire \tms1x00.RAM[43][2] ;
 wire \tms1x00.RAM[43][3] ;
 wire \tms1x00.RAM[44][0] ;
 wire \tms1x00.RAM[44][1] ;
 wire \tms1x00.RAM[44][2] ;
 wire \tms1x00.RAM[44][3] ;
 wire \tms1x00.RAM[45][0] ;
 wire \tms1x00.RAM[45][1] ;
 wire \tms1x00.RAM[45][2] ;
 wire \tms1x00.RAM[45][3] ;
 wire \tms1x00.RAM[46][0] ;
 wire \tms1x00.RAM[46][1] ;
 wire \tms1x00.RAM[46][2] ;
 wire \tms1x00.RAM[46][3] ;
 wire \tms1x00.RAM[47][0] ;
 wire \tms1x00.RAM[47][1] ;
 wire \tms1x00.RAM[47][2] ;
 wire \tms1x00.RAM[47][3] ;
 wire \tms1x00.RAM[48][0] ;
 wire \tms1x00.RAM[48][1] ;
 wire \tms1x00.RAM[48][2] ;
 wire \tms1x00.RAM[48][3] ;
 wire \tms1x00.RAM[49][0] ;
 wire \tms1x00.RAM[49][1] ;
 wire \tms1x00.RAM[49][2] ;
 wire \tms1x00.RAM[49][3] ;
 wire \tms1x00.RAM[4][0] ;
 wire \tms1x00.RAM[4][1] ;
 wire \tms1x00.RAM[4][2] ;
 wire \tms1x00.RAM[4][3] ;
 wire \tms1x00.RAM[50][0] ;
 wire \tms1x00.RAM[50][1] ;
 wire \tms1x00.RAM[50][2] ;
 wire \tms1x00.RAM[50][3] ;
 wire \tms1x00.RAM[51][0] ;
 wire \tms1x00.RAM[51][1] ;
 wire \tms1x00.RAM[51][2] ;
 wire \tms1x00.RAM[51][3] ;
 wire \tms1x00.RAM[52][0] ;
 wire \tms1x00.RAM[52][1] ;
 wire \tms1x00.RAM[52][2] ;
 wire \tms1x00.RAM[52][3] ;
 wire \tms1x00.RAM[53][0] ;
 wire \tms1x00.RAM[53][1] ;
 wire \tms1x00.RAM[53][2] ;
 wire \tms1x00.RAM[53][3] ;
 wire \tms1x00.RAM[54][0] ;
 wire \tms1x00.RAM[54][1] ;
 wire \tms1x00.RAM[54][2] ;
 wire \tms1x00.RAM[54][3] ;
 wire \tms1x00.RAM[55][0] ;
 wire \tms1x00.RAM[55][1] ;
 wire \tms1x00.RAM[55][2] ;
 wire \tms1x00.RAM[55][3] ;
 wire \tms1x00.RAM[56][0] ;
 wire \tms1x00.RAM[56][1] ;
 wire \tms1x00.RAM[56][2] ;
 wire \tms1x00.RAM[56][3] ;
 wire \tms1x00.RAM[57][0] ;
 wire \tms1x00.RAM[57][1] ;
 wire \tms1x00.RAM[57][2] ;
 wire \tms1x00.RAM[57][3] ;
 wire \tms1x00.RAM[58][0] ;
 wire \tms1x00.RAM[58][1] ;
 wire \tms1x00.RAM[58][2] ;
 wire \tms1x00.RAM[58][3] ;
 wire \tms1x00.RAM[59][0] ;
 wire \tms1x00.RAM[59][1] ;
 wire \tms1x00.RAM[59][2] ;
 wire \tms1x00.RAM[59][3] ;
 wire \tms1x00.RAM[5][0] ;
 wire \tms1x00.RAM[5][1] ;
 wire \tms1x00.RAM[5][2] ;
 wire \tms1x00.RAM[5][3] ;
 wire \tms1x00.RAM[60][0] ;
 wire \tms1x00.RAM[60][1] ;
 wire \tms1x00.RAM[60][2] ;
 wire \tms1x00.RAM[60][3] ;
 wire \tms1x00.RAM[61][0] ;
 wire \tms1x00.RAM[61][1] ;
 wire \tms1x00.RAM[61][2] ;
 wire \tms1x00.RAM[61][3] ;
 wire \tms1x00.RAM[62][0] ;
 wire \tms1x00.RAM[62][1] ;
 wire \tms1x00.RAM[62][2] ;
 wire \tms1x00.RAM[62][3] ;
 wire \tms1x00.RAM[63][0] ;
 wire \tms1x00.RAM[63][1] ;
 wire \tms1x00.RAM[63][2] ;
 wire \tms1x00.RAM[63][3] ;
 wire \tms1x00.RAM[64][0] ;
 wire \tms1x00.RAM[64][1] ;
 wire \tms1x00.RAM[64][2] ;
 wire \tms1x00.RAM[64][3] ;
 wire \tms1x00.RAM[65][0] ;
 wire \tms1x00.RAM[65][1] ;
 wire \tms1x00.RAM[65][2] ;
 wire \tms1x00.RAM[65][3] ;
 wire \tms1x00.RAM[66][0] ;
 wire \tms1x00.RAM[66][1] ;
 wire \tms1x00.RAM[66][2] ;
 wire \tms1x00.RAM[66][3] ;
 wire \tms1x00.RAM[67][0] ;
 wire \tms1x00.RAM[67][1] ;
 wire \tms1x00.RAM[67][2] ;
 wire \tms1x00.RAM[67][3] ;
 wire \tms1x00.RAM[68][0] ;
 wire \tms1x00.RAM[68][1] ;
 wire \tms1x00.RAM[68][2] ;
 wire \tms1x00.RAM[68][3] ;
 wire \tms1x00.RAM[69][0] ;
 wire \tms1x00.RAM[69][1] ;
 wire \tms1x00.RAM[69][2] ;
 wire \tms1x00.RAM[69][3] ;
 wire \tms1x00.RAM[6][0] ;
 wire \tms1x00.RAM[6][1] ;
 wire \tms1x00.RAM[6][2] ;
 wire \tms1x00.RAM[6][3] ;
 wire \tms1x00.RAM[70][0] ;
 wire \tms1x00.RAM[70][1] ;
 wire \tms1x00.RAM[70][2] ;
 wire \tms1x00.RAM[70][3] ;
 wire \tms1x00.RAM[71][0] ;
 wire \tms1x00.RAM[71][1] ;
 wire \tms1x00.RAM[71][2] ;
 wire \tms1x00.RAM[71][3] ;
 wire \tms1x00.RAM[72][0] ;
 wire \tms1x00.RAM[72][1] ;
 wire \tms1x00.RAM[72][2] ;
 wire \tms1x00.RAM[72][3] ;
 wire \tms1x00.RAM[73][0] ;
 wire \tms1x00.RAM[73][1] ;
 wire \tms1x00.RAM[73][2] ;
 wire \tms1x00.RAM[73][3] ;
 wire \tms1x00.RAM[74][0] ;
 wire \tms1x00.RAM[74][1] ;
 wire \tms1x00.RAM[74][2] ;
 wire \tms1x00.RAM[74][3] ;
 wire \tms1x00.RAM[75][0] ;
 wire \tms1x00.RAM[75][1] ;
 wire \tms1x00.RAM[75][2] ;
 wire \tms1x00.RAM[75][3] ;
 wire \tms1x00.RAM[76][0] ;
 wire \tms1x00.RAM[76][1] ;
 wire \tms1x00.RAM[76][2] ;
 wire \tms1x00.RAM[76][3] ;
 wire \tms1x00.RAM[77][0] ;
 wire \tms1x00.RAM[77][1] ;
 wire \tms1x00.RAM[77][2] ;
 wire \tms1x00.RAM[77][3] ;
 wire \tms1x00.RAM[78][0] ;
 wire \tms1x00.RAM[78][1] ;
 wire \tms1x00.RAM[78][2] ;
 wire \tms1x00.RAM[78][3] ;
 wire \tms1x00.RAM[79][0] ;
 wire \tms1x00.RAM[79][1] ;
 wire \tms1x00.RAM[79][2] ;
 wire \tms1x00.RAM[79][3] ;
 wire \tms1x00.RAM[7][0] ;
 wire \tms1x00.RAM[7][1] ;
 wire \tms1x00.RAM[7][2] ;
 wire \tms1x00.RAM[7][3] ;
 wire \tms1x00.RAM[80][0] ;
 wire \tms1x00.RAM[80][1] ;
 wire \tms1x00.RAM[80][2] ;
 wire \tms1x00.RAM[80][3] ;
 wire \tms1x00.RAM[81][0] ;
 wire \tms1x00.RAM[81][1] ;
 wire \tms1x00.RAM[81][2] ;
 wire \tms1x00.RAM[81][3] ;
 wire \tms1x00.RAM[82][0] ;
 wire \tms1x00.RAM[82][1] ;
 wire \tms1x00.RAM[82][2] ;
 wire \tms1x00.RAM[82][3] ;
 wire \tms1x00.RAM[83][0] ;
 wire \tms1x00.RAM[83][1] ;
 wire \tms1x00.RAM[83][2] ;
 wire \tms1x00.RAM[83][3] ;
 wire \tms1x00.RAM[84][0] ;
 wire \tms1x00.RAM[84][1] ;
 wire \tms1x00.RAM[84][2] ;
 wire \tms1x00.RAM[84][3] ;
 wire \tms1x00.RAM[85][0] ;
 wire \tms1x00.RAM[85][1] ;
 wire \tms1x00.RAM[85][2] ;
 wire \tms1x00.RAM[85][3] ;
 wire \tms1x00.RAM[86][0] ;
 wire \tms1x00.RAM[86][1] ;
 wire \tms1x00.RAM[86][2] ;
 wire \tms1x00.RAM[86][3] ;
 wire \tms1x00.RAM[87][0] ;
 wire \tms1x00.RAM[87][1] ;
 wire \tms1x00.RAM[87][2] ;
 wire \tms1x00.RAM[87][3] ;
 wire \tms1x00.RAM[88][0] ;
 wire \tms1x00.RAM[88][1] ;
 wire \tms1x00.RAM[88][2] ;
 wire \tms1x00.RAM[88][3] ;
 wire \tms1x00.RAM[89][0] ;
 wire \tms1x00.RAM[89][1] ;
 wire \tms1x00.RAM[89][2] ;
 wire \tms1x00.RAM[89][3] ;
 wire \tms1x00.RAM[8][0] ;
 wire \tms1x00.RAM[8][1] ;
 wire \tms1x00.RAM[8][2] ;
 wire \tms1x00.RAM[8][3] ;
 wire \tms1x00.RAM[90][0] ;
 wire \tms1x00.RAM[90][1] ;
 wire \tms1x00.RAM[90][2] ;
 wire \tms1x00.RAM[90][3] ;
 wire \tms1x00.RAM[91][0] ;
 wire \tms1x00.RAM[91][1] ;
 wire \tms1x00.RAM[91][2] ;
 wire \tms1x00.RAM[91][3] ;
 wire \tms1x00.RAM[92][0] ;
 wire \tms1x00.RAM[92][1] ;
 wire \tms1x00.RAM[92][2] ;
 wire \tms1x00.RAM[92][3] ;
 wire \tms1x00.RAM[93][0] ;
 wire \tms1x00.RAM[93][1] ;
 wire \tms1x00.RAM[93][2] ;
 wire \tms1x00.RAM[93][3] ;
 wire \tms1x00.RAM[94][0] ;
 wire \tms1x00.RAM[94][1] ;
 wire \tms1x00.RAM[94][2] ;
 wire \tms1x00.RAM[94][3] ;
 wire \tms1x00.RAM[95][0] ;
 wire \tms1x00.RAM[95][1] ;
 wire \tms1x00.RAM[95][2] ;
 wire \tms1x00.RAM[95][3] ;
 wire \tms1x00.RAM[96][0] ;
 wire \tms1x00.RAM[96][1] ;
 wire \tms1x00.RAM[96][2] ;
 wire \tms1x00.RAM[96][3] ;
 wire \tms1x00.RAM[97][0] ;
 wire \tms1x00.RAM[97][1] ;
 wire \tms1x00.RAM[97][2] ;
 wire \tms1x00.RAM[97][3] ;
 wire \tms1x00.RAM[98][0] ;
 wire \tms1x00.RAM[98][1] ;
 wire \tms1x00.RAM[98][2] ;
 wire \tms1x00.RAM[98][3] ;
 wire \tms1x00.RAM[99][0] ;
 wire \tms1x00.RAM[99][1] ;
 wire \tms1x00.RAM[99][2] ;
 wire \tms1x00.RAM[99][3] ;
 wire \tms1x00.RAM[9][0] ;
 wire \tms1x00.RAM[9][1] ;
 wire \tms1x00.RAM[9][2] ;
 wire \tms1x00.RAM[9][3] ;
 wire \tms1x00.SR[0] ;
 wire \tms1x00.SR[1] ;
 wire \tms1x00.SR[2] ;
 wire \tms1x00.SR[3] ;
 wire \tms1x00.SR[4] ;
 wire \tms1x00.SR[5] ;
 wire \tms1x00.X[0] ;
 wire \tms1x00.X[1] ;
 wire \tms1x00.X[2] ;
 wire \tms1x00.Y[0] ;
 wire \tms1x00.Y[1] ;
 wire \tms1x00.Y[2] ;
 wire \tms1x00.Y[3] ;
 wire \tms1x00.ins_in[0] ;
 wire \tms1x00.ins_in[1] ;
 wire \tms1x00.ins_in[2] ;
 wire \tms1x00.ins_in[3] ;
 wire \tms1x00.ins_in[4] ;
 wire \tms1x00.ins_in[5] ;
 wire \tms1x00.ins_in[6] ;
 wire \tms1x00.ins_in[7] ;
 wire \tms1x00.ram_addr_buff[0] ;
 wire \tms1x00.ram_addr_buff[1] ;
 wire \tms1x00.ram_addr_buff[2] ;
 wire \tms1x00.ram_addr_buff[3] ;
 wire \tms1x00.ram_addr_buff[4] ;
 wire \tms1x00.ram_addr_buff[5] ;
 wire \tms1x00.ram_addr_buff[6] ;
 wire \tms1x00.rom_addr[0] ;
 wire \tms1x00.rom_addr[1] ;
 wire \tms1x00.status ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire clknet_leaf_1_wb_clk_i;
 wire clknet_leaf_2_wb_clk_i;
 wire clknet_leaf_3_wb_clk_i;
 wire clknet_leaf_4_wb_clk_i;
 wire clknet_leaf_5_wb_clk_i;
 wire clknet_leaf_6_wb_clk_i;
 wire clknet_leaf_7_wb_clk_i;
 wire clknet_leaf_8_wb_clk_i;
 wire clknet_leaf_9_wb_clk_i;
 wire clknet_leaf_10_wb_clk_i;
 wire clknet_leaf_11_wb_clk_i;
 wire clknet_leaf_12_wb_clk_i;
 wire clknet_leaf_13_wb_clk_i;
 wire clknet_leaf_14_wb_clk_i;
 wire clknet_leaf_15_wb_clk_i;
 wire clknet_leaf_16_wb_clk_i;
 wire clknet_leaf_17_wb_clk_i;
 wire clknet_leaf_18_wb_clk_i;
 wire clknet_leaf_19_wb_clk_i;
 wire clknet_leaf_20_wb_clk_i;
 wire clknet_leaf_21_wb_clk_i;
 wire clknet_leaf_22_wb_clk_i;
 wire clknet_leaf_23_wb_clk_i;
 wire clknet_leaf_24_wb_clk_i;
 wire clknet_leaf_25_wb_clk_i;
 wire clknet_leaf_26_wb_clk_i;
 wire clknet_leaf_27_wb_clk_i;
 wire clknet_leaf_28_wb_clk_i;
 wire clknet_leaf_29_wb_clk_i;
 wire clknet_leaf_30_wb_clk_i;
 wire clknet_leaf_31_wb_clk_i;
 wire clknet_leaf_32_wb_clk_i;
 wire clknet_leaf_33_wb_clk_i;
 wire clknet_leaf_34_wb_clk_i;
 wire clknet_leaf_35_wb_clk_i;
 wire clknet_leaf_37_wb_clk_i;
 wire clknet_0_wb_clk_i;
 wire clknet_2_0__leaf_wb_clk_i;
 wire clknet_2_1__leaf_wb_clk_i;
 wire clknet_2_2__leaf_wb_clk_i;
 wire clknet_2_3__leaf_wb_clk_i;

 sky130_fd_sc_hd__buf_2 _2074_ (.A(\tms1x00.Y[0] ),
    .X(_0616_));
 sky130_fd_sc_hd__buf_2 _2075_ (.A(\tms1x00.ram_addr_buff[0] ),
    .X(_0617_));
 sky130_fd_sc_hd__inv_2 _2076_ (.A(net16),
    .Y(_0618_));
 sky130_fd_sc_hd__nand2b_1 _2077_ (.A_N(net33),
    .B(net35),
    .Y(_0619_));
 sky130_fd_sc_hd__nor2_4 _2078_ (.A(net34),
    .B(_0619_),
    .Y(_0620_));
 sky130_fd_sc_hd__nand2_2 _2079_ (.A(_0618_),
    .B(_0620_),
    .Y(_0621_));
 sky130_fd_sc_hd__buf_4 _2080_ (.A(_0621_),
    .X(_0622_));
 sky130_fd_sc_hd__mux2_1 _2081_ (.A0(_0616_),
    .A1(_0617_),
    .S(_0622_),
    .X(_0623_));
 sky130_fd_sc_hd__clkbuf_1 _2082_ (.A(_0623_),
    .X(_0007_));
 sky130_fd_sc_hd__buf_2 _2083_ (.A(\tms1x00.Y[1] ),
    .X(_0624_));
 sky130_fd_sc_hd__buf_2 _2084_ (.A(\tms1x00.ram_addr_buff[1] ),
    .X(_0625_));
 sky130_fd_sc_hd__mux2_1 _2085_ (.A0(_0624_),
    .A1(_0625_),
    .S(_0622_),
    .X(_0626_));
 sky130_fd_sc_hd__clkbuf_1 _2086_ (.A(_0626_),
    .X(_0008_));
 sky130_fd_sc_hd__buf_2 _2087_ (.A(\tms1x00.Y[2] ),
    .X(_0627_));
 sky130_fd_sc_hd__mux2_1 _2088_ (.A0(_0627_),
    .A1(\tms1x00.ram_addr_buff[2] ),
    .S(_0622_),
    .X(_0628_));
 sky130_fd_sc_hd__clkbuf_1 _2089_ (.A(_0628_),
    .X(_0009_));
 sky130_fd_sc_hd__clkbuf_4 _2090_ (.A(\tms1x00.Y[3] ),
    .X(_0629_));
 sky130_fd_sc_hd__clkbuf_4 _2091_ (.A(_0629_),
    .X(_0630_));
 sky130_fd_sc_hd__mux2_1 _2092_ (.A0(_0630_),
    .A1(\tms1x00.ram_addr_buff[3] ),
    .S(_0622_),
    .X(_0631_));
 sky130_fd_sc_hd__clkbuf_1 _2093_ (.A(_0631_),
    .X(_0010_));
 sky130_fd_sc_hd__mux2_1 _2094_ (.A0(\tms1x00.X[2] ),
    .A1(\tms1x00.ram_addr_buff[4] ),
    .S(_0622_),
    .X(_0632_));
 sky130_fd_sc_hd__clkbuf_1 _2095_ (.A(_0632_),
    .X(_0011_));
 sky130_fd_sc_hd__mux2_1 _2096_ (.A0(\tms1x00.X[0] ),
    .A1(\tms1x00.ram_addr_buff[5] ),
    .S(_0622_),
    .X(_0633_));
 sky130_fd_sc_hd__clkbuf_1 _2097_ (.A(_0633_),
    .X(_0012_));
 sky130_fd_sc_hd__mux2_1 _2098_ (.A0(\tms1x00.X[1] ),
    .A1(\tms1x00.ram_addr_buff[6] ),
    .S(_0622_),
    .X(_0634_));
 sky130_fd_sc_hd__clkbuf_1 _2099_ (.A(_0634_),
    .X(_0013_));
 sky130_fd_sc_hd__inv_2 _2100_ (.A(net18),
    .Y(net70));
 sky130_fd_sc_hd__inv_2 _2101_ (.A(net27),
    .Y(net71));
 sky130_fd_sc_hd__or3_1 _2102_ (.A(_0627_),
    .B(_0624_),
    .C(_0616_),
    .X(_0635_));
 sky130_fd_sc_hd__clkbuf_4 _2103_ (.A(\tms1x00.ins_in[7] ),
    .X(_0636_));
 sky130_fd_sc_hd__clkbuf_4 _2104_ (.A(\tms1x00.ins_in[6] ),
    .X(_0637_));
 sky130_fd_sc_hd__or4_1 _2105_ (.A(\tms1x00.ins_in[3] ),
    .B(\tms1x00.ins_in[2] ),
    .C(\tms1x00.ins_in[1] ),
    .D(\tms1x00.ins_in[0] ),
    .X(_0638_));
 sky130_fd_sc_hd__nand2_1 _2106_ (.A(\tms1x00.ins_in[5] ),
    .B(\tms1x00.ins_in[4] ),
    .Y(_0639_));
 sky130_fd_sc_hd__or2_2 _2107_ (.A(_0638_),
    .B(_0639_),
    .X(_0640_));
 sky130_fd_sc_hd__nand3b_2 _2108_ (.A_N(net35),
    .B(net33),
    .C(net34),
    .Y(_0641_));
 sky130_fd_sc_hd__or4_4 _2109_ (.A(_0636_),
    .B(_0637_),
    .C(_0640_),
    .D(_0641_),
    .X(_0642_));
 sky130_fd_sc_hd__buf_2 _2110_ (.A(_0642_),
    .X(_0643_));
 sky130_fd_sc_hd__inv_2 _2111_ (.A(\tms1x00.Y[3] ),
    .Y(_0644_));
 sky130_fd_sc_hd__buf_2 _2112_ (.A(_0644_),
    .X(_0645_));
 sky130_fd_sc_hd__nor3_1 _2113_ (.A(_0627_),
    .B(_0624_),
    .C(_0616_),
    .Y(_0646_));
 sky130_fd_sc_hd__or2b_1 _2114_ (.A(\tms1x00.ins_in[6] ),
    .B_N(\tms1x00.ins_in[7] ),
    .X(_0647_));
 sky130_fd_sc_hd__or2_2 _2115_ (.A(_0641_),
    .B(_0647_),
    .X(_0648_));
 sky130_fd_sc_hd__nor2_4 _2116_ (.A(_0640_),
    .B(_0648_),
    .Y(_0649_));
 sky130_fd_sc_hd__buf_2 _2117_ (.A(_0649_),
    .X(_0650_));
 sky130_fd_sc_hd__a31o_1 _2118_ (.A1(_0645_),
    .A2(_0646_),
    .A3(_0650_),
    .B1(net36),
    .X(_0651_));
 sky130_fd_sc_hd__clkbuf_4 _2119_ (.A(_0618_),
    .X(_0652_));
 sky130_fd_sc_hd__o311a_1 _2120_ (.A1(_0630_),
    .A2(_0635_),
    .A3(_0643_),
    .B1(_0651_),
    .C1(_0652_),
    .X(_0014_));
 sky130_fd_sc_hd__and4b_1 _2121_ (.A_N(\tms1x00.ins_in[5] ),
    .B(\tms1x00.ins_in[4] ),
    .C(\tms1x00.ins_in[7] ),
    .D(\tms1x00.ins_in[6] ),
    .X(_0653_));
 sky130_fd_sc_hd__nand3b_1 _2122_ (.A_N(\tms1x00.ins_in[3] ),
    .B(\tms1x00.ins_in[2] ),
    .C(_0653_),
    .Y(_0654_));
 sky130_fd_sc_hd__or3b_1 _2123_ (.A(\tms1x00.ins_in[1] ),
    .B(net33),
    .C_N(net34),
    .X(_0655_));
 sky130_fd_sc_hd__or4_2 _2124_ (.A(net35),
    .B(net16),
    .C(_0654_),
    .D(_0655_),
    .X(_0656_));
 sky130_fd_sc_hd__clkbuf_4 _2125_ (.A(_0005_),
    .X(_0657_));
 sky130_fd_sc_hd__buf_4 _2126_ (.A(_0001_),
    .X(_0658_));
 sky130_fd_sc_hd__clkbuf_4 _2127_ (.A(_0658_),
    .X(_0659_));
 sky130_fd_sc_hd__clkbuf_4 _2128_ (.A(_0659_),
    .X(_0660_));
 sky130_fd_sc_hd__buf_6 _2129_ (.A(_0000_),
    .X(_0661_));
 sky130_fd_sc_hd__mux2_1 _2130_ (.A0(\tms1x00.RAM[92][0] ),
    .A1(\tms1x00.RAM[93][0] ),
    .S(_0661_),
    .X(_0662_));
 sky130_fd_sc_hd__inv_2 _2131_ (.A(_0662_),
    .Y(_0663_));
 sky130_fd_sc_hd__clkbuf_4 _2132_ (.A(_0659_),
    .X(_0664_));
 sky130_fd_sc_hd__buf_6 _2133_ (.A(_0000_),
    .X(_0665_));
 sky130_fd_sc_hd__buf_6 _2134_ (.A(_0665_),
    .X(_0666_));
 sky130_fd_sc_hd__mux2_1 _2135_ (.A0(\tms1x00.RAM[94][0] ),
    .A1(\tms1x00.RAM[95][0] ),
    .S(_0666_),
    .X(_0667_));
 sky130_fd_sc_hd__nand2_1 _2136_ (.A(_0664_),
    .B(_0667_),
    .Y(_0668_));
 sky130_fd_sc_hd__clkbuf_4 _2137_ (.A(_0002_),
    .X(_0669_));
 sky130_fd_sc_hd__o211a_1 _2138_ (.A1(_0660_),
    .A2(_0663_),
    .B1(_0668_),
    .C1(_0669_),
    .X(_0670_));
 sky130_fd_sc_hd__buf_2 _2139_ (.A(_0002_),
    .X(_0671_));
 sky130_fd_sc_hd__clkbuf_4 _2140_ (.A(_0671_),
    .X(_0672_));
 sky130_fd_sc_hd__buf_6 _2141_ (.A(_0665_),
    .X(_0673_));
 sky130_fd_sc_hd__buf_4 _2142_ (.A(_0658_),
    .X(_0674_));
 sky130_fd_sc_hd__mux4_1 _2143_ (.A0(\tms1x00.RAM[88][0] ),
    .A1(\tms1x00.RAM[89][0] ),
    .A2(\tms1x00.RAM[90][0] ),
    .A3(\tms1x00.RAM[91][0] ),
    .S0(_0673_),
    .S1(_0674_),
    .X(_0675_));
 sky130_fd_sc_hd__clkbuf_4 _2144_ (.A(_0003_),
    .X(_0676_));
 sky130_fd_sc_hd__o21ai_1 _2145_ (.A1(_0672_),
    .A2(_0675_),
    .B1(_0676_),
    .Y(_0677_));
 sky130_fd_sc_hd__clkbuf_4 _2146_ (.A(_0671_),
    .X(_0678_));
 sky130_fd_sc_hd__buf_6 _2147_ (.A(_0000_),
    .X(_0679_));
 sky130_fd_sc_hd__buf_6 _2148_ (.A(_0679_),
    .X(_0680_));
 sky130_fd_sc_hd__buf_6 _2149_ (.A(_0001_),
    .X(_0681_));
 sky130_fd_sc_hd__buf_6 _2150_ (.A(_0681_),
    .X(_0682_));
 sky130_fd_sc_hd__mux4_1 _2151_ (.A0(\tms1x00.RAM[80][0] ),
    .A1(\tms1x00.RAM[81][0] ),
    .A2(\tms1x00.RAM[82][0] ),
    .A3(\tms1x00.RAM[83][0] ),
    .S0(_0680_),
    .S1(_0682_),
    .X(_0683_));
 sky130_fd_sc_hd__nor2_1 _2152_ (.A(_0678_),
    .B(_0683_),
    .Y(_0684_));
 sky130_fd_sc_hd__inv_2 _2153_ (.A(_0002_),
    .Y(_0685_));
 sky130_fd_sc_hd__clkbuf_4 _2154_ (.A(_0685_),
    .X(_0686_));
 sky130_fd_sc_hd__buf_4 _2155_ (.A(_0661_),
    .X(_0687_));
 sky130_fd_sc_hd__buf_4 _2156_ (.A(_0658_),
    .X(_0688_));
 sky130_fd_sc_hd__mux4_1 _2157_ (.A0(\tms1x00.RAM[84][0] ),
    .A1(\tms1x00.RAM[85][0] ),
    .A2(\tms1x00.RAM[86][0] ),
    .A3(\tms1x00.RAM[87][0] ),
    .S0(_0687_),
    .S1(_0688_),
    .X(_0689_));
 sky130_fd_sc_hd__clkinv_2 _2158_ (.A(_0003_),
    .Y(_0690_));
 sky130_fd_sc_hd__clkbuf_4 _2159_ (.A(_0690_),
    .X(_0691_));
 sky130_fd_sc_hd__o21ai_1 _2160_ (.A1(_0686_),
    .A2(_0689_),
    .B1(_0691_),
    .Y(_0692_));
 sky130_fd_sc_hd__clkbuf_4 _2161_ (.A(_0004_),
    .X(_0693_));
 sky130_fd_sc_hd__o221a_1 _2162_ (.A1(_0670_),
    .A2(_0677_),
    .B1(_0684_),
    .B2(_0692_),
    .C1(_0693_),
    .X(_0694_));
 sky130_fd_sc_hd__buf_2 _2163_ (.A(_0004_),
    .X(_0695_));
 sky130_fd_sc_hd__buf_4 _2164_ (.A(_0001_),
    .X(_0696_));
 sky130_fd_sc_hd__buf_4 _2165_ (.A(_0696_),
    .X(_0697_));
 sky130_fd_sc_hd__buf_6 _2166_ (.A(_0665_),
    .X(_0698_));
 sky130_fd_sc_hd__mux2_1 _2167_ (.A0(\tms1x00.RAM[76][0] ),
    .A1(\tms1x00.RAM[77][0] ),
    .S(_0698_),
    .X(_0699_));
 sky130_fd_sc_hd__and2b_1 _2168_ (.A_N(_0697_),
    .B(_0699_),
    .X(_0700_));
 sky130_fd_sc_hd__buf_6 _2169_ (.A(_0001_),
    .X(_0701_));
 sky130_fd_sc_hd__clkbuf_4 _2170_ (.A(_0701_),
    .X(_0702_));
 sky130_fd_sc_hd__buf_6 _2171_ (.A(_0665_),
    .X(_0703_));
 sky130_fd_sc_hd__mux2_1 _2172_ (.A0(\tms1x00.RAM[78][0] ),
    .A1(\tms1x00.RAM[79][0] ),
    .S(_0703_),
    .X(_0704_));
 sky130_fd_sc_hd__clkbuf_4 _2173_ (.A(_0685_),
    .X(_0705_));
 sky130_fd_sc_hd__a21o_1 _2174_ (.A1(_0702_),
    .A2(_0704_),
    .B1(_0705_),
    .X(_0706_));
 sky130_fd_sc_hd__mux4_1 _2175_ (.A0(\tms1x00.RAM[72][0] ),
    .A1(\tms1x00.RAM[73][0] ),
    .A2(\tms1x00.RAM[74][0] ),
    .A3(\tms1x00.RAM[75][0] ),
    .S0(_0687_),
    .S1(_0688_),
    .X(_0707_));
 sky130_fd_sc_hd__clkbuf_4 _2176_ (.A(_0671_),
    .X(_0708_));
 sky130_fd_sc_hd__clkbuf_4 _2177_ (.A(_0003_),
    .X(_0709_));
 sky130_fd_sc_hd__o221a_1 _2178_ (.A1(_0700_),
    .A2(_0706_),
    .B1(_0707_),
    .B2(_0708_),
    .C1(_0709_),
    .X(_0710_));
 sky130_fd_sc_hd__mux2_1 _2179_ (.A0(\tms1x00.RAM[68][0] ),
    .A1(\tms1x00.RAM[69][0] ),
    .S(_0666_),
    .X(_0711_));
 sky130_fd_sc_hd__and2b_1 _2180_ (.A_N(_0702_),
    .B(_0711_),
    .X(_0712_));
 sky130_fd_sc_hd__buf_4 _2181_ (.A(_0665_),
    .X(_0713_));
 sky130_fd_sc_hd__mux2_1 _2182_ (.A0(\tms1x00.RAM[70][0] ),
    .A1(\tms1x00.RAM[71][0] ),
    .S(_0713_),
    .X(_0714_));
 sky130_fd_sc_hd__clkbuf_4 _2183_ (.A(_0685_),
    .X(_0715_));
 sky130_fd_sc_hd__a21o_1 _2184_ (.A1(_0664_),
    .A2(_0714_),
    .B1(_0715_),
    .X(_0716_));
 sky130_fd_sc_hd__buf_8 _2185_ (.A(_0000_),
    .X(_0717_));
 sky130_fd_sc_hd__buf_6 _2186_ (.A(_0717_),
    .X(_0718_));
 sky130_fd_sc_hd__mux4_2 _2187_ (.A0(\tms1x00.RAM[64][0] ),
    .A1(\tms1x00.RAM[65][0] ),
    .A2(\tms1x00.RAM[66][0] ),
    .A3(\tms1x00.RAM[67][0] ),
    .S0(_0718_),
    .S1(_0682_),
    .X(_0719_));
 sky130_fd_sc_hd__clkbuf_4 _2188_ (.A(_0002_),
    .X(_0720_));
 sky130_fd_sc_hd__clkbuf_4 _2189_ (.A(_0720_),
    .X(_0721_));
 sky130_fd_sc_hd__buf_2 _2190_ (.A(_0690_),
    .X(_0722_));
 sky130_fd_sc_hd__clkbuf_4 _2191_ (.A(_0722_),
    .X(_0723_));
 sky130_fd_sc_hd__o221a_1 _2192_ (.A1(_0712_),
    .A2(_0716_),
    .B1(_0719_),
    .B2(_0721_),
    .C1(_0723_),
    .X(_0724_));
 sky130_fd_sc_hd__nor3_1 _2193_ (.A(_0695_),
    .B(_0710_),
    .C(_0724_),
    .Y(_0725_));
 sky130_fd_sc_hd__mux2_1 _2194_ (.A0(\tms1x00.RAM[118][0] ),
    .A1(\tms1x00.RAM[119][0] ),
    .S(_0713_),
    .X(_0726_));
 sky130_fd_sc_hd__nand2_1 _2195_ (.A(_0660_),
    .B(_0726_),
    .Y(_0727_));
 sky130_fd_sc_hd__mux2_1 _2196_ (.A0(\tms1x00.RAM[116][0] ),
    .A1(\tms1x00.RAM[117][0] ),
    .S(_0679_),
    .X(_0728_));
 sky130_fd_sc_hd__or2b_1 _2197_ (.A(_0674_),
    .B_N(_0728_),
    .X(_0729_));
 sky130_fd_sc_hd__buf_6 _2198_ (.A(_0001_),
    .X(_0730_));
 sky130_fd_sc_hd__mux4_1 _2199_ (.A0(\tms1x00.RAM[112][0] ),
    .A1(\tms1x00.RAM[113][0] ),
    .A2(\tms1x00.RAM[114][0] ),
    .A3(\tms1x00.RAM[115][0] ),
    .S0(_0679_),
    .S1(_0730_),
    .X(_0731_));
 sky130_fd_sc_hd__o21ai_1 _2200_ (.A1(_0671_),
    .A2(_0731_),
    .B1(_0722_),
    .Y(_0732_));
 sky130_fd_sc_hd__a31o_1 _2201_ (.A1(_0672_),
    .A2(_0727_),
    .A3(_0729_),
    .B1(_0732_),
    .X(_0733_));
 sky130_fd_sc_hd__buf_4 _2202_ (.A(_0705_),
    .X(_0734_));
 sky130_fd_sc_hd__mux4_1 _2203_ (.A0(\tms1x00.RAM[124][0] ),
    .A1(\tms1x00.RAM[125][0] ),
    .A2(\tms1x00.RAM[126][0] ),
    .A3(\tms1x00.RAM[127][0] ),
    .S0(_0718_),
    .S1(_0682_),
    .X(_0735_));
 sky130_fd_sc_hd__buf_4 _2204_ (.A(_0002_),
    .X(_0736_));
 sky130_fd_sc_hd__buf_6 _2205_ (.A(_0000_),
    .X(_0737_));
 sky130_fd_sc_hd__buf_4 _2206_ (.A(_0001_),
    .X(_0738_));
 sky130_fd_sc_hd__mux4_1 _2207_ (.A0(\tms1x00.RAM[120][0] ),
    .A1(\tms1x00.RAM[121][0] ),
    .A2(\tms1x00.RAM[122][0] ),
    .A3(\tms1x00.RAM[123][0] ),
    .S0(_0737_),
    .S1(_0738_),
    .X(_0739_));
 sky130_fd_sc_hd__buf_2 _2208_ (.A(_0003_),
    .X(_0740_));
 sky130_fd_sc_hd__o21a_1 _2209_ (.A1(_0736_),
    .A2(_0739_),
    .B1(_0740_),
    .X(_0741_));
 sky130_fd_sc_hd__o21ai_1 _2210_ (.A1(_0734_),
    .A2(_0735_),
    .B1(_0741_),
    .Y(_0742_));
 sky130_fd_sc_hd__clkinv_2 _2211_ (.A(_0005_),
    .Y(_0743_));
 sky130_fd_sc_hd__buf_6 _2212_ (.A(_0000_),
    .X(_0744_));
 sky130_fd_sc_hd__mux4_1 _2213_ (.A0(\tms1x00.RAM[108][0] ),
    .A1(\tms1x00.RAM[109][0] ),
    .A2(\tms1x00.RAM[110][0] ),
    .A3(\tms1x00.RAM[111][0] ),
    .S0(_0744_),
    .S1(_0681_),
    .X(_0745_));
 sky130_fd_sc_hd__nor2_1 _2214_ (.A(_0715_),
    .B(_0745_),
    .Y(_0746_));
 sky130_fd_sc_hd__mux4_2 _2215_ (.A0(\tms1x00.RAM[104][0] ),
    .A1(\tms1x00.RAM[105][0] ),
    .A2(\tms1x00.RAM[106][0] ),
    .A3(\tms1x00.RAM[107][0] ),
    .S0(_0661_),
    .S1(_0658_),
    .X(_0747_));
 sky130_fd_sc_hd__o21ai_1 _2216_ (.A1(_0671_),
    .A2(_0747_),
    .B1(_0740_),
    .Y(_0748_));
 sky130_fd_sc_hd__mux4_1 _2217_ (.A0(\tms1x00.RAM[96][0] ),
    .A1(\tms1x00.RAM[97][0] ),
    .A2(\tms1x00.RAM[98][0] ),
    .A3(\tms1x00.RAM[99][0] ),
    .S0(_0737_),
    .S1(_0696_),
    .X(_0749_));
 sky130_fd_sc_hd__nor2_1 _2218_ (.A(_0736_),
    .B(_0749_),
    .Y(_0750_));
 sky130_fd_sc_hd__clkbuf_4 _2219_ (.A(_0685_),
    .X(_0751_));
 sky130_fd_sc_hd__mux4_1 _2220_ (.A0(\tms1x00.RAM[100][0] ),
    .A1(\tms1x00.RAM[101][0] ),
    .A2(\tms1x00.RAM[102][0] ),
    .A3(\tms1x00.RAM[103][0] ),
    .S0(_0679_),
    .S1(_0730_),
    .X(_0752_));
 sky130_fd_sc_hd__o21ai_1 _2221_ (.A1(_0751_),
    .A2(_0752_),
    .B1(_0722_),
    .Y(_0753_));
 sky130_fd_sc_hd__clkinv_2 _2222_ (.A(_0004_),
    .Y(_0754_));
 sky130_fd_sc_hd__o221a_1 _2223_ (.A1(_0746_),
    .A2(_0748_),
    .B1(_0750_),
    .B2(_0753_),
    .C1(_0754_),
    .X(_0755_));
 sky130_fd_sc_hd__a311o_1 _2224_ (.A1(_0693_),
    .A2(_0733_),
    .A3(_0742_),
    .B1(_0743_),
    .C1(_0755_),
    .X(_0756_));
 sky130_fd_sc_hd__o311a_2 _2225_ (.A1(_0657_),
    .A2(_0694_),
    .A3(_0725_),
    .B1(_0756_),
    .C1(_0006_),
    .X(_0757_));
 sky130_fd_sc_hd__buf_4 _2226_ (.A(_0659_),
    .X(_0758_));
 sky130_fd_sc_hd__buf_6 _2227_ (.A(_0000_),
    .X(_0759_));
 sky130_fd_sc_hd__buf_6 _2228_ (.A(_0759_),
    .X(_0760_));
 sky130_fd_sc_hd__mux2_1 _2229_ (.A0(\tms1x00.RAM[6][0] ),
    .A1(\tms1x00.RAM[7][0] ),
    .S(_0760_),
    .X(_0761_));
 sky130_fd_sc_hd__mux2_1 _2230_ (.A0(\tms1x00.RAM[4][0] ),
    .A1(\tms1x00.RAM[5][0] ),
    .S(_0698_),
    .X(_0762_));
 sky130_fd_sc_hd__and2b_1 _2231_ (.A_N(_0697_),
    .B(_0762_),
    .X(_0763_));
 sky130_fd_sc_hd__a211o_1 _2232_ (.A1(_0758_),
    .A2(_0761_),
    .B1(_0763_),
    .C1(_0734_),
    .X(_0764_));
 sky130_fd_sc_hd__mux4_1 _2233_ (.A0(\tms1x00.RAM[0][0] ),
    .A1(\tms1x00.RAM[1][0] ),
    .A2(\tms1x00.RAM[2][0] ),
    .A3(\tms1x00.RAM[3][0] ),
    .S0(_0687_),
    .S1(_0688_),
    .X(_0765_));
 sky130_fd_sc_hd__or2_1 _2234_ (.A(_0708_),
    .B(_0765_),
    .X(_0766_));
 sky130_fd_sc_hd__buf_4 _2235_ (.A(_0658_),
    .X(_0767_));
 sky130_fd_sc_hd__mux2_1 _2236_ (.A0(\tms1x00.RAM[12][0] ),
    .A1(\tms1x00.RAM[13][0] ),
    .S(_0703_),
    .X(_0768_));
 sky130_fd_sc_hd__and2b_1 _2237_ (.A_N(_0767_),
    .B(_0768_),
    .X(_0769_));
 sky130_fd_sc_hd__mux2_1 _2238_ (.A0(\tms1x00.RAM[14][0] ),
    .A1(\tms1x00.RAM[15][0] ),
    .S(_0713_),
    .X(_0770_));
 sky130_fd_sc_hd__a21o_1 _2239_ (.A1(_0664_),
    .A2(_0770_),
    .B1(_0751_),
    .X(_0771_));
 sky130_fd_sc_hd__mux4_1 _2240_ (.A0(\tms1x00.RAM[8][0] ),
    .A1(\tms1x00.RAM[9][0] ),
    .A2(\tms1x00.RAM[10][0] ),
    .A3(\tms1x00.RAM[11][0] ),
    .S0(_0680_),
    .S1(_0682_),
    .X(_0772_));
 sky130_fd_sc_hd__o221a_1 _2241_ (.A1(_0769_),
    .A2(_0771_),
    .B1(_0772_),
    .B2(_0721_),
    .C1(_0709_),
    .X(_0773_));
 sky130_fd_sc_hd__a311oi_1 _2242_ (.A1(_0723_),
    .A2(_0764_),
    .A3(_0766_),
    .B1(_0695_),
    .C1(_0773_),
    .Y(_0774_));
 sky130_fd_sc_hd__buf_4 _2243_ (.A(_0730_),
    .X(_0775_));
 sky130_fd_sc_hd__mux2_1 _2244_ (.A0(\tms1x00.RAM[28][0] ),
    .A1(\tms1x00.RAM[29][0] ),
    .S(_0759_),
    .X(_0776_));
 sky130_fd_sc_hd__or2b_1 _2245_ (.A(_0775_),
    .B_N(_0776_),
    .X(_0777_));
 sky130_fd_sc_hd__mux2_1 _2246_ (.A0(\tms1x00.RAM[30][0] ),
    .A1(\tms1x00.RAM[31][0] ),
    .S(_0673_),
    .X(_0778_));
 sky130_fd_sc_hd__nand2_1 _2247_ (.A(_0758_),
    .B(_0778_),
    .Y(_0779_));
 sky130_fd_sc_hd__mux4_1 _2248_ (.A0(\tms1x00.RAM[24][0] ),
    .A1(\tms1x00.RAM[25][0] ),
    .A2(\tms1x00.RAM[26][0] ),
    .A3(\tms1x00.RAM[27][0] ),
    .S0(_0759_),
    .S1(_0738_),
    .X(_0780_));
 sky130_fd_sc_hd__o21ai_2 _2249_ (.A1(_0736_),
    .A2(_0780_),
    .B1(_0676_),
    .Y(_0781_));
 sky130_fd_sc_hd__a31o_1 _2250_ (.A1(_0708_),
    .A2(_0777_),
    .A3(_0779_),
    .B1(_0781_),
    .X(_0782_));
 sky130_fd_sc_hd__mux4_1 _2251_ (.A0(\tms1x00.RAM[16][0] ),
    .A1(\tms1x00.RAM[17][0] ),
    .A2(\tms1x00.RAM[18][0] ),
    .A3(\tms1x00.RAM[19][0] ),
    .S0(_0760_),
    .S1(_0702_),
    .X(_0783_));
 sky130_fd_sc_hd__mux4_1 _2252_ (.A0(\tms1x00.RAM[20][0] ),
    .A1(\tms1x00.RAM[21][0] ),
    .A2(\tms1x00.RAM[22][0] ),
    .A3(\tms1x00.RAM[23][0] ),
    .S0(_0703_),
    .S1(_0659_),
    .X(_0784_));
 sky130_fd_sc_hd__o21a_1 _2253_ (.A1(_0686_),
    .A2(_0784_),
    .B1(_0691_),
    .X(_0785_));
 sky130_fd_sc_hd__o21ai_1 _2254_ (.A1(_0721_),
    .A2(_0783_),
    .B1(_0785_),
    .Y(_0786_));
 sky130_fd_sc_hd__a31o_1 _2255_ (.A1(_0695_),
    .A2(_0782_),
    .A3(_0786_),
    .B1(_0657_),
    .X(_0787_));
 sky130_fd_sc_hd__inv_2 _2256_ (.A(_0006_),
    .Y(_0788_));
 sky130_fd_sc_hd__mux2_1 _2257_ (.A0(\tms1x00.RAM[54][0] ),
    .A1(\tms1x00.RAM[55][0] ),
    .S(_0673_),
    .X(_0789_));
 sky130_fd_sc_hd__nand2_1 _2258_ (.A(_0758_),
    .B(_0789_),
    .Y(_0790_));
 sky130_fd_sc_hd__mux2_1 _2259_ (.A0(\tms1x00.RAM[52][0] ),
    .A1(\tms1x00.RAM[53][0] ),
    .S(_0759_),
    .X(_0791_));
 sky130_fd_sc_hd__or2b_1 _2260_ (.A(_0775_),
    .B_N(_0791_),
    .X(_0792_));
 sky130_fd_sc_hd__mux4_1 _2261_ (.A0(\tms1x00.RAM[48][0] ),
    .A1(\tms1x00.RAM[49][0] ),
    .A2(\tms1x00.RAM[50][0] ),
    .A3(\tms1x00.RAM[51][0] ),
    .S0(_0737_),
    .S1(_0738_),
    .X(_0793_));
 sky130_fd_sc_hd__o21ai_1 _2262_ (.A1(_0736_),
    .A2(_0793_),
    .B1(_0691_),
    .Y(_0794_));
 sky130_fd_sc_hd__a31o_1 _2263_ (.A1(_0708_),
    .A2(_0790_),
    .A3(_0792_),
    .B1(_0794_),
    .X(_0795_));
 sky130_fd_sc_hd__mux4_2 _2264_ (.A0(\tms1x00.RAM[60][0] ),
    .A1(\tms1x00.RAM[61][0] ),
    .A2(\tms1x00.RAM[62][0] ),
    .A3(\tms1x00.RAM[63][0] ),
    .S0(_0760_),
    .S1(_0767_),
    .X(_0796_));
 sky130_fd_sc_hd__buf_6 _2265_ (.A(_0665_),
    .X(_0797_));
 sky130_fd_sc_hd__mux4_1 _2266_ (.A0(\tms1x00.RAM[56][0] ),
    .A1(\tms1x00.RAM[57][0] ),
    .A2(\tms1x00.RAM[58][0] ),
    .A3(\tms1x00.RAM[59][0] ),
    .S0(_0797_),
    .S1(_0701_),
    .X(_0798_));
 sky130_fd_sc_hd__o21a_1 _2267_ (.A1(_0669_),
    .A2(_0798_),
    .B1(_0676_),
    .X(_0799_));
 sky130_fd_sc_hd__o21ai_1 _2268_ (.A1(_0734_),
    .A2(_0796_),
    .B1(_0799_),
    .Y(_0800_));
 sky130_fd_sc_hd__mux4_1 _2269_ (.A0(\tms1x00.RAM[44][0] ),
    .A1(\tms1x00.RAM[45][0] ),
    .A2(\tms1x00.RAM[46][0] ),
    .A3(\tms1x00.RAM[47][0] ),
    .S0(_0698_),
    .S1(_0701_),
    .X(_0801_));
 sky130_fd_sc_hd__nor2_1 _2270_ (.A(_0686_),
    .B(_0801_),
    .Y(_0802_));
 sky130_fd_sc_hd__mux4_1 _2271_ (.A0(\tms1x00.RAM[40][0] ),
    .A1(\tms1x00.RAM[41][0] ),
    .A2(\tms1x00.RAM[42][0] ),
    .A3(\tms1x00.RAM[43][0] ),
    .S0(_0717_),
    .S1(_0681_),
    .X(_0803_));
 sky130_fd_sc_hd__o21ai_1 _2272_ (.A1(_0720_),
    .A2(_0803_),
    .B1(_0740_),
    .Y(_0804_));
 sky130_fd_sc_hd__mux4_1 _2273_ (.A0(\tms1x00.RAM[32][0] ),
    .A1(\tms1x00.RAM[33][0] ),
    .A2(\tms1x00.RAM[34][0] ),
    .A3(\tms1x00.RAM[35][0] ),
    .S0(_0797_),
    .S1(_0701_),
    .X(_0805_));
 sky130_fd_sc_hd__nor2_1 _2274_ (.A(_0669_),
    .B(_0805_),
    .Y(_0806_));
 sky130_fd_sc_hd__mux4_1 _2275_ (.A0(\tms1x00.RAM[36][0] ),
    .A1(\tms1x00.RAM[37][0] ),
    .A2(\tms1x00.RAM[38][0] ),
    .A3(\tms1x00.RAM[39][0] ),
    .S0(_0737_),
    .S1(_0696_),
    .X(_0807_));
 sky130_fd_sc_hd__o21ai_1 _2276_ (.A1(_0715_),
    .A2(_0807_),
    .B1(_0691_),
    .Y(_0808_));
 sky130_fd_sc_hd__o221a_1 _2277_ (.A1(_0802_),
    .A2(_0804_),
    .B1(_0806_),
    .B2(_0808_),
    .C1(_0754_),
    .X(_0809_));
 sky130_fd_sc_hd__a311o_1 _2278_ (.A1(_0693_),
    .A2(_0795_),
    .A3(_0800_),
    .B1(_0743_),
    .C1(_0809_),
    .X(_0810_));
 sky130_fd_sc_hd__o211a_1 _2279_ (.A1(_0774_),
    .A2(_0787_),
    .B1(_0788_),
    .C1(_0810_),
    .X(_0811_));
 sky130_fd_sc_hd__o22ai_1 _2280_ (.A1(\tms1x00.ins_in[7] ),
    .A2(_0637_),
    .B1(_0757_),
    .B2(_0811_),
    .Y(_0812_));
 sky130_fd_sc_hd__nor2_1 _2281_ (.A(\tms1x00.ins_in[1] ),
    .B(\tms1x00.ins_in[0] ),
    .Y(_0813_));
 sky130_fd_sc_hd__and3_1 _2282_ (.A(\tms1x00.ins_in[3] ),
    .B(\tms1x00.ins_in[2] ),
    .C(_0813_),
    .X(_0814_));
 sky130_fd_sc_hd__or4b_1 _2283_ (.A(\tms1x00.ins_in[4] ),
    .B(net16),
    .C(_0641_),
    .D_N(_0814_),
    .X(_0815_));
 sky130_fd_sc_hd__nor2_1 _2284_ (.A(\tms1x00.ins_in[5] ),
    .B(_0815_),
    .Y(_0816_));
 sky130_fd_sc_hd__or3_1 _2285_ (.A(\tms1x00.ins_in[7] ),
    .B(\tms1x00.ins_in[6] ),
    .C(_0816_),
    .X(_0817_));
 sky130_fd_sc_hd__nor3_2 _2286_ (.A(\tms1x00.ins_in[1] ),
    .B(\tms1x00.ins_in[0] ),
    .C(_0656_),
    .Y(_0818_));
 sky130_fd_sc_hd__a32o_1 _2287_ (.A1(_0656_),
    .A2(_0812_),
    .A3(_0817_),
    .B1(_0818_),
    .B2(\tms1x00.A[0] ),
    .X(_0819_));
 sky130_fd_sc_hd__buf_4 _2288_ (.A(_0819_),
    .X(_0820_));
 sky130_fd_sc_hd__buf_4 _2289_ (.A(_0820_),
    .X(_0821_));
 sky130_fd_sc_hd__nand3b_4 _2290_ (.A_N(\tms1x00.ram_addr_buff[4] ),
    .B(\tms1x00.ram_addr_buff[5] ),
    .C(\tms1x00.ram_addr_buff[6] ),
    .Y(_0822_));
 sky130_fd_sc_hd__buf_4 _2291_ (.A(_0822_),
    .X(_0823_));
 sky130_fd_sc_hd__nand2_1 _2292_ (.A(\tms1x00.ram_addr_buff[0] ),
    .B(\tms1x00.ram_addr_buff[1] ),
    .Y(_0824_));
 sky130_fd_sc_hd__and2_2 _2293_ (.A(_0815_),
    .B(_0656_),
    .X(_0825_));
 sky130_fd_sc_hd__or3_1 _2294_ (.A(\tms1x00.ram_addr_buff[2] ),
    .B(\tms1x00.ram_addr_buff[3] ),
    .C(_0825_),
    .X(_0826_));
 sky130_fd_sc_hd__or2_4 _2295_ (.A(_0824_),
    .B(_0826_),
    .X(_0827_));
 sky130_fd_sc_hd__or2_2 _2296_ (.A(_0823_),
    .B(_0827_),
    .X(_0828_));
 sky130_fd_sc_hd__mux2_1 _2297_ (.A0(_0821_),
    .A1(\tms1x00.RAM[99][0] ),
    .S(_0828_),
    .X(_0829_));
 sky130_fd_sc_hd__clkbuf_1 _2298_ (.A(_0829_),
    .X(_0015_));
 sky130_fd_sc_hd__mux2_1 _2299_ (.A0(\tms1x00.RAM[92][1] ),
    .A1(\tms1x00.RAM[93][1] ),
    .S(_0665_),
    .X(_0830_));
 sky130_fd_sc_hd__inv_2 _2300_ (.A(_0830_),
    .Y(_0831_));
 sky130_fd_sc_hd__mux2_1 _2301_ (.A0(\tms1x00.RAM[94][1] ),
    .A1(\tms1x00.RAM[95][1] ),
    .S(_0703_),
    .X(_0832_));
 sky130_fd_sc_hd__nand2_1 _2302_ (.A(_0664_),
    .B(_0832_),
    .Y(_0833_));
 sky130_fd_sc_hd__o211a_1 _2303_ (.A1(_0660_),
    .A2(_0831_),
    .B1(_0833_),
    .C1(_0669_),
    .X(_0834_));
 sky130_fd_sc_hd__mux4_1 _2304_ (.A0(\tms1x00.RAM[88][1] ),
    .A1(\tms1x00.RAM[89][1] ),
    .A2(\tms1x00.RAM[90][1] ),
    .A3(\tms1x00.RAM[91][1] ),
    .S0(_0673_),
    .S1(_0674_),
    .X(_0835_));
 sky130_fd_sc_hd__o21ai_1 _2305_ (.A1(_0672_),
    .A2(_0835_),
    .B1(_0676_),
    .Y(_0836_));
 sky130_fd_sc_hd__mux4_2 _2306_ (.A0(\tms1x00.RAM[80][1] ),
    .A1(\tms1x00.RAM[81][1] ),
    .A2(\tms1x00.RAM[82][1] ),
    .A3(\tms1x00.RAM[83][1] ),
    .S0(_0680_),
    .S1(_0775_),
    .X(_0837_));
 sky130_fd_sc_hd__nor2_1 _2307_ (.A(_0678_),
    .B(_0837_),
    .Y(_0838_));
 sky130_fd_sc_hd__mux4_1 _2308_ (.A0(\tms1x00.RAM[84][1] ),
    .A1(\tms1x00.RAM[85][1] ),
    .A2(\tms1x00.RAM[86][1] ),
    .A3(\tms1x00.RAM[87][1] ),
    .S0(_0687_),
    .S1(_0674_),
    .X(_0839_));
 sky130_fd_sc_hd__o21ai_1 _2309_ (.A1(_0686_),
    .A2(_0839_),
    .B1(_0691_),
    .Y(_0840_));
 sky130_fd_sc_hd__o221a_1 _2310_ (.A1(_0834_),
    .A2(_0836_),
    .B1(_0838_),
    .B2(_0840_),
    .C1(_0004_),
    .X(_0841_));
 sky130_fd_sc_hd__mux2_1 _2311_ (.A0(\tms1x00.RAM[76][1] ),
    .A1(\tms1x00.RAM[77][1] ),
    .S(_0698_),
    .X(_0842_));
 sky130_fd_sc_hd__and2b_1 _2312_ (.A_N(_0697_),
    .B(_0842_),
    .X(_0843_));
 sky130_fd_sc_hd__mux2_1 _2313_ (.A0(\tms1x00.RAM[78][1] ),
    .A1(\tms1x00.RAM[79][1] ),
    .S(_0703_),
    .X(_0844_));
 sky130_fd_sc_hd__a21o_1 _2314_ (.A1(_0702_),
    .A2(_0844_),
    .B1(_0705_),
    .X(_0845_));
 sky130_fd_sc_hd__mux4_1 _2315_ (.A0(\tms1x00.RAM[72][1] ),
    .A1(\tms1x00.RAM[73][1] ),
    .A2(\tms1x00.RAM[74][1] ),
    .A3(\tms1x00.RAM[75][1] ),
    .S0(_0687_),
    .S1(_0688_),
    .X(_0846_));
 sky130_fd_sc_hd__o221a_1 _2316_ (.A1(_0843_),
    .A2(_0845_),
    .B1(_0846_),
    .B2(_0708_),
    .C1(_0709_),
    .X(_0847_));
 sky130_fd_sc_hd__mux2_1 _2317_ (.A0(\tms1x00.RAM[68][1] ),
    .A1(\tms1x00.RAM[69][1] ),
    .S(_0703_),
    .X(_0848_));
 sky130_fd_sc_hd__and2b_1 _2318_ (.A_N(_0767_),
    .B(_0848_),
    .X(_0849_));
 sky130_fd_sc_hd__mux2_1 _2319_ (.A0(\tms1x00.RAM[70][1] ),
    .A1(\tms1x00.RAM[71][1] ),
    .S(_0713_),
    .X(_0850_));
 sky130_fd_sc_hd__a21o_1 _2320_ (.A1(_0664_),
    .A2(_0850_),
    .B1(_0751_),
    .X(_0851_));
 sky130_fd_sc_hd__mux4_1 _2321_ (.A0(\tms1x00.RAM[64][1] ),
    .A1(\tms1x00.RAM[65][1] ),
    .A2(\tms1x00.RAM[66][1] ),
    .A3(\tms1x00.RAM[67][1] ),
    .S0(_0680_),
    .S1(_0775_),
    .X(_0852_));
 sky130_fd_sc_hd__o221a_1 _2322_ (.A1(_0849_),
    .A2(_0851_),
    .B1(_0852_),
    .B2(_0678_),
    .C1(_0723_),
    .X(_0853_));
 sky130_fd_sc_hd__nor3_1 _2323_ (.A(_0695_),
    .B(_0847_),
    .C(_0853_),
    .Y(_0854_));
 sky130_fd_sc_hd__mux2_1 _2324_ (.A0(\tms1x00.RAM[118][1] ),
    .A1(\tms1x00.RAM[119][1] ),
    .S(_0713_),
    .X(_0855_));
 sky130_fd_sc_hd__nand2_1 _2325_ (.A(_0660_),
    .B(_0855_),
    .Y(_0856_));
 sky130_fd_sc_hd__mux2_1 _2326_ (.A0(\tms1x00.RAM[116][1] ),
    .A1(\tms1x00.RAM[117][1] ),
    .S(_0679_),
    .X(_0857_));
 sky130_fd_sc_hd__or2b_1 _2327_ (.A(_0659_),
    .B_N(_0857_),
    .X(_0858_));
 sky130_fd_sc_hd__mux4_1 _2328_ (.A0(\tms1x00.RAM[112][1] ),
    .A1(\tms1x00.RAM[113][1] ),
    .A2(\tms1x00.RAM[114][1] ),
    .A3(\tms1x00.RAM[115][1] ),
    .S0(_0679_),
    .S1(_0730_),
    .X(_0859_));
 sky130_fd_sc_hd__o21ai_1 _2329_ (.A1(_0671_),
    .A2(_0859_),
    .B1(_0722_),
    .Y(_0860_));
 sky130_fd_sc_hd__a31o_1 _2330_ (.A1(_0672_),
    .A2(_0856_),
    .A3(_0858_),
    .B1(_0860_),
    .X(_0861_));
 sky130_fd_sc_hd__mux4_1 _2331_ (.A0(\tms1x00.RAM[124][1] ),
    .A1(\tms1x00.RAM[125][1] ),
    .A2(\tms1x00.RAM[126][1] ),
    .A3(\tms1x00.RAM[127][1] ),
    .S0(_0718_),
    .S1(_0682_),
    .X(_0862_));
 sky130_fd_sc_hd__mux4_1 _2332_ (.A0(\tms1x00.RAM[120][1] ),
    .A1(\tms1x00.RAM[121][1] ),
    .A2(\tms1x00.RAM[122][1] ),
    .A3(\tms1x00.RAM[123][1] ),
    .S0(_0737_),
    .S1(_0738_),
    .X(_0863_));
 sky130_fd_sc_hd__o21a_1 _2333_ (.A1(_0736_),
    .A2(_0863_),
    .B1(_0740_),
    .X(_0864_));
 sky130_fd_sc_hd__o21ai_1 _2334_ (.A1(_0734_),
    .A2(_0862_),
    .B1(_0864_),
    .Y(_0865_));
 sky130_fd_sc_hd__mux4_1 _2335_ (.A0(\tms1x00.RAM[108][1] ),
    .A1(\tms1x00.RAM[109][1] ),
    .A2(\tms1x00.RAM[110][1] ),
    .A3(\tms1x00.RAM[111][1] ),
    .S0(_0744_),
    .S1(_0681_),
    .X(_0866_));
 sky130_fd_sc_hd__nor2_1 _2336_ (.A(_0715_),
    .B(_0866_),
    .Y(_0867_));
 sky130_fd_sc_hd__mux4_2 _2337_ (.A0(\tms1x00.RAM[104][1] ),
    .A1(\tms1x00.RAM[105][1] ),
    .A2(\tms1x00.RAM[106][1] ),
    .A3(\tms1x00.RAM[107][1] ),
    .S0(_0661_),
    .S1(_0658_),
    .X(_0868_));
 sky130_fd_sc_hd__o21ai_1 _2338_ (.A1(_0671_),
    .A2(_0868_),
    .B1(_0740_),
    .Y(_0869_));
 sky130_fd_sc_hd__mux4_1 _2339_ (.A0(\tms1x00.RAM[96][1] ),
    .A1(\tms1x00.RAM[97][1] ),
    .A2(\tms1x00.RAM[98][1] ),
    .A3(\tms1x00.RAM[99][1] ),
    .S0(_0744_),
    .S1(_0696_),
    .X(_0870_));
 sky130_fd_sc_hd__nor2_1 _2340_ (.A(_0720_),
    .B(_0870_),
    .Y(_0871_));
 sky130_fd_sc_hd__mux4_1 _2341_ (.A0(\tms1x00.RAM[100][1] ),
    .A1(\tms1x00.RAM[101][1] ),
    .A2(\tms1x00.RAM[102][1] ),
    .A3(\tms1x00.RAM[103][1] ),
    .S0(_0679_),
    .S1(_0730_),
    .X(_0872_));
 sky130_fd_sc_hd__o21ai_1 _2342_ (.A1(_0705_),
    .A2(_0872_),
    .B1(_0722_),
    .Y(_0873_));
 sky130_fd_sc_hd__o221a_1 _2343_ (.A1(_0867_),
    .A2(_0869_),
    .B1(_0871_),
    .B2(_0873_),
    .C1(_0754_),
    .X(_0874_));
 sky130_fd_sc_hd__a311o_1 _2344_ (.A1(_0693_),
    .A2(_0861_),
    .A3(_0865_),
    .B1(_0743_),
    .C1(_0874_),
    .X(_0875_));
 sky130_fd_sc_hd__o311a_2 _2345_ (.A1(_0657_),
    .A2(_0841_),
    .A3(_0854_),
    .B1(_0875_),
    .C1(_0006_),
    .X(_0876_));
 sky130_fd_sc_hd__mux2_1 _2346_ (.A0(\tms1x00.RAM[6][1] ),
    .A1(\tms1x00.RAM[7][1] ),
    .S(_0760_),
    .X(_0877_));
 sky130_fd_sc_hd__mux2_1 _2347_ (.A0(\tms1x00.RAM[4][1] ),
    .A1(\tms1x00.RAM[5][1] ),
    .S(_0698_),
    .X(_0878_));
 sky130_fd_sc_hd__and2b_1 _2348_ (.A_N(_0697_),
    .B(_0878_),
    .X(_0879_));
 sky130_fd_sc_hd__a211o_1 _2349_ (.A1(_0758_),
    .A2(_0877_),
    .B1(_0879_),
    .C1(_0734_),
    .X(_0880_));
 sky130_fd_sc_hd__mux4_1 _2350_ (.A0(\tms1x00.RAM[0][1] ),
    .A1(\tms1x00.RAM[1][1] ),
    .A2(\tms1x00.RAM[2][1] ),
    .A3(\tms1x00.RAM[3][1] ),
    .S0(_0687_),
    .S1(_0674_),
    .X(_0881_));
 sky130_fd_sc_hd__or2_1 _2351_ (.A(_0708_),
    .B(_0881_),
    .X(_0882_));
 sky130_fd_sc_hd__mux2_1 _2352_ (.A0(\tms1x00.RAM[12][1] ),
    .A1(\tms1x00.RAM[13][1] ),
    .S(_0797_),
    .X(_0883_));
 sky130_fd_sc_hd__and2b_1 _2353_ (.A_N(_0767_),
    .B(_0883_),
    .X(_0884_));
 sky130_fd_sc_hd__mux2_1 _2354_ (.A0(\tms1x00.RAM[14][1] ),
    .A1(\tms1x00.RAM[15][1] ),
    .S(_0713_),
    .X(_0885_));
 sky130_fd_sc_hd__a21o_1 _2355_ (.A1(_0664_),
    .A2(_0885_),
    .B1(_0751_),
    .X(_0886_));
 sky130_fd_sc_hd__mux4_1 _2356_ (.A0(\tms1x00.RAM[8][1] ),
    .A1(\tms1x00.RAM[9][1] ),
    .A2(\tms1x00.RAM[10][1] ),
    .A3(\tms1x00.RAM[11][1] ),
    .S0(_0680_),
    .S1(_0775_),
    .X(_0887_));
 sky130_fd_sc_hd__o221a_1 _2357_ (.A1(_0884_),
    .A2(_0886_),
    .B1(_0887_),
    .B2(_0678_),
    .C1(_0709_),
    .X(_0888_));
 sky130_fd_sc_hd__a311oi_1 _2358_ (.A1(_0723_),
    .A2(_0880_),
    .A3(_0882_),
    .B1(_0695_),
    .C1(_0888_),
    .Y(_0889_));
 sky130_fd_sc_hd__mux2_1 _2359_ (.A0(\tms1x00.RAM[28][1] ),
    .A1(\tms1x00.RAM[29][1] ),
    .S(_0759_),
    .X(_0890_));
 sky130_fd_sc_hd__or2b_1 _2360_ (.A(_0775_),
    .B_N(_0890_),
    .X(_0891_));
 sky130_fd_sc_hd__mux2_1 _2361_ (.A0(\tms1x00.RAM[30][1] ),
    .A1(\tms1x00.RAM[31][1] ),
    .S(_0673_),
    .X(_0892_));
 sky130_fd_sc_hd__nand2_1 _2362_ (.A(_0758_),
    .B(_0892_),
    .Y(_0893_));
 sky130_fd_sc_hd__mux4_1 _2363_ (.A0(\tms1x00.RAM[24][1] ),
    .A1(\tms1x00.RAM[25][1] ),
    .A2(\tms1x00.RAM[26][1] ),
    .A3(\tms1x00.RAM[27][1] ),
    .S0(_0737_),
    .S1(_0738_),
    .X(_0894_));
 sky130_fd_sc_hd__o21ai_1 _2364_ (.A1(_0736_),
    .A2(_0894_),
    .B1(_0676_),
    .Y(_0895_));
 sky130_fd_sc_hd__a31o_1 _2365_ (.A1(_0708_),
    .A2(_0891_),
    .A3(_0893_),
    .B1(_0895_),
    .X(_0896_));
 sky130_fd_sc_hd__mux4_2 _2366_ (.A0(\tms1x00.RAM[16][1] ),
    .A1(\tms1x00.RAM[17][1] ),
    .A2(\tms1x00.RAM[18][1] ),
    .A3(\tms1x00.RAM[19][1] ),
    .S0(_0760_),
    .S1(_0767_),
    .X(_0897_));
 sky130_fd_sc_hd__mux4_1 _2367_ (.A0(\tms1x00.RAM[20][1] ),
    .A1(\tms1x00.RAM[21][1] ),
    .A2(\tms1x00.RAM[22][1] ),
    .A3(\tms1x00.RAM[23][1] ),
    .S0(_0703_),
    .S1(_0701_),
    .X(_0898_));
 sky130_fd_sc_hd__o21a_1 _2368_ (.A1(_0686_),
    .A2(_0898_),
    .B1(_0691_),
    .X(_0899_));
 sky130_fd_sc_hd__o21ai_1 _2369_ (.A1(_0721_),
    .A2(_0897_),
    .B1(_0899_),
    .Y(_0900_));
 sky130_fd_sc_hd__a31o_1 _2370_ (.A1(_0693_),
    .A2(_0896_),
    .A3(_0900_),
    .B1(_0657_),
    .X(_0901_));
 sky130_fd_sc_hd__mux2_1 _2371_ (.A0(\tms1x00.RAM[54][1] ),
    .A1(\tms1x00.RAM[55][1] ),
    .S(_0713_),
    .X(_0902_));
 sky130_fd_sc_hd__nand2_1 _2372_ (.A(_0660_),
    .B(_0902_),
    .Y(_0903_));
 sky130_fd_sc_hd__mux2_1 _2373_ (.A0(\tms1x00.RAM[52][1] ),
    .A1(\tms1x00.RAM[53][1] ),
    .S(_0744_),
    .X(_0904_));
 sky130_fd_sc_hd__or2b_1 _2374_ (.A(_0674_),
    .B_N(_0904_),
    .X(_0905_));
 sky130_fd_sc_hd__mux4_1 _2375_ (.A0(\tms1x00.RAM[48][1] ),
    .A1(\tms1x00.RAM[49][1] ),
    .A2(\tms1x00.RAM[50][1] ),
    .A3(\tms1x00.RAM[51][1] ),
    .S0(_0717_),
    .S1(_0681_),
    .X(_0906_));
 sky130_fd_sc_hd__o21ai_1 _2376_ (.A1(_0720_),
    .A2(_0906_),
    .B1(_0722_),
    .Y(_0907_));
 sky130_fd_sc_hd__a31o_1 _2377_ (.A1(_0672_),
    .A2(_0903_),
    .A3(_0905_),
    .B1(_0907_),
    .X(_0908_));
 sky130_fd_sc_hd__mux4_2 _2378_ (.A0(\tms1x00.RAM[60][1] ),
    .A1(\tms1x00.RAM[61][1] ),
    .A2(\tms1x00.RAM[62][1] ),
    .A3(\tms1x00.RAM[63][1] ),
    .S0(_0718_),
    .S1(_0697_),
    .X(_0909_));
 sky130_fd_sc_hd__mux4_1 _2379_ (.A0(\tms1x00.RAM[56][1] ),
    .A1(\tms1x00.RAM[57][1] ),
    .A2(\tms1x00.RAM[58][1] ),
    .A3(\tms1x00.RAM[59][1] ),
    .S0(_0759_),
    .S1(_0738_),
    .X(_0910_));
 sky130_fd_sc_hd__o21a_1 _2380_ (.A1(_0736_),
    .A2(_0910_),
    .B1(_0740_),
    .X(_0911_));
 sky130_fd_sc_hd__o21ai_1 _2381_ (.A1(_0734_),
    .A2(_0909_),
    .B1(_0911_),
    .Y(_0912_));
 sky130_fd_sc_hd__mux4_1 _2382_ (.A0(\tms1x00.RAM[44][1] ),
    .A1(\tms1x00.RAM[45][1] ),
    .A2(\tms1x00.RAM[46][1] ),
    .A3(\tms1x00.RAM[47][1] ),
    .S0(_0717_),
    .S1(_0681_),
    .X(_0913_));
 sky130_fd_sc_hd__nor2_1 _2383_ (.A(_0751_),
    .B(_0913_),
    .Y(_0914_));
 sky130_fd_sc_hd__mux4_2 _2384_ (.A0(\tms1x00.RAM[40][1] ),
    .A1(\tms1x00.RAM[41][1] ),
    .A2(\tms1x00.RAM[42][1] ),
    .A3(\tms1x00.RAM[43][1] ),
    .S0(_0661_),
    .S1(_0658_),
    .X(_0915_));
 sky130_fd_sc_hd__o21ai_1 _2385_ (.A1(_0671_),
    .A2(_0915_),
    .B1(_0003_),
    .Y(_0916_));
 sky130_fd_sc_hd__mux4_2 _2386_ (.A0(\tms1x00.RAM[32][1] ),
    .A1(\tms1x00.RAM[33][1] ),
    .A2(\tms1x00.RAM[34][1] ),
    .A3(\tms1x00.RAM[35][1] ),
    .S0(_0744_),
    .S1(_0696_),
    .X(_0917_));
 sky130_fd_sc_hd__nor2_1 _2387_ (.A(_0720_),
    .B(_0917_),
    .Y(_0918_));
 sky130_fd_sc_hd__mux4_1 _2388_ (.A0(\tms1x00.RAM[36][1] ),
    .A1(\tms1x00.RAM[37][1] ),
    .A2(\tms1x00.RAM[38][1] ),
    .A3(\tms1x00.RAM[39][1] ),
    .S0(_0679_),
    .S1(_0730_),
    .X(_0919_));
 sky130_fd_sc_hd__o21ai_1 _2389_ (.A1(_0705_),
    .A2(_0919_),
    .B1(_0690_),
    .Y(_0920_));
 sky130_fd_sc_hd__o221a_1 _2390_ (.A1(_0914_),
    .A2(_0916_),
    .B1(_0918_),
    .B2(_0920_),
    .C1(_0754_),
    .X(_0921_));
 sky130_fd_sc_hd__a311o_1 _2391_ (.A1(_0693_),
    .A2(_0908_),
    .A3(_0912_),
    .B1(_0921_),
    .C1(_0743_),
    .X(_0922_));
 sky130_fd_sc_hd__o211a_2 _2392_ (.A1(_0889_),
    .A2(_0901_),
    .B1(_0922_),
    .C1(_0788_),
    .X(_0923_));
 sky130_fd_sc_hd__and2b_1 _2393_ (.A_N(\tms1x00.ins_in[7] ),
    .B(\tms1x00.ins_in[6] ),
    .X(_0924_));
 sky130_fd_sc_hd__o21bai_1 _2394_ (.A1(_0876_),
    .A2(_0923_),
    .B1_N(_0924_),
    .Y(_0925_));
 sky130_fd_sc_hd__clkbuf_4 _2395_ (.A(\tms1x00.ins_in[5] ),
    .X(_0926_));
 sky130_fd_sc_hd__o21ai_1 _2396_ (.A1(_0926_),
    .A2(_0815_),
    .B1(_0924_),
    .Y(_0927_));
 sky130_fd_sc_hd__a32o_1 _2397_ (.A1(_0656_),
    .A2(_0925_),
    .A3(_0927_),
    .B1(_0818_),
    .B2(\tms1x00.A[1] ),
    .X(_0928_));
 sky130_fd_sc_hd__buf_4 _2398_ (.A(_0928_),
    .X(_0929_));
 sky130_fd_sc_hd__buf_4 _2399_ (.A(_0929_),
    .X(_0930_));
 sky130_fd_sc_hd__mux2_1 _2400_ (.A0(_0930_),
    .A1(\tms1x00.RAM[99][1] ),
    .S(_0828_),
    .X(_0931_));
 sky130_fd_sc_hd__clkbuf_1 _2401_ (.A(_0931_),
    .X(_0016_));
 sky130_fd_sc_hd__mux2_1 _2402_ (.A0(\tms1x00.RAM[92][2] ),
    .A1(\tms1x00.RAM[93][2] ),
    .S(_0661_),
    .X(_0932_));
 sky130_fd_sc_hd__inv_2 _2403_ (.A(_0932_),
    .Y(_0933_));
 sky130_fd_sc_hd__mux2_1 _2404_ (.A0(\tms1x00.RAM[94][2] ),
    .A1(\tms1x00.RAM[95][2] ),
    .S(_0666_),
    .X(_0934_));
 sky130_fd_sc_hd__nand2_1 _2405_ (.A(_0664_),
    .B(_0934_),
    .Y(_0935_));
 sky130_fd_sc_hd__o211a_1 _2406_ (.A1(_0660_),
    .A2(_0933_),
    .B1(_0935_),
    .C1(_0669_),
    .X(_0936_));
 sky130_fd_sc_hd__mux4_1 _2407_ (.A0(\tms1x00.RAM[88][2] ),
    .A1(\tms1x00.RAM[89][2] ),
    .A2(\tms1x00.RAM[90][2] ),
    .A3(\tms1x00.RAM[91][2] ),
    .S0(_0673_),
    .S1(_0674_),
    .X(_0937_));
 sky130_fd_sc_hd__o21ai_1 _2408_ (.A1(_0672_),
    .A2(_0937_),
    .B1(_0676_),
    .Y(_0938_));
 sky130_fd_sc_hd__mux4_1 _2409_ (.A0(\tms1x00.RAM[80][2] ),
    .A1(\tms1x00.RAM[81][2] ),
    .A2(\tms1x00.RAM[82][2] ),
    .A3(\tms1x00.RAM[83][2] ),
    .S0(_0680_),
    .S1(_0775_),
    .X(_0939_));
 sky130_fd_sc_hd__nor2_1 _2410_ (.A(_0678_),
    .B(_0939_),
    .Y(_0940_));
 sky130_fd_sc_hd__mux4_1 _2411_ (.A0(\tms1x00.RAM[84][2] ),
    .A1(\tms1x00.RAM[85][2] ),
    .A2(\tms1x00.RAM[86][2] ),
    .A3(\tms1x00.RAM[87][2] ),
    .S0(_0687_),
    .S1(_0674_),
    .X(_0941_));
 sky130_fd_sc_hd__o21ai_1 _2412_ (.A1(_0686_),
    .A2(_0941_),
    .B1(_0691_),
    .Y(_0942_));
 sky130_fd_sc_hd__o221a_1 _2413_ (.A1(_0936_),
    .A2(_0938_),
    .B1(_0940_),
    .B2(_0942_),
    .C1(_0693_),
    .X(_0943_));
 sky130_fd_sc_hd__mux2_1 _2414_ (.A0(\tms1x00.RAM[76][2] ),
    .A1(\tms1x00.RAM[77][2] ),
    .S(_0698_),
    .X(_0944_));
 sky130_fd_sc_hd__and2b_1 _2415_ (.A_N(_0697_),
    .B(_0944_),
    .X(_0945_));
 sky130_fd_sc_hd__mux2_1 _2416_ (.A0(\tms1x00.RAM[78][2] ),
    .A1(\tms1x00.RAM[79][2] ),
    .S(_0703_),
    .X(_0946_));
 sky130_fd_sc_hd__a21o_1 _2417_ (.A1(_0702_),
    .A2(_0946_),
    .B1(_0705_),
    .X(_0947_));
 sky130_fd_sc_hd__mux4_1 _2418_ (.A0(\tms1x00.RAM[72][2] ),
    .A1(\tms1x00.RAM[73][2] ),
    .A2(\tms1x00.RAM[74][2] ),
    .A3(\tms1x00.RAM[75][2] ),
    .S0(_0687_),
    .S1(_0688_),
    .X(_0948_));
 sky130_fd_sc_hd__o221a_1 _2419_ (.A1(_0945_),
    .A2(_0947_),
    .B1(_0948_),
    .B2(_0708_),
    .C1(_0709_),
    .X(_0949_));
 sky130_fd_sc_hd__mux2_1 _2420_ (.A0(\tms1x00.RAM[68][2] ),
    .A1(\tms1x00.RAM[69][2] ),
    .S(_0666_),
    .X(_0950_));
 sky130_fd_sc_hd__and2b_1 _2421_ (.A_N(_0702_),
    .B(_0950_),
    .X(_0951_));
 sky130_fd_sc_hd__mux2_1 _2422_ (.A0(\tms1x00.RAM[70][2] ),
    .A1(\tms1x00.RAM[71][2] ),
    .S(_0713_),
    .X(_0952_));
 sky130_fd_sc_hd__a21o_1 _2423_ (.A1(_0664_),
    .A2(_0952_),
    .B1(_0751_),
    .X(_0953_));
 sky130_fd_sc_hd__mux4_2 _2424_ (.A0(\tms1x00.RAM[64][2] ),
    .A1(\tms1x00.RAM[65][2] ),
    .A2(\tms1x00.RAM[66][2] ),
    .A3(\tms1x00.RAM[67][2] ),
    .S0(_0718_),
    .S1(_0682_),
    .X(_0954_));
 sky130_fd_sc_hd__o221a_1 _2425_ (.A1(_0951_),
    .A2(_0953_),
    .B1(_0954_),
    .B2(_0721_),
    .C1(_0723_),
    .X(_0955_));
 sky130_fd_sc_hd__nor3_1 _2426_ (.A(_0695_),
    .B(_0949_),
    .C(_0955_),
    .Y(_0956_));
 sky130_fd_sc_hd__mux2_1 _2427_ (.A0(\tms1x00.RAM[118][2] ),
    .A1(\tms1x00.RAM[119][2] ),
    .S(_0673_),
    .X(_0957_));
 sky130_fd_sc_hd__nand2_1 _2428_ (.A(_0660_),
    .B(_0957_),
    .Y(_0958_));
 sky130_fd_sc_hd__mux2_1 _2429_ (.A0(\tms1x00.RAM[116][2] ),
    .A1(\tms1x00.RAM[117][2] ),
    .S(_0744_),
    .X(_0959_));
 sky130_fd_sc_hd__or2b_1 _2430_ (.A(_0688_),
    .B_N(_0959_),
    .X(_0960_));
 sky130_fd_sc_hd__mux4_1 _2431_ (.A0(\tms1x00.RAM[112][2] ),
    .A1(\tms1x00.RAM[113][2] ),
    .A2(\tms1x00.RAM[114][2] ),
    .A3(\tms1x00.RAM[115][2] ),
    .S0(_0717_),
    .S1(_0681_),
    .X(_0961_));
 sky130_fd_sc_hd__o21ai_1 _2432_ (.A1(_0720_),
    .A2(_0961_),
    .B1(_0722_),
    .Y(_0962_));
 sky130_fd_sc_hd__a31o_1 _2433_ (.A1(_0672_),
    .A2(_0958_),
    .A3(_0960_),
    .B1(_0962_),
    .X(_0963_));
 sky130_fd_sc_hd__mux4_1 _2434_ (.A0(\tms1x00.RAM[124][2] ),
    .A1(\tms1x00.RAM[125][2] ),
    .A2(\tms1x00.RAM[126][2] ),
    .A3(\tms1x00.RAM[127][2] ),
    .S0(_0718_),
    .S1(_0697_),
    .X(_0964_));
 sky130_fd_sc_hd__mux4_1 _2435_ (.A0(\tms1x00.RAM[120][2] ),
    .A1(\tms1x00.RAM[121][2] ),
    .A2(\tms1x00.RAM[122][2] ),
    .A3(\tms1x00.RAM[123][2] ),
    .S0(_0698_),
    .S1(_0701_),
    .X(_0965_));
 sky130_fd_sc_hd__o21a_1 _2436_ (.A1(_0669_),
    .A2(_0965_),
    .B1(_0740_),
    .X(_0966_));
 sky130_fd_sc_hd__o21ai_1 _2437_ (.A1(_0734_),
    .A2(_0964_),
    .B1(_0966_),
    .Y(_0967_));
 sky130_fd_sc_hd__mux4_1 _2438_ (.A0(\tms1x00.RAM[108][2] ),
    .A1(\tms1x00.RAM[109][2] ),
    .A2(\tms1x00.RAM[110][2] ),
    .A3(\tms1x00.RAM[111][2] ),
    .S0(_0717_),
    .S1(_0681_),
    .X(_0968_));
 sky130_fd_sc_hd__nor2_1 _2439_ (.A(_0715_),
    .B(_0968_),
    .Y(_0969_));
 sky130_fd_sc_hd__mux4_2 _2440_ (.A0(\tms1x00.RAM[104][2] ),
    .A1(\tms1x00.RAM[105][2] ),
    .A2(\tms1x00.RAM[106][2] ),
    .A3(\tms1x00.RAM[107][2] ),
    .S0(_0661_),
    .S1(_0658_),
    .X(_0970_));
 sky130_fd_sc_hd__o21ai_1 _2441_ (.A1(_0671_),
    .A2(_0970_),
    .B1(_0740_),
    .Y(_0971_));
 sky130_fd_sc_hd__mux4_1 _2442_ (.A0(\tms1x00.RAM[96][2] ),
    .A1(\tms1x00.RAM[97][2] ),
    .A2(\tms1x00.RAM[98][2] ),
    .A3(\tms1x00.RAM[99][2] ),
    .S0(_0744_),
    .S1(_0696_),
    .X(_0972_));
 sky130_fd_sc_hd__nor2_1 _2443_ (.A(_0720_),
    .B(_0972_),
    .Y(_0973_));
 sky130_fd_sc_hd__mux4_1 _2444_ (.A0(\tms1x00.RAM[100][2] ),
    .A1(\tms1x00.RAM[101][2] ),
    .A2(\tms1x00.RAM[102][2] ),
    .A3(\tms1x00.RAM[103][2] ),
    .S0(_0679_),
    .S1(_0730_),
    .X(_0974_));
 sky130_fd_sc_hd__o21ai_1 _2445_ (.A1(_0705_),
    .A2(_0974_),
    .B1(_0690_),
    .Y(_0975_));
 sky130_fd_sc_hd__o221a_1 _2446_ (.A1(_0969_),
    .A2(_0971_),
    .B1(_0973_),
    .B2(_0975_),
    .C1(_0754_),
    .X(_0976_));
 sky130_fd_sc_hd__a311o_1 _2447_ (.A1(_0693_),
    .A2(_0963_),
    .A3(_0967_),
    .B1(_0976_),
    .C1(_0743_),
    .X(_0977_));
 sky130_fd_sc_hd__o311a_2 _2448_ (.A1(_0657_),
    .A2(_0943_),
    .A3(_0956_),
    .B1(_0006_),
    .C1(_0977_),
    .X(_0978_));
 sky130_fd_sc_hd__mux2_1 _2449_ (.A0(\tms1x00.RAM[6][2] ),
    .A1(\tms1x00.RAM[7][2] ),
    .S(_0760_),
    .X(_0979_));
 sky130_fd_sc_hd__mux2_1 _2450_ (.A0(\tms1x00.RAM[4][2] ),
    .A1(\tms1x00.RAM[5][2] ),
    .S(_0698_),
    .X(_0980_));
 sky130_fd_sc_hd__and2b_1 _2451_ (.A_N(_0682_),
    .B(_0980_),
    .X(_0981_));
 sky130_fd_sc_hd__a211o_1 _2452_ (.A1(_0758_),
    .A2(_0979_),
    .B1(_0981_),
    .C1(_0686_),
    .X(_0982_));
 sky130_fd_sc_hd__mux4_1 _2453_ (.A0(\tms1x00.RAM[0][2] ),
    .A1(\tms1x00.RAM[1][2] ),
    .A2(\tms1x00.RAM[2][2] ),
    .A3(\tms1x00.RAM[3][2] ),
    .S0(_0687_),
    .S1(_0674_),
    .X(_0983_));
 sky130_fd_sc_hd__or2_1 _2454_ (.A(_0708_),
    .B(_0983_),
    .X(_0984_));
 sky130_fd_sc_hd__mux2_1 _2455_ (.A0(\tms1x00.RAM[12][2] ),
    .A1(\tms1x00.RAM[13][2] ),
    .S(_0797_),
    .X(_0985_));
 sky130_fd_sc_hd__and2b_1 _2456_ (.A_N(_0767_),
    .B(_0985_),
    .X(_0986_));
 sky130_fd_sc_hd__mux2_1 _2457_ (.A0(\tms1x00.RAM[14][2] ),
    .A1(\tms1x00.RAM[15][2] ),
    .S(_0666_),
    .X(_0987_));
 sky130_fd_sc_hd__a21o_1 _2458_ (.A1(_0664_),
    .A2(_0987_),
    .B1(_0751_),
    .X(_0988_));
 sky130_fd_sc_hd__mux4_1 _2459_ (.A0(\tms1x00.RAM[8][2] ),
    .A1(\tms1x00.RAM[9][2] ),
    .A2(\tms1x00.RAM[10][2] ),
    .A3(\tms1x00.RAM[11][2] ),
    .S0(_0680_),
    .S1(_0775_),
    .X(_0989_));
 sky130_fd_sc_hd__o221a_1 _2460_ (.A1(_0986_),
    .A2(_0988_),
    .B1(_0989_),
    .B2(_0678_),
    .C1(_0709_),
    .X(_0990_));
 sky130_fd_sc_hd__a311oi_1 _2461_ (.A1(_0723_),
    .A2(_0982_),
    .A3(_0984_),
    .B1(_0695_),
    .C1(_0990_),
    .Y(_0991_));
 sky130_fd_sc_hd__mux2_1 _2462_ (.A0(\tms1x00.RAM[28][2] ),
    .A1(\tms1x00.RAM[29][2] ),
    .S(_0759_),
    .X(_0992_));
 sky130_fd_sc_hd__or2b_1 _2463_ (.A(_0775_),
    .B_N(_0992_),
    .X(_0993_));
 sky130_fd_sc_hd__mux2_1 _2464_ (.A0(\tms1x00.RAM[30][2] ),
    .A1(\tms1x00.RAM[31][2] ),
    .S(_0673_),
    .X(_0994_));
 sky130_fd_sc_hd__nand2_1 _2465_ (.A(_0758_),
    .B(_0994_),
    .Y(_0995_));
 sky130_fd_sc_hd__mux4_1 _2466_ (.A0(\tms1x00.RAM[24][2] ),
    .A1(\tms1x00.RAM[25][2] ),
    .A2(\tms1x00.RAM[26][2] ),
    .A3(\tms1x00.RAM[27][2] ),
    .S0(_0737_),
    .S1(_0738_),
    .X(_0996_));
 sky130_fd_sc_hd__o21ai_2 _2467_ (.A1(_0736_),
    .A2(_0996_),
    .B1(_0676_),
    .Y(_0997_));
 sky130_fd_sc_hd__a31o_1 _2468_ (.A1(_0672_),
    .A2(_0993_),
    .A3(_0995_),
    .B1(_0997_),
    .X(_0998_));
 sky130_fd_sc_hd__mux4_2 _2469_ (.A0(\tms1x00.RAM[16][2] ),
    .A1(\tms1x00.RAM[17][2] ),
    .A2(\tms1x00.RAM[18][2] ),
    .A3(\tms1x00.RAM[19][2] ),
    .S0(_0718_),
    .S1(_0767_),
    .X(_0999_));
 sky130_fd_sc_hd__mux4_1 _2470_ (.A0(\tms1x00.RAM[20][2] ),
    .A1(\tms1x00.RAM[21][2] ),
    .A2(\tms1x00.RAM[22][2] ),
    .A3(\tms1x00.RAM[23][2] ),
    .S0(_0797_),
    .S1(_0701_),
    .X(_1000_));
 sky130_fd_sc_hd__o21a_1 _2471_ (.A1(_0686_),
    .A2(_1000_),
    .B1(_0691_),
    .X(_1001_));
 sky130_fd_sc_hd__o21ai_1 _2472_ (.A1(_0721_),
    .A2(_0999_),
    .B1(_1001_),
    .Y(_1002_));
 sky130_fd_sc_hd__a31o_1 _2473_ (.A1(_0693_),
    .A2(_0998_),
    .A3(_1002_),
    .B1(_0657_),
    .X(_1003_));
 sky130_fd_sc_hd__mux2_1 _2474_ (.A0(\tms1x00.RAM[54][2] ),
    .A1(\tms1x00.RAM[55][2] ),
    .S(_0673_),
    .X(_1004_));
 sky130_fd_sc_hd__nand2_1 _2475_ (.A(_0660_),
    .B(_1004_),
    .Y(_1005_));
 sky130_fd_sc_hd__mux2_1 _2476_ (.A0(\tms1x00.RAM[52][2] ),
    .A1(\tms1x00.RAM[53][2] ),
    .S(_0737_),
    .X(_1006_));
 sky130_fd_sc_hd__or2b_1 _2477_ (.A(_0688_),
    .B_N(_1006_),
    .X(_1007_));
 sky130_fd_sc_hd__mux4_1 _2478_ (.A0(\tms1x00.RAM[48][2] ),
    .A1(\tms1x00.RAM[49][2] ),
    .A2(\tms1x00.RAM[50][2] ),
    .A3(\tms1x00.RAM[51][2] ),
    .S0(_0744_),
    .S1(_0696_),
    .X(_1008_));
 sky130_fd_sc_hd__o21ai_1 _2479_ (.A1(_0736_),
    .A2(_1008_),
    .B1(_0722_),
    .Y(_1009_));
 sky130_fd_sc_hd__a31o_1 _2480_ (.A1(_0672_),
    .A2(_1005_),
    .A3(_1007_),
    .B1(_1009_),
    .X(_1010_));
 sky130_fd_sc_hd__mux4_2 _2481_ (.A0(\tms1x00.RAM[60][2] ),
    .A1(\tms1x00.RAM[61][2] ),
    .A2(\tms1x00.RAM[62][2] ),
    .A3(\tms1x00.RAM[63][2] ),
    .S0(_0718_),
    .S1(_0767_),
    .X(_1011_));
 sky130_fd_sc_hd__mux4_1 _2482_ (.A0(\tms1x00.RAM[56][2] ),
    .A1(\tms1x00.RAM[57][2] ),
    .A2(\tms1x00.RAM[58][2] ),
    .A3(\tms1x00.RAM[59][2] ),
    .S0(_0797_),
    .S1(_0701_),
    .X(_1012_));
 sky130_fd_sc_hd__o21a_1 _2483_ (.A1(_0669_),
    .A2(_1012_),
    .B1(_0676_),
    .X(_1013_));
 sky130_fd_sc_hd__o21ai_1 _2484_ (.A1(_0734_),
    .A2(_1011_),
    .B1(_1013_),
    .Y(_1014_));
 sky130_fd_sc_hd__mux4_1 _2485_ (.A0(\tms1x00.RAM[44][2] ),
    .A1(\tms1x00.RAM[45][2] ),
    .A2(\tms1x00.RAM[46][2] ),
    .A3(\tms1x00.RAM[47][2] ),
    .S0(_0759_),
    .S1(_0738_),
    .X(_1015_));
 sky130_fd_sc_hd__nor2_1 _2486_ (.A(_0715_),
    .B(_1015_),
    .Y(_1016_));
 sky130_fd_sc_hd__mux4_2 _2487_ (.A0(\tms1x00.RAM[40][2] ),
    .A1(\tms1x00.RAM[41][2] ),
    .A2(\tms1x00.RAM[42][2] ),
    .A3(\tms1x00.RAM[43][2] ),
    .S0(_0717_),
    .S1(_0730_),
    .X(_1017_));
 sky130_fd_sc_hd__o21ai_1 _2488_ (.A1(_0720_),
    .A2(_1017_),
    .B1(_0740_),
    .Y(_1018_));
 sky130_fd_sc_hd__mux4_1 _2489_ (.A0(\tms1x00.RAM[32][2] ),
    .A1(\tms1x00.RAM[33][2] ),
    .A2(\tms1x00.RAM[34][2] ),
    .A3(\tms1x00.RAM[35][2] ),
    .S0(_0797_),
    .S1(_0701_),
    .X(_1019_));
 sky130_fd_sc_hd__nor2_1 _2490_ (.A(_0669_),
    .B(_1019_),
    .Y(_1020_));
 sky130_fd_sc_hd__mux4_1 _2491_ (.A0(\tms1x00.RAM[36][2] ),
    .A1(\tms1x00.RAM[37][2] ),
    .A2(\tms1x00.RAM[38][2] ),
    .A3(\tms1x00.RAM[39][2] ),
    .S0(_0744_),
    .S1(_0696_),
    .X(_1021_));
 sky130_fd_sc_hd__o21ai_1 _2492_ (.A1(_0715_),
    .A2(_1021_),
    .B1(_0722_),
    .Y(_1022_));
 sky130_fd_sc_hd__o221a_1 _2493_ (.A1(_1016_),
    .A2(_1018_),
    .B1(_1020_),
    .B2(_1022_),
    .C1(_0754_),
    .X(_1023_));
 sky130_fd_sc_hd__a311o_1 _2494_ (.A1(_0693_),
    .A2(_1010_),
    .A3(_1014_),
    .B1(_0743_),
    .C1(_1023_),
    .X(_1024_));
 sky130_fd_sc_hd__o211a_1 _2495_ (.A1(_0991_),
    .A2(_1003_),
    .B1(_0788_),
    .C1(_1024_),
    .X(_1025_));
 sky130_fd_sc_hd__o21ai_1 _2496_ (.A1(_0978_),
    .A2(_1025_),
    .B1(_0647_),
    .Y(_1026_));
 sky130_fd_sc_hd__or3b_1 _2497_ (.A(_0637_),
    .B(_0816_),
    .C_N(\tms1x00.ins_in[7] ),
    .X(_1027_));
 sky130_fd_sc_hd__a32o_1 _2498_ (.A1(_0656_),
    .A2(_1026_),
    .A3(_1027_),
    .B1(_0818_),
    .B2(\tms1x00.A[2] ),
    .X(_1028_));
 sky130_fd_sc_hd__buf_4 _2499_ (.A(_1028_),
    .X(_1029_));
 sky130_fd_sc_hd__buf_4 _2500_ (.A(_1029_),
    .X(_1030_));
 sky130_fd_sc_hd__mux2_1 _2501_ (.A0(_1030_),
    .A1(\tms1x00.RAM[99][2] ),
    .S(_0828_),
    .X(_1031_));
 sky130_fd_sc_hd__clkbuf_1 _2502_ (.A(_1031_),
    .X(_0017_));
 sky130_fd_sc_hd__mux2_1 _2503_ (.A0(\tms1x00.RAM[116][3] ),
    .A1(\tms1x00.RAM[117][3] ),
    .S(_0665_),
    .X(_1032_));
 sky130_fd_sc_hd__and2b_1 _2504_ (.A_N(_0659_),
    .B(_1032_),
    .X(_1033_));
 sky130_fd_sc_hd__mux2_1 _2505_ (.A0(\tms1x00.RAM[118][3] ),
    .A1(\tms1x00.RAM[119][3] ),
    .S(_0661_),
    .X(_1034_));
 sky130_fd_sc_hd__a21o_1 _2506_ (.A1(_0659_),
    .A2(_1034_),
    .B1(_0685_),
    .X(_1035_));
 sky130_fd_sc_hd__mux4_1 _2507_ (.A0(\tms1x00.RAM[112][3] ),
    .A1(\tms1x00.RAM[113][3] ),
    .A2(\tms1x00.RAM[114][3] ),
    .A3(\tms1x00.RAM[115][3] ),
    .S0(_0759_),
    .S1(_0738_),
    .X(_1036_));
 sky130_fd_sc_hd__o221a_1 _2508_ (.A1(_1033_),
    .A2(_1035_),
    .B1(_1036_),
    .B2(_0669_),
    .C1(_0691_),
    .X(_1037_));
 sky130_fd_sc_hd__mux4_1 _2509_ (.A0(\tms1x00.RAM[120][3] ),
    .A1(\tms1x00.RAM[121][3] ),
    .A2(\tms1x00.RAM[122][3] ),
    .A3(\tms1x00.RAM[123][3] ),
    .S0(_0703_),
    .S1(_0659_),
    .X(_1038_));
 sky130_fd_sc_hd__mux4_1 _2510_ (.A0(\tms1x00.RAM[124][3] ),
    .A1(\tms1x00.RAM[125][3] ),
    .A2(\tms1x00.RAM[126][3] ),
    .A3(\tms1x00.RAM[127][3] ),
    .S0(_0665_),
    .S1(_0001_),
    .X(_1039_));
 sky130_fd_sc_hd__or2_1 _2511_ (.A(_0685_),
    .B(_1039_),
    .X(_1040_));
 sky130_fd_sc_hd__o211a_1 _2512_ (.A1(_0669_),
    .A2(_1038_),
    .B1(_1040_),
    .C1(_0676_),
    .X(_1041_));
 sky130_fd_sc_hd__o31a_1 _2513_ (.A1(_0754_),
    .A2(_1037_),
    .A3(_1041_),
    .B1(_0657_),
    .X(_1042_));
 sky130_fd_sc_hd__mux4_1 _2514_ (.A0(\tms1x00.RAM[100][3] ),
    .A1(\tms1x00.RAM[101][3] ),
    .A2(\tms1x00.RAM[102][3] ),
    .A3(\tms1x00.RAM[103][3] ),
    .S0(_0698_),
    .S1(_0701_),
    .X(_1043_));
 sky130_fd_sc_hd__or2_1 _2515_ (.A(_0686_),
    .B(_1043_),
    .X(_1044_));
 sky130_fd_sc_hd__mux4_1 _2516_ (.A0(\tms1x00.RAM[96][3] ),
    .A1(\tms1x00.RAM[97][3] ),
    .A2(\tms1x00.RAM[98][3] ),
    .A3(\tms1x00.RAM[99][3] ),
    .S0(_0759_),
    .S1(_0738_),
    .X(_1045_));
 sky130_fd_sc_hd__or2_1 _2517_ (.A(_0736_),
    .B(_1045_),
    .X(_1046_));
 sky130_fd_sc_hd__mux4_2 _2518_ (.A0(\tms1x00.RAM[108][3] ),
    .A1(\tms1x00.RAM[109][3] ),
    .A2(\tms1x00.RAM[110][3] ),
    .A3(\tms1x00.RAM[111][3] ),
    .S0(_0666_),
    .S1(_0659_),
    .X(_1047_));
 sky130_fd_sc_hd__mux4_2 _2519_ (.A0(\tms1x00.RAM[104][3] ),
    .A1(\tms1x00.RAM[105][3] ),
    .A2(\tms1x00.RAM[106][3] ),
    .A3(\tms1x00.RAM[107][3] ),
    .S0(_0665_),
    .S1(_0658_),
    .X(_1048_));
 sky130_fd_sc_hd__or2_1 _2520_ (.A(_0002_),
    .B(_1048_),
    .X(_1049_));
 sky130_fd_sc_hd__o211a_1 _2521_ (.A1(_0686_),
    .A2(_1047_),
    .B1(_1049_),
    .C1(_0676_),
    .X(_1050_));
 sky130_fd_sc_hd__a311o_1 _2522_ (.A1(_0723_),
    .A2(_1044_),
    .A3(_1046_),
    .B1(_0004_),
    .C1(_1050_),
    .X(_1051_));
 sky130_fd_sc_hd__mux2_1 _2523_ (.A0(\tms1x00.RAM[92][3] ),
    .A1(\tms1x00.RAM[93][3] ),
    .S(_0661_),
    .X(_1052_));
 sky130_fd_sc_hd__or2b_1 _2524_ (.A(_0659_),
    .B_N(_1052_),
    .X(_1053_));
 sky130_fd_sc_hd__mux2_1 _2525_ (.A0(\tms1x00.RAM[94][3] ),
    .A1(\tms1x00.RAM[95][3] ),
    .S(_0713_),
    .X(_1054_));
 sky130_fd_sc_hd__nand2_1 _2526_ (.A(_0660_),
    .B(_1054_),
    .Y(_1055_));
 sky130_fd_sc_hd__mux4_1 _2527_ (.A0(\tms1x00.RAM[88][3] ),
    .A1(\tms1x00.RAM[89][3] ),
    .A2(\tms1x00.RAM[90][3] ),
    .A3(\tms1x00.RAM[91][3] ),
    .S0(_0661_),
    .S1(_0658_),
    .X(_1056_));
 sky130_fd_sc_hd__o21ai_1 _2528_ (.A1(_0671_),
    .A2(_1056_),
    .B1(_0003_),
    .Y(_1057_));
 sky130_fd_sc_hd__a31o_1 _2529_ (.A1(_0672_),
    .A2(_1053_),
    .A3(_1055_),
    .B1(_1057_),
    .X(_1058_));
 sky130_fd_sc_hd__mux4_2 _2530_ (.A0(\tms1x00.RAM[80][3] ),
    .A1(\tms1x00.RAM[81][3] ),
    .A2(\tms1x00.RAM[82][3] ),
    .A3(\tms1x00.RAM[83][3] ),
    .S0(_0680_),
    .S1(_0688_),
    .X(_1059_));
 sky130_fd_sc_hd__mux4_1 _2531_ (.A0(\tms1x00.RAM[84][3] ),
    .A1(\tms1x00.RAM[85][3] ),
    .A2(\tms1x00.RAM[86][3] ),
    .A3(\tms1x00.RAM[87][3] ),
    .S0(_0717_),
    .S1(_0681_),
    .X(_1060_));
 sky130_fd_sc_hd__o21a_1 _2532_ (.A1(_0715_),
    .A2(_1060_),
    .B1(_0690_),
    .X(_1061_));
 sky130_fd_sc_hd__o21ai_1 _2533_ (.A1(_0678_),
    .A2(_1059_),
    .B1(_1061_),
    .Y(_1062_));
 sky130_fd_sc_hd__a31o_1 _2534_ (.A1(_0004_),
    .A2(_1058_),
    .A3(_1062_),
    .B1(_0657_),
    .X(_1063_));
 sky130_fd_sc_hd__mux2_1 _2535_ (.A0(\tms1x00.RAM[76][3] ),
    .A1(\tms1x00.RAM[77][3] ),
    .S(_0737_),
    .X(_1064_));
 sky130_fd_sc_hd__and2b_1 _2536_ (.A_N(_0682_),
    .B(_1064_),
    .X(_1065_));
 sky130_fd_sc_hd__mux2_1 _2537_ (.A0(\tms1x00.RAM[78][3] ),
    .A1(\tms1x00.RAM[79][3] ),
    .S(_0698_),
    .X(_1066_));
 sky130_fd_sc_hd__a21o_1 _2538_ (.A1(_0697_),
    .A2(_1066_),
    .B1(_0705_),
    .X(_1067_));
 sky130_fd_sc_hd__mux4_1 _2539_ (.A0(\tms1x00.RAM[72][3] ),
    .A1(\tms1x00.RAM[73][3] ),
    .A2(\tms1x00.RAM[74][3] ),
    .A3(\tms1x00.RAM[75][3] ),
    .S0(_0673_),
    .S1(_0674_),
    .X(_1068_));
 sky130_fd_sc_hd__o221a_1 _2540_ (.A1(_1065_),
    .A2(_1067_),
    .B1(_1068_),
    .B2(_0708_),
    .C1(_0709_),
    .X(_1069_));
 sky130_fd_sc_hd__mux2_1 _2541_ (.A0(\tms1x00.RAM[68][3] ),
    .A1(\tms1x00.RAM[69][3] ),
    .S(_0797_),
    .X(_1070_));
 sky130_fd_sc_hd__and2b_1 _2542_ (.A_N(_0697_),
    .B(_1070_),
    .X(_1071_));
 sky130_fd_sc_hd__mux2_1 _2543_ (.A0(\tms1x00.RAM[70][3] ),
    .A1(\tms1x00.RAM[71][3] ),
    .S(_0666_),
    .X(_1072_));
 sky130_fd_sc_hd__a21o_1 _2544_ (.A1(_0702_),
    .A2(_1072_),
    .B1(_0705_),
    .X(_1073_));
 sky130_fd_sc_hd__mux4_1 _2545_ (.A0(\tms1x00.RAM[64][3] ),
    .A1(\tms1x00.RAM[65][3] ),
    .A2(\tms1x00.RAM[66][3] ),
    .A3(\tms1x00.RAM[67][3] ),
    .S0(_0680_),
    .S1(_0688_),
    .X(_1074_));
 sky130_fd_sc_hd__o221a_1 _2546_ (.A1(_1071_),
    .A2(_1073_),
    .B1(_1074_),
    .B2(_0678_),
    .C1(_0723_),
    .X(_1075_));
 sky130_fd_sc_hd__nor3_1 _2547_ (.A(_0695_),
    .B(_1069_),
    .C(_1075_),
    .Y(_1076_));
 sky130_fd_sc_hd__o2bb2a_1 _2548_ (.A1_N(_1042_),
    .A2_N(_1051_),
    .B1(_1063_),
    .B2(_1076_),
    .X(_1077_));
 sky130_fd_sc_hd__mux4_2 _2549_ (.A0(\tms1x00.RAM[24][3] ),
    .A1(\tms1x00.RAM[25][3] ),
    .A2(\tms1x00.RAM[26][3] ),
    .A3(\tms1x00.RAM[27][3] ),
    .S0(_0760_),
    .S1(_0758_),
    .X(_1078_));
 sky130_fd_sc_hd__mux2_1 _2550_ (.A0(\tms1x00.RAM[30][3] ),
    .A1(\tms1x00.RAM[31][3] ),
    .S(_0760_),
    .X(_1079_));
 sky130_fd_sc_hd__mux2_1 _2551_ (.A0(\tms1x00.RAM[28][3] ),
    .A1(\tms1x00.RAM[29][3] ),
    .S(_0703_),
    .X(_1080_));
 sky130_fd_sc_hd__and2b_1 _2552_ (.A_N(_0767_),
    .B(_1080_),
    .X(_1081_));
 sky130_fd_sc_hd__a211o_1 _2553_ (.A1(_0758_),
    .A2(_1079_),
    .B1(_1081_),
    .C1(_0734_),
    .X(_1082_));
 sky130_fd_sc_hd__o211ai_1 _2554_ (.A1(_0721_),
    .A2(_1078_),
    .B1(_1082_),
    .C1(_0709_),
    .Y(_1083_));
 sky130_fd_sc_hd__mux4_2 _2555_ (.A0(\tms1x00.RAM[16][3] ),
    .A1(\tms1x00.RAM[17][3] ),
    .A2(\tms1x00.RAM[18][3] ),
    .A3(\tms1x00.RAM[19][3] ),
    .S0(_0760_),
    .S1(_0758_),
    .X(_1084_));
 sky130_fd_sc_hd__mux4_1 _2556_ (.A0(\tms1x00.RAM[20][3] ),
    .A1(\tms1x00.RAM[21][3] ),
    .A2(\tms1x00.RAM[22][3] ),
    .A3(\tms1x00.RAM[23][3] ),
    .S0(_0760_),
    .S1(_0702_),
    .X(_1085_));
 sky130_fd_sc_hd__o21a_1 _2557_ (.A1(_0734_),
    .A2(_1085_),
    .B1(_0723_),
    .X(_1086_));
 sky130_fd_sc_hd__o21ai_1 _2558_ (.A1(_0721_),
    .A2(_1084_),
    .B1(_1086_),
    .Y(_1087_));
 sky130_fd_sc_hd__mux2_1 _2559_ (.A0(\tms1x00.RAM[12][3] ),
    .A1(\tms1x00.RAM[13][3] ),
    .S(_0797_),
    .X(_1088_));
 sky130_fd_sc_hd__and2b_1 _2560_ (.A_N(_0767_),
    .B(_1088_),
    .X(_1089_));
 sky130_fd_sc_hd__mux2_1 _2561_ (.A0(\tms1x00.RAM[14][3] ),
    .A1(\tms1x00.RAM[15][3] ),
    .S(_0666_),
    .X(_1090_));
 sky130_fd_sc_hd__a21o_1 _2562_ (.A1(_0664_),
    .A2(_1090_),
    .B1(_0751_),
    .X(_1091_));
 sky130_fd_sc_hd__mux4_1 _2563_ (.A0(\tms1x00.RAM[8][3] ),
    .A1(\tms1x00.RAM[9][3] ),
    .A2(\tms1x00.RAM[10][3] ),
    .A3(\tms1x00.RAM[11][3] ),
    .S0(_0680_),
    .S1(_0775_),
    .X(_1092_));
 sky130_fd_sc_hd__o221a_1 _2564_ (.A1(_1089_),
    .A2(_1091_),
    .B1(_1092_),
    .B2(_0678_),
    .C1(_0709_),
    .X(_1093_));
 sky130_fd_sc_hd__mux2_1 _2565_ (.A0(\tms1x00.RAM[4][3] ),
    .A1(\tms1x00.RAM[5][3] ),
    .S(_0666_),
    .X(_1094_));
 sky130_fd_sc_hd__and2b_1 _2566_ (.A_N(_0702_),
    .B(_1094_),
    .X(_1095_));
 sky130_fd_sc_hd__mux2_1 _2567_ (.A0(\tms1x00.RAM[6][3] ),
    .A1(\tms1x00.RAM[7][3] ),
    .S(_0713_),
    .X(_1096_));
 sky130_fd_sc_hd__a21o_1 _2568_ (.A1(_0660_),
    .A2(_1096_),
    .B1(_0715_),
    .X(_1097_));
 sky130_fd_sc_hd__mux4_1 _2569_ (.A0(\tms1x00.RAM[0][3] ),
    .A1(\tms1x00.RAM[1][3] ),
    .A2(\tms1x00.RAM[2][3] ),
    .A3(\tms1x00.RAM[3][3] ),
    .S0(_0718_),
    .S1(_0682_),
    .X(_1098_));
 sky130_fd_sc_hd__o221a_1 _2570_ (.A1(_1095_),
    .A2(_1097_),
    .B1(_1098_),
    .B2(_0721_),
    .C1(_0723_),
    .X(_1099_));
 sky130_fd_sc_hd__nor3_1 _2571_ (.A(_0695_),
    .B(_1093_),
    .C(_1099_),
    .Y(_1100_));
 sky130_fd_sc_hd__a311o_1 _2572_ (.A1(_0695_),
    .A2(_1083_),
    .A3(_1087_),
    .B1(_1100_),
    .C1(_0657_),
    .X(_1101_));
 sky130_fd_sc_hd__mux2_1 _2573_ (.A0(\tms1x00.RAM[52][3] ),
    .A1(\tms1x00.RAM[53][3] ),
    .S(_0797_),
    .X(_1102_));
 sky130_fd_sc_hd__and2b_1 _2574_ (.A_N(_0697_),
    .B(_1102_),
    .X(_1103_));
 sky130_fd_sc_hd__mux2_1 _2575_ (.A0(\tms1x00.RAM[54][3] ),
    .A1(\tms1x00.RAM[55][3] ),
    .S(_0666_),
    .X(_1104_));
 sky130_fd_sc_hd__a21o_1 _2576_ (.A1(_0702_),
    .A2(_1104_),
    .B1(_0705_),
    .X(_1105_));
 sky130_fd_sc_hd__mux4_1 _2577_ (.A0(\tms1x00.RAM[48][3] ),
    .A1(\tms1x00.RAM[49][3] ),
    .A2(\tms1x00.RAM[50][3] ),
    .A3(\tms1x00.RAM[51][3] ),
    .S0(_0687_),
    .S1(_0688_),
    .X(_1106_));
 sky130_fd_sc_hd__o221a_1 _2578_ (.A1(_1103_),
    .A2(_1105_),
    .B1(_1106_),
    .B2(_0678_),
    .C1(_0691_),
    .X(_1107_));
 sky130_fd_sc_hd__mux4_2 _2579_ (.A0(\tms1x00.RAM[56][3] ),
    .A1(\tms1x00.RAM[57][3] ),
    .A2(\tms1x00.RAM[58][3] ),
    .A3(\tms1x00.RAM[59][3] ),
    .S0(_0718_),
    .S1(_0682_),
    .X(_1108_));
 sky130_fd_sc_hd__mux4_1 _2580_ (.A0(\tms1x00.RAM[60][3] ),
    .A1(\tms1x00.RAM[61][3] ),
    .A2(\tms1x00.RAM[62][3] ),
    .A3(\tms1x00.RAM[63][3] ),
    .S0(_0679_),
    .S1(_0730_),
    .X(_1109_));
 sky130_fd_sc_hd__or2_1 _2581_ (.A(_0751_),
    .B(_1109_),
    .X(_1110_));
 sky130_fd_sc_hd__o211a_1 _2582_ (.A1(_0721_),
    .A2(_1108_),
    .B1(_1110_),
    .C1(_0709_),
    .X(_1111_));
 sky130_fd_sc_hd__mux4_1 _2583_ (.A0(\tms1x00.RAM[44][3] ),
    .A1(\tms1x00.RAM[45][3] ),
    .A2(\tms1x00.RAM[46][3] ),
    .A3(\tms1x00.RAM[47][3] ),
    .S0(_0717_),
    .S1(_0730_),
    .X(_1112_));
 sky130_fd_sc_hd__or2_1 _2584_ (.A(_0751_),
    .B(_1112_),
    .X(_1113_));
 sky130_fd_sc_hd__mux4_1 _2585_ (.A0(\tms1x00.RAM[40][3] ),
    .A1(\tms1x00.RAM[41][3] ),
    .A2(\tms1x00.RAM[42][3] ),
    .A3(\tms1x00.RAM[43][3] ),
    .S0(_0744_),
    .S1(_0696_),
    .X(_1114_));
 sky130_fd_sc_hd__o21a_1 _2586_ (.A1(_0720_),
    .A2(_1114_),
    .B1(_0740_),
    .X(_1115_));
 sky130_fd_sc_hd__mux4_1 _2587_ (.A0(\tms1x00.RAM[32][3] ),
    .A1(\tms1x00.RAM[33][3] ),
    .A2(\tms1x00.RAM[34][3] ),
    .A3(\tms1x00.RAM[35][3] ),
    .S0(_0717_),
    .S1(_0681_),
    .X(_1116_));
 sky130_fd_sc_hd__or2_1 _2588_ (.A(_0720_),
    .B(_1116_),
    .X(_1117_));
 sky130_fd_sc_hd__mux4_1 _2589_ (.A0(\tms1x00.RAM[36][3] ),
    .A1(\tms1x00.RAM[37][3] ),
    .A2(\tms1x00.RAM[38][3] ),
    .A3(\tms1x00.RAM[39][3] ),
    .S0(_0737_),
    .S1(_0696_),
    .X(_1118_));
 sky130_fd_sc_hd__o21a_1 _2590_ (.A1(_0715_),
    .A2(_1118_),
    .B1(_0722_),
    .X(_1119_));
 sky130_fd_sc_hd__a221o_1 _2591_ (.A1(_1113_),
    .A2(_1115_),
    .B1(_1117_),
    .B2(_1119_),
    .C1(_0004_),
    .X(_1120_));
 sky130_fd_sc_hd__o311a_1 _2592_ (.A1(_0754_),
    .A2(_1107_),
    .A3(_1111_),
    .B1(_1120_),
    .C1(_0657_),
    .X(_1121_));
 sky130_fd_sc_hd__nor2_1 _2593_ (.A(_0006_),
    .B(_1121_),
    .Y(_1122_));
 sky130_fd_sc_hd__a22oi_4 _2594_ (.A1(_0006_),
    .A2(_1077_),
    .B1(_1101_),
    .B2(_1122_),
    .Y(_1123_));
 sky130_fd_sc_hd__nand2_1 _2595_ (.A(\tms1x00.ins_in[7] ),
    .B(\tms1x00.ins_in[6] ),
    .Y(_1124_));
 sky130_fd_sc_hd__and3_1 _2596_ (.A(\tms1x00.ins_in[7] ),
    .B(_0637_),
    .C(_0816_),
    .X(_1125_));
 sky130_fd_sc_hd__a221o_1 _2597_ (.A1(\tms1x00.A[3] ),
    .A2(_0818_),
    .B1(_1123_),
    .B2(_1124_),
    .C1(_1125_),
    .X(_1126_));
 sky130_fd_sc_hd__buf_4 _2598_ (.A(_1126_),
    .X(_1127_));
 sky130_fd_sc_hd__buf_4 _2599_ (.A(_1127_),
    .X(_1128_));
 sky130_fd_sc_hd__mux2_1 _2600_ (.A0(_1128_),
    .A1(\tms1x00.RAM[99][3] ),
    .S(_0828_),
    .X(_1129_));
 sky130_fd_sc_hd__clkbuf_1 _2601_ (.A(_1129_),
    .X(_0018_));
 sky130_fd_sc_hd__clkbuf_4 _2602_ (.A(_0820_),
    .X(_1130_));
 sky130_fd_sc_hd__nand3b_4 _2603_ (.A_N(\tms1x00.ram_addr_buff[5] ),
    .B(\tms1x00.ram_addr_buff[6] ),
    .C(\tms1x00.ram_addr_buff[4] ),
    .Y(_1131_));
 sky130_fd_sc_hd__buf_4 _2604_ (.A(_1131_),
    .X(_1132_));
 sky130_fd_sc_hd__or3b_1 _2605_ (.A(\tms1x00.ram_addr_buff[2] ),
    .B(_0825_),
    .C_N(\tms1x00.ram_addr_buff[3] ),
    .X(_1133_));
 sky130_fd_sc_hd__or3b_1 _2606_ (.A(\tms1x00.ram_addr_buff[1] ),
    .B(_1133_),
    .C_N(\tms1x00.ram_addr_buff[0] ),
    .X(_1134_));
 sky130_fd_sc_hd__buf_4 _2607_ (.A(_1134_),
    .X(_1135_));
 sky130_fd_sc_hd__nor2_2 _2608_ (.A(_1132_),
    .B(_1135_),
    .Y(_1136_));
 sky130_fd_sc_hd__mux2_1 _2609_ (.A0(\tms1x00.RAM[89][0] ),
    .A1(_1130_),
    .S(_1136_),
    .X(_1137_));
 sky130_fd_sc_hd__clkbuf_1 _2610_ (.A(_1137_),
    .X(_0019_));
 sky130_fd_sc_hd__clkbuf_4 _2611_ (.A(_0929_),
    .X(_1138_));
 sky130_fd_sc_hd__mux2_1 _2612_ (.A0(\tms1x00.RAM[89][1] ),
    .A1(_1138_),
    .S(_1136_),
    .X(_1139_));
 sky130_fd_sc_hd__clkbuf_1 _2613_ (.A(_1139_),
    .X(_0020_));
 sky130_fd_sc_hd__clkbuf_4 _2614_ (.A(_1029_),
    .X(_1140_));
 sky130_fd_sc_hd__mux2_1 _2615_ (.A0(\tms1x00.RAM[89][2] ),
    .A1(_1140_),
    .S(_1136_),
    .X(_1141_));
 sky130_fd_sc_hd__clkbuf_1 _2616_ (.A(_1141_),
    .X(_0021_));
 sky130_fd_sc_hd__clkbuf_4 _2617_ (.A(_1127_),
    .X(_1142_));
 sky130_fd_sc_hd__mux2_1 _2618_ (.A0(\tms1x00.RAM[89][3] ),
    .A1(_1142_),
    .S(_1136_),
    .X(_1143_));
 sky130_fd_sc_hd__clkbuf_1 _2619_ (.A(_1143_),
    .X(_0022_));
 sky130_fd_sc_hd__nand3b_2 _2620_ (.A_N(\tms1x00.ram_addr_buff[6] ),
    .B(\tms1x00.ram_addr_buff[5] ),
    .C(\tms1x00.ram_addr_buff[4] ),
    .Y(_1144_));
 sky130_fd_sc_hd__buf_4 _2621_ (.A(_1144_),
    .X(_1145_));
 sky130_fd_sc_hd__or2_1 _2622_ (.A(_0824_),
    .B(_1133_),
    .X(_1146_));
 sky130_fd_sc_hd__buf_6 _2623_ (.A(_1146_),
    .X(_1147_));
 sky130_fd_sc_hd__nor2_2 _2624_ (.A(_1145_),
    .B(_1147_),
    .Y(_1148_));
 sky130_fd_sc_hd__mux2_1 _2625_ (.A0(\tms1x00.RAM[59][0] ),
    .A1(_1130_),
    .S(_1148_),
    .X(_1149_));
 sky130_fd_sc_hd__clkbuf_1 _2626_ (.A(_1149_),
    .X(_0023_));
 sky130_fd_sc_hd__mux2_1 _2627_ (.A0(\tms1x00.RAM[59][1] ),
    .A1(_1138_),
    .S(_1148_),
    .X(_1150_));
 sky130_fd_sc_hd__clkbuf_1 _2628_ (.A(_1150_),
    .X(_0024_));
 sky130_fd_sc_hd__mux2_1 _2629_ (.A0(\tms1x00.RAM[59][2] ),
    .A1(_1140_),
    .S(_1148_),
    .X(_1151_));
 sky130_fd_sc_hd__clkbuf_1 _2630_ (.A(_1151_),
    .X(_0025_));
 sky130_fd_sc_hd__mux2_1 _2631_ (.A0(\tms1x00.RAM[59][3] ),
    .A1(_1142_),
    .S(_1148_),
    .X(_1152_));
 sky130_fd_sc_hd__clkbuf_1 _2632_ (.A(_1152_),
    .X(_0026_));
 sky130_fd_sc_hd__and3b_2 _2633_ (.A_N(_0825_),
    .B(\tms1x00.ram_addr_buff[3] ),
    .C(\tms1x00.ram_addr_buff[2] ),
    .X(_1153_));
 sky130_fd_sc_hd__nand3b_4 _2634_ (.A_N(_0625_),
    .B(_1153_),
    .C(_0617_),
    .Y(_1154_));
 sky130_fd_sc_hd__or2_2 _2635_ (.A(_0823_),
    .B(_1154_),
    .X(_1155_));
 sky130_fd_sc_hd__mux2_1 _2636_ (.A0(_0821_),
    .A1(\tms1x00.RAM[109][0] ),
    .S(_1155_),
    .X(_1156_));
 sky130_fd_sc_hd__clkbuf_1 _2637_ (.A(_1156_),
    .X(_0027_));
 sky130_fd_sc_hd__mux2_1 _2638_ (.A0(_0930_),
    .A1(\tms1x00.RAM[109][1] ),
    .S(_1155_),
    .X(_1157_));
 sky130_fd_sc_hd__clkbuf_1 _2639_ (.A(_1157_),
    .X(_0028_));
 sky130_fd_sc_hd__mux2_1 _2640_ (.A0(_1030_),
    .A1(\tms1x00.RAM[109][2] ),
    .S(_1155_),
    .X(_1158_));
 sky130_fd_sc_hd__clkbuf_1 _2641_ (.A(_1158_),
    .X(_0029_));
 sky130_fd_sc_hd__mux2_1 _2642_ (.A0(_1128_),
    .A1(\tms1x00.RAM[109][3] ),
    .S(_1155_),
    .X(_1159_));
 sky130_fd_sc_hd__clkbuf_1 _2643_ (.A(_1159_),
    .X(_0030_));
 sky130_fd_sc_hd__or3b_4 _2644_ (.A(\tms1x00.ram_addr_buff[4] ),
    .B(\tms1x00.ram_addr_buff[5] ),
    .C_N(\tms1x00.ram_addr_buff[6] ),
    .X(_1160_));
 sky130_fd_sc_hd__buf_4 _2645_ (.A(_1160_),
    .X(_1161_));
 sky130_fd_sc_hd__or2b_1 _2646_ (.A(\tms1x00.ram_addr_buff[3] ),
    .B_N(\tms1x00.ram_addr_buff[2] ),
    .X(_1162_));
 sky130_fd_sc_hd__or4b_4 _2647_ (.A(\tms1x00.ram_addr_buff[1] ),
    .B(_0825_),
    .C(_1162_),
    .D_N(\tms1x00.ram_addr_buff[0] ),
    .X(_1163_));
 sky130_fd_sc_hd__or2_2 _2648_ (.A(_1161_),
    .B(_1163_),
    .X(_1164_));
 sky130_fd_sc_hd__mux2_1 _2649_ (.A0(_0821_),
    .A1(\tms1x00.RAM[69][0] ),
    .S(_1164_),
    .X(_1165_));
 sky130_fd_sc_hd__clkbuf_1 _2650_ (.A(_1165_),
    .X(_0031_));
 sky130_fd_sc_hd__mux2_1 _2651_ (.A0(_0930_),
    .A1(\tms1x00.RAM[69][1] ),
    .S(_1164_),
    .X(_1166_));
 sky130_fd_sc_hd__clkbuf_1 _2652_ (.A(_1166_),
    .X(_0032_));
 sky130_fd_sc_hd__mux2_1 _2653_ (.A0(_1030_),
    .A1(\tms1x00.RAM[69][2] ),
    .S(_1164_),
    .X(_1167_));
 sky130_fd_sc_hd__clkbuf_1 _2654_ (.A(_1167_),
    .X(_0033_));
 sky130_fd_sc_hd__mux2_1 _2655_ (.A0(_1128_),
    .A1(\tms1x00.RAM[69][3] ),
    .S(_1164_),
    .X(_1168_));
 sky130_fd_sc_hd__clkbuf_1 _2656_ (.A(_1168_),
    .X(_0034_));
 sky130_fd_sc_hd__or2b_4 _2657_ (.A(_0824_),
    .B_N(_1153_),
    .X(_1169_));
 sky130_fd_sc_hd__or2_2 _2658_ (.A(_1161_),
    .B(_1169_),
    .X(_1170_));
 sky130_fd_sc_hd__mux2_1 _2659_ (.A0(_0821_),
    .A1(\tms1x00.RAM[79][0] ),
    .S(_1170_),
    .X(_1171_));
 sky130_fd_sc_hd__clkbuf_1 _2660_ (.A(_1171_),
    .X(_0035_));
 sky130_fd_sc_hd__mux2_1 _2661_ (.A0(_0930_),
    .A1(\tms1x00.RAM[79][1] ),
    .S(_1170_),
    .X(_1172_));
 sky130_fd_sc_hd__clkbuf_1 _2662_ (.A(_1172_),
    .X(_0036_));
 sky130_fd_sc_hd__mux2_1 _2663_ (.A0(_1030_),
    .A1(\tms1x00.RAM[79][2] ),
    .S(_1170_),
    .X(_1173_));
 sky130_fd_sc_hd__clkbuf_1 _2664_ (.A(_1173_),
    .X(_0037_));
 sky130_fd_sc_hd__mux2_1 _2665_ (.A0(_1128_),
    .A1(\tms1x00.RAM[79][3] ),
    .S(_1170_),
    .X(_1174_));
 sky130_fd_sc_hd__clkbuf_1 _2666_ (.A(_1174_),
    .X(_0038_));
 sky130_fd_sc_hd__nand3_4 _2667_ (.A(\tms1x00.ram_addr_buff[4] ),
    .B(\tms1x00.ram_addr_buff[5] ),
    .C(\tms1x00.ram_addr_buff[6] ),
    .Y(_1175_));
 sky130_fd_sc_hd__clkbuf_4 _2668_ (.A(_1175_),
    .X(_1176_));
 sky130_fd_sc_hd__or2_2 _2669_ (.A(_1169_),
    .B(_1176_),
    .X(_1177_));
 sky130_fd_sc_hd__mux2_1 _2670_ (.A0(_0821_),
    .A1(\tms1x00.RAM[127][0] ),
    .S(_1177_),
    .X(_1178_));
 sky130_fd_sc_hd__clkbuf_1 _2671_ (.A(_1178_),
    .X(_0039_));
 sky130_fd_sc_hd__mux2_1 _2672_ (.A0(_0930_),
    .A1(\tms1x00.RAM[127][1] ),
    .S(_1177_),
    .X(_1179_));
 sky130_fd_sc_hd__clkbuf_1 _2673_ (.A(_1179_),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_1 _2674_ (.A0(_1030_),
    .A1(\tms1x00.RAM[127][2] ),
    .S(_1177_),
    .X(_1180_));
 sky130_fd_sc_hd__clkbuf_1 _2675_ (.A(_1180_),
    .X(_0041_));
 sky130_fd_sc_hd__mux2_1 _2676_ (.A0(_1128_),
    .A1(\tms1x00.RAM[127][3] ),
    .S(_1177_),
    .X(_1181_));
 sky130_fd_sc_hd__clkbuf_1 _2677_ (.A(_1181_),
    .X(_0042_));
 sky130_fd_sc_hd__or3b_4 _2678_ (.A(_0625_),
    .B(_0826_),
    .C_N(_0617_),
    .X(_1182_));
 sky130_fd_sc_hd__or2_2 _2679_ (.A(_1145_),
    .B(_1182_),
    .X(_1183_));
 sky130_fd_sc_hd__mux2_1 _2680_ (.A0(_0821_),
    .A1(\tms1x00.RAM[49][0] ),
    .S(_1183_),
    .X(_1184_));
 sky130_fd_sc_hd__clkbuf_1 _2681_ (.A(_1184_),
    .X(_0043_));
 sky130_fd_sc_hd__mux2_1 _2682_ (.A0(_0930_),
    .A1(\tms1x00.RAM[49][1] ),
    .S(_1183_),
    .X(_1185_));
 sky130_fd_sc_hd__clkbuf_1 _2683_ (.A(_1185_),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _2684_ (.A0(_1030_),
    .A1(\tms1x00.RAM[49][2] ),
    .S(_1183_),
    .X(_1186_));
 sky130_fd_sc_hd__clkbuf_1 _2685_ (.A(_1186_),
    .X(_0045_));
 sky130_fd_sc_hd__mux2_1 _2686_ (.A0(_1128_),
    .A1(\tms1x00.RAM[49][3] ),
    .S(_1183_),
    .X(_1187_));
 sky130_fd_sc_hd__clkbuf_1 _2687_ (.A(_1187_),
    .X(_0046_));
 sky130_fd_sc_hd__or3b_4 _2688_ (.A(\tms1x00.ram_addr_buff[5] ),
    .B(\tms1x00.ram_addr_buff[6] ),
    .C_N(\tms1x00.ram_addr_buff[4] ),
    .X(_1188_));
 sky130_fd_sc_hd__or2_2 _2689_ (.A(_0827_),
    .B(_1188_),
    .X(_1189_));
 sky130_fd_sc_hd__mux2_1 _2690_ (.A0(_0821_),
    .A1(\tms1x00.RAM[19][0] ),
    .S(_1189_),
    .X(_1190_));
 sky130_fd_sc_hd__clkbuf_1 _2691_ (.A(_1190_),
    .X(_0047_));
 sky130_fd_sc_hd__mux2_1 _2692_ (.A0(_0930_),
    .A1(\tms1x00.RAM[19][1] ),
    .S(_1189_),
    .X(_1191_));
 sky130_fd_sc_hd__clkbuf_1 _2693_ (.A(_1191_),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _2694_ (.A0(_1030_),
    .A1(\tms1x00.RAM[19][2] ),
    .S(_1189_),
    .X(_1192_));
 sky130_fd_sc_hd__clkbuf_1 _2695_ (.A(_1192_),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_1 _2696_ (.A0(_1128_),
    .A1(\tms1x00.RAM[19][3] ),
    .S(_1189_),
    .X(_1193_));
 sky130_fd_sc_hd__clkbuf_1 _2697_ (.A(_1193_),
    .X(_0050_));
 sky130_fd_sc_hd__or2_2 _2698_ (.A(_1132_),
    .B(_1169_),
    .X(_1194_));
 sky130_fd_sc_hd__mux2_1 _2699_ (.A0(_0821_),
    .A1(\tms1x00.RAM[95][0] ),
    .S(_1194_),
    .X(_1195_));
 sky130_fd_sc_hd__clkbuf_1 _2700_ (.A(_1195_),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _2701_ (.A0(_0930_),
    .A1(\tms1x00.RAM[95][1] ),
    .S(_1194_),
    .X(_1196_));
 sky130_fd_sc_hd__clkbuf_1 _2702_ (.A(_1196_),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _2703_ (.A0(_1030_),
    .A1(\tms1x00.RAM[95][2] ),
    .S(_1194_),
    .X(_1197_));
 sky130_fd_sc_hd__clkbuf_1 _2704_ (.A(_1197_),
    .X(_0053_));
 sky130_fd_sc_hd__mux2_1 _2705_ (.A0(_1128_),
    .A1(\tms1x00.RAM[95][3] ),
    .S(_1194_),
    .X(_1198_));
 sky130_fd_sc_hd__clkbuf_1 _2706_ (.A(_1198_),
    .X(_0054_));
 sky130_fd_sc_hd__nand3b_4 _2707_ (.A_N(_0617_),
    .B(_0625_),
    .C(_1153_),
    .Y(_1199_));
 sky130_fd_sc_hd__or2_2 _2708_ (.A(_1132_),
    .B(_1199_),
    .X(_1200_));
 sky130_fd_sc_hd__mux2_1 _2709_ (.A0(_0821_),
    .A1(\tms1x00.RAM[94][0] ),
    .S(_1200_),
    .X(_1201_));
 sky130_fd_sc_hd__clkbuf_1 _2710_ (.A(_1201_),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _2711_ (.A0(_0930_),
    .A1(\tms1x00.RAM[94][1] ),
    .S(_1200_),
    .X(_1202_));
 sky130_fd_sc_hd__clkbuf_1 _2712_ (.A(_1202_),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _2713_ (.A0(_1030_),
    .A1(\tms1x00.RAM[94][2] ),
    .S(_1200_),
    .X(_1203_));
 sky130_fd_sc_hd__clkbuf_1 _2714_ (.A(_1203_),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _2715_ (.A0(_1128_),
    .A1(\tms1x00.RAM[94][3] ),
    .S(_1200_),
    .X(_1204_));
 sky130_fd_sc_hd__clkbuf_1 _2716_ (.A(_1204_),
    .X(_0058_));
 sky130_fd_sc_hd__or2_2 _2717_ (.A(_1132_),
    .B(_1154_),
    .X(_1205_));
 sky130_fd_sc_hd__mux2_1 _2718_ (.A0(_0821_),
    .A1(\tms1x00.RAM[93][0] ),
    .S(_1205_),
    .X(_1206_));
 sky130_fd_sc_hd__clkbuf_1 _2719_ (.A(_1206_),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _2720_ (.A0(_0930_),
    .A1(\tms1x00.RAM[93][1] ),
    .S(_1205_),
    .X(_1207_));
 sky130_fd_sc_hd__clkbuf_1 _2721_ (.A(_1207_),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _2722_ (.A0(_1030_),
    .A1(\tms1x00.RAM[93][2] ),
    .S(_1205_),
    .X(_1208_));
 sky130_fd_sc_hd__clkbuf_1 _2723_ (.A(_1208_),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _2724_ (.A0(_1128_),
    .A1(\tms1x00.RAM[93][3] ),
    .S(_1205_),
    .X(_1209_));
 sky130_fd_sc_hd__clkbuf_1 _2725_ (.A(_1209_),
    .X(_0062_));
 sky130_fd_sc_hd__buf_4 _2726_ (.A(_0820_),
    .X(_1210_));
 sky130_fd_sc_hd__or3b_4 _2727_ (.A(_0617_),
    .B(_0625_),
    .C_N(_1153_),
    .X(_1211_));
 sky130_fd_sc_hd__or2_2 _2728_ (.A(_1132_),
    .B(_1211_),
    .X(_1212_));
 sky130_fd_sc_hd__mux2_1 _2729_ (.A0(_1210_),
    .A1(\tms1x00.RAM[92][0] ),
    .S(_1212_),
    .X(_1213_));
 sky130_fd_sc_hd__clkbuf_1 _2730_ (.A(_1213_),
    .X(_0063_));
 sky130_fd_sc_hd__buf_4 _2731_ (.A(_0929_),
    .X(_1214_));
 sky130_fd_sc_hd__mux2_1 _2732_ (.A0(_1214_),
    .A1(\tms1x00.RAM[92][1] ),
    .S(_1212_),
    .X(_1215_));
 sky130_fd_sc_hd__clkbuf_1 _2733_ (.A(_1215_),
    .X(_0064_));
 sky130_fd_sc_hd__buf_4 _2734_ (.A(_1029_),
    .X(_1216_));
 sky130_fd_sc_hd__mux2_1 _2735_ (.A0(_1216_),
    .A1(\tms1x00.RAM[92][2] ),
    .S(_1212_),
    .X(_1217_));
 sky130_fd_sc_hd__clkbuf_1 _2736_ (.A(_1217_),
    .X(_0065_));
 sky130_fd_sc_hd__clkbuf_4 _2737_ (.A(_1127_),
    .X(_1218_));
 sky130_fd_sc_hd__mux2_1 _2738_ (.A0(_1218_),
    .A1(\tms1x00.RAM[92][3] ),
    .S(_1212_),
    .X(_1219_));
 sky130_fd_sc_hd__clkbuf_1 _2739_ (.A(_1219_),
    .X(_0066_));
 sky130_fd_sc_hd__nor2_2 _2740_ (.A(_1132_),
    .B(_1147_),
    .Y(_1220_));
 sky130_fd_sc_hd__mux2_1 _2741_ (.A0(\tms1x00.RAM[91][0] ),
    .A1(_1130_),
    .S(_1220_),
    .X(_1221_));
 sky130_fd_sc_hd__clkbuf_1 _2742_ (.A(_1221_),
    .X(_0067_));
 sky130_fd_sc_hd__mux2_1 _2743_ (.A0(\tms1x00.RAM[91][1] ),
    .A1(_1138_),
    .S(_1220_),
    .X(_1222_));
 sky130_fd_sc_hd__clkbuf_1 _2744_ (.A(_1222_),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _2745_ (.A0(\tms1x00.RAM[91][2] ),
    .A1(_1140_),
    .S(_1220_),
    .X(_1223_));
 sky130_fd_sc_hd__clkbuf_1 _2746_ (.A(_1223_),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_1 _2747_ (.A0(\tms1x00.RAM[91][3] ),
    .A1(_1142_),
    .S(_1220_),
    .X(_1224_));
 sky130_fd_sc_hd__clkbuf_1 _2748_ (.A(_1224_),
    .X(_0070_));
 sky130_fd_sc_hd__or3b_1 _2749_ (.A(_1133_),
    .B(\tms1x00.ram_addr_buff[0] ),
    .C_N(\tms1x00.ram_addr_buff[1] ),
    .X(_1225_));
 sky130_fd_sc_hd__buf_4 _2750_ (.A(_1225_),
    .X(_1226_));
 sky130_fd_sc_hd__nor2_2 _2751_ (.A(_1132_),
    .B(_1226_),
    .Y(_1227_));
 sky130_fd_sc_hd__mux2_1 _2752_ (.A0(\tms1x00.RAM[90][0] ),
    .A1(_1130_),
    .S(_1227_),
    .X(_1228_));
 sky130_fd_sc_hd__clkbuf_1 _2753_ (.A(_1228_),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _2754_ (.A0(\tms1x00.RAM[90][1] ),
    .A1(_1138_),
    .S(_1227_),
    .X(_1229_));
 sky130_fd_sc_hd__clkbuf_1 _2755_ (.A(_1229_),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_1 _2756_ (.A0(\tms1x00.RAM[90][2] ),
    .A1(_1140_),
    .S(_1227_),
    .X(_1230_));
 sky130_fd_sc_hd__clkbuf_1 _2757_ (.A(_1230_),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _2758_ (.A0(\tms1x00.RAM[90][3] ),
    .A1(_1142_),
    .S(_1227_),
    .X(_1231_));
 sky130_fd_sc_hd__clkbuf_1 _2759_ (.A(_1231_),
    .X(_0074_));
 sky130_fd_sc_hd__or3_4 _2760_ (.A(\tms1x00.ram_addr_buff[4] ),
    .B(\tms1x00.ram_addr_buff[5] ),
    .C(\tms1x00.ram_addr_buff[6] ),
    .X(_1232_));
 sky130_fd_sc_hd__buf_4 _2761_ (.A(_1232_),
    .X(_1233_));
 sky130_fd_sc_hd__or3_1 _2762_ (.A(\tms1x00.ram_addr_buff[0] ),
    .B(\tms1x00.ram_addr_buff[1] ),
    .C(_1133_),
    .X(_1234_));
 sky130_fd_sc_hd__buf_4 _2763_ (.A(_1234_),
    .X(_1235_));
 sky130_fd_sc_hd__nor2_2 _2764_ (.A(_1233_),
    .B(_1235_),
    .Y(_1236_));
 sky130_fd_sc_hd__mux2_1 _2765_ (.A0(\tms1x00.RAM[8][0] ),
    .A1(_1130_),
    .S(_1236_),
    .X(_1237_));
 sky130_fd_sc_hd__clkbuf_1 _2766_ (.A(_1237_),
    .X(_0075_));
 sky130_fd_sc_hd__mux2_1 _2767_ (.A0(\tms1x00.RAM[8][1] ),
    .A1(_1138_),
    .S(_1236_),
    .X(_1238_));
 sky130_fd_sc_hd__clkbuf_1 _2768_ (.A(_1238_),
    .X(_0076_));
 sky130_fd_sc_hd__mux2_1 _2769_ (.A0(\tms1x00.RAM[8][2] ),
    .A1(_1140_),
    .S(_1236_),
    .X(_1239_));
 sky130_fd_sc_hd__clkbuf_1 _2770_ (.A(_1239_),
    .X(_0077_));
 sky130_fd_sc_hd__mux2_1 _2771_ (.A0(\tms1x00.RAM[8][3] ),
    .A1(_1142_),
    .S(_1236_),
    .X(_1240_));
 sky130_fd_sc_hd__clkbuf_1 _2772_ (.A(_1240_),
    .X(_0078_));
 sky130_fd_sc_hd__nor2_2 _2773_ (.A(_1132_),
    .B(_1235_),
    .Y(_1241_));
 sky130_fd_sc_hd__mux2_1 _2774_ (.A0(\tms1x00.RAM[88][0] ),
    .A1(_1130_),
    .S(_1241_),
    .X(_1242_));
 sky130_fd_sc_hd__clkbuf_1 _2775_ (.A(_1242_),
    .X(_0079_));
 sky130_fd_sc_hd__mux2_1 _2776_ (.A0(\tms1x00.RAM[88][1] ),
    .A1(_1138_),
    .S(_1241_),
    .X(_1243_));
 sky130_fd_sc_hd__clkbuf_1 _2777_ (.A(_1243_),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _2778_ (.A0(\tms1x00.RAM[88][2] ),
    .A1(_1140_),
    .S(_1241_),
    .X(_1244_));
 sky130_fd_sc_hd__clkbuf_1 _2779_ (.A(_1244_),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_1 _2780_ (.A0(\tms1x00.RAM[88][3] ),
    .A1(_1142_),
    .S(_1241_),
    .X(_1245_));
 sky130_fd_sc_hd__clkbuf_1 _2781_ (.A(_1245_),
    .X(_0082_));
 sky130_fd_sc_hd__or3_1 _2782_ (.A(_0824_),
    .B(_0825_),
    .C(_1162_),
    .X(_1246_));
 sky130_fd_sc_hd__buf_6 _2783_ (.A(_1246_),
    .X(_1247_));
 sky130_fd_sc_hd__nor2_2 _2784_ (.A(_1132_),
    .B(_1247_),
    .Y(_1248_));
 sky130_fd_sc_hd__mux2_1 _2785_ (.A0(\tms1x00.RAM[87][0] ),
    .A1(_1130_),
    .S(_1248_),
    .X(_1249_));
 sky130_fd_sc_hd__clkbuf_1 _2786_ (.A(_1249_),
    .X(_0083_));
 sky130_fd_sc_hd__mux2_1 _2787_ (.A0(\tms1x00.RAM[87][1] ),
    .A1(_1138_),
    .S(_1248_),
    .X(_1250_));
 sky130_fd_sc_hd__clkbuf_1 _2788_ (.A(_1250_),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_1 _2789_ (.A0(\tms1x00.RAM[87][2] ),
    .A1(_1140_),
    .S(_1248_),
    .X(_1251_));
 sky130_fd_sc_hd__clkbuf_1 _2790_ (.A(_1251_),
    .X(_0085_));
 sky130_fd_sc_hd__mux2_1 _2791_ (.A0(\tms1x00.RAM[87][3] ),
    .A1(_1142_),
    .S(_1248_),
    .X(_1252_));
 sky130_fd_sc_hd__clkbuf_1 _2792_ (.A(_1252_),
    .X(_0086_));
 sky130_fd_sc_hd__or2_1 _2793_ (.A(_0825_),
    .B(_1162_),
    .X(_1253_));
 sky130_fd_sc_hd__or3b_4 _2794_ (.A(_1253_),
    .B(_0617_),
    .C_N(_0625_),
    .X(_1254_));
 sky130_fd_sc_hd__or2_2 _2795_ (.A(_1132_),
    .B(_1254_),
    .X(_1255_));
 sky130_fd_sc_hd__mux2_1 _2796_ (.A0(_1210_),
    .A1(\tms1x00.RAM[86][0] ),
    .S(_1255_),
    .X(_1256_));
 sky130_fd_sc_hd__clkbuf_1 _2797_ (.A(_1256_),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_1 _2798_ (.A0(_1214_),
    .A1(\tms1x00.RAM[86][1] ),
    .S(_1255_),
    .X(_1257_));
 sky130_fd_sc_hd__clkbuf_1 _2799_ (.A(_1257_),
    .X(_0088_));
 sky130_fd_sc_hd__mux2_1 _2800_ (.A0(_1216_),
    .A1(\tms1x00.RAM[86][2] ),
    .S(_1255_),
    .X(_1258_));
 sky130_fd_sc_hd__clkbuf_1 _2801_ (.A(_1258_),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _2802_ (.A0(_1218_),
    .A1(\tms1x00.RAM[86][3] ),
    .S(_1255_),
    .X(_1259_));
 sky130_fd_sc_hd__clkbuf_1 _2803_ (.A(_1259_),
    .X(_0090_));
 sky130_fd_sc_hd__nor2_2 _2804_ (.A(_0823_),
    .B(_1135_),
    .Y(_1260_));
 sky130_fd_sc_hd__mux2_1 _2805_ (.A0(\tms1x00.RAM[105][0] ),
    .A1(_1130_),
    .S(_1260_),
    .X(_1261_));
 sky130_fd_sc_hd__clkbuf_1 _2806_ (.A(_1261_),
    .X(_0091_));
 sky130_fd_sc_hd__mux2_1 _2807_ (.A0(\tms1x00.RAM[105][1] ),
    .A1(_1138_),
    .S(_1260_),
    .X(_1262_));
 sky130_fd_sc_hd__clkbuf_1 _2808_ (.A(_1262_),
    .X(_0092_));
 sky130_fd_sc_hd__mux2_1 _2809_ (.A0(\tms1x00.RAM[105][2] ),
    .A1(_1140_),
    .S(_1260_),
    .X(_1263_));
 sky130_fd_sc_hd__clkbuf_1 _2810_ (.A(_1263_),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _2811_ (.A0(\tms1x00.RAM[105][3] ),
    .A1(_1142_),
    .S(_1260_),
    .X(_1264_));
 sky130_fd_sc_hd__clkbuf_1 _2812_ (.A(_1264_),
    .X(_0094_));
 sky130_fd_sc_hd__clkbuf_4 _2813_ (.A(_0819_),
    .X(_1265_));
 sky130_fd_sc_hd__buf_4 _2814_ (.A(_1265_),
    .X(_1266_));
 sky130_fd_sc_hd__nor2_2 _2815_ (.A(_0823_),
    .B(_1235_),
    .Y(_1267_));
 sky130_fd_sc_hd__mux2_1 _2816_ (.A0(\tms1x00.RAM[104][0] ),
    .A1(_1266_),
    .S(_1267_),
    .X(_1268_));
 sky130_fd_sc_hd__clkbuf_1 _2817_ (.A(_1268_),
    .X(_0095_));
 sky130_fd_sc_hd__buf_4 _2818_ (.A(_0928_),
    .X(_1269_));
 sky130_fd_sc_hd__clkbuf_4 _2819_ (.A(_1269_),
    .X(_1270_));
 sky130_fd_sc_hd__mux2_1 _2820_ (.A0(\tms1x00.RAM[104][1] ),
    .A1(_1270_),
    .S(_1267_),
    .X(_1271_));
 sky130_fd_sc_hd__clkbuf_1 _2821_ (.A(_1271_),
    .X(_0096_));
 sky130_fd_sc_hd__buf_4 _2822_ (.A(_1028_),
    .X(_1272_));
 sky130_fd_sc_hd__buf_4 _2823_ (.A(_1272_),
    .X(_1273_));
 sky130_fd_sc_hd__mux2_1 _2824_ (.A0(\tms1x00.RAM[104][2] ),
    .A1(_1273_),
    .S(_1267_),
    .X(_1274_));
 sky130_fd_sc_hd__clkbuf_1 _2825_ (.A(_1274_),
    .X(_0097_));
 sky130_fd_sc_hd__buf_4 _2826_ (.A(_1126_),
    .X(_1275_));
 sky130_fd_sc_hd__clkbuf_4 _2827_ (.A(_1275_),
    .X(_1276_));
 sky130_fd_sc_hd__mux2_1 _2828_ (.A0(\tms1x00.RAM[104][3] ),
    .A1(_1276_),
    .S(_1267_),
    .X(_1277_));
 sky130_fd_sc_hd__clkbuf_1 _2829_ (.A(_1277_),
    .X(_0098_));
 sky130_fd_sc_hd__nor2_2 _2830_ (.A(_0823_),
    .B(_1247_),
    .Y(_1278_));
 sky130_fd_sc_hd__mux2_1 _2831_ (.A0(\tms1x00.RAM[103][0] ),
    .A1(_1266_),
    .S(_1278_),
    .X(_1279_));
 sky130_fd_sc_hd__clkbuf_1 _2832_ (.A(_1279_),
    .X(_0099_));
 sky130_fd_sc_hd__mux2_1 _2833_ (.A0(\tms1x00.RAM[103][1] ),
    .A1(_1270_),
    .S(_1278_),
    .X(_1280_));
 sky130_fd_sc_hd__clkbuf_1 _2834_ (.A(_1280_),
    .X(_0100_));
 sky130_fd_sc_hd__mux2_1 _2835_ (.A0(\tms1x00.RAM[103][2] ),
    .A1(_1273_),
    .S(_1278_),
    .X(_1281_));
 sky130_fd_sc_hd__clkbuf_1 _2836_ (.A(_1281_),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _2837_ (.A0(\tms1x00.RAM[103][3] ),
    .A1(_1276_),
    .S(_1278_),
    .X(_1282_));
 sky130_fd_sc_hd__clkbuf_1 _2838_ (.A(_1282_),
    .X(_0102_));
 sky130_fd_sc_hd__or2_2 _2839_ (.A(_0823_),
    .B(_1254_),
    .X(_1283_));
 sky130_fd_sc_hd__mux2_1 _2840_ (.A0(_1210_),
    .A1(\tms1x00.RAM[102][0] ),
    .S(_1283_),
    .X(_1284_));
 sky130_fd_sc_hd__clkbuf_1 _2841_ (.A(_1284_),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _2842_ (.A0(_1214_),
    .A1(\tms1x00.RAM[102][1] ),
    .S(_1283_),
    .X(_1285_));
 sky130_fd_sc_hd__clkbuf_1 _2843_ (.A(_1285_),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _2844_ (.A0(_1216_),
    .A1(\tms1x00.RAM[102][2] ),
    .S(_1283_),
    .X(_1286_));
 sky130_fd_sc_hd__clkbuf_1 _2845_ (.A(_1286_),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _2846_ (.A0(_1218_),
    .A1(\tms1x00.RAM[102][3] ),
    .S(_1283_),
    .X(_1287_));
 sky130_fd_sc_hd__clkbuf_1 _2847_ (.A(_1287_),
    .X(_0106_));
 sky130_fd_sc_hd__or2_2 _2848_ (.A(_0823_),
    .B(_1163_),
    .X(_1288_));
 sky130_fd_sc_hd__mux2_1 _2849_ (.A0(_1210_),
    .A1(\tms1x00.RAM[101][0] ),
    .S(_1288_),
    .X(_1289_));
 sky130_fd_sc_hd__clkbuf_1 _2850_ (.A(_1289_),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _2851_ (.A0(_1214_),
    .A1(\tms1x00.RAM[101][1] ),
    .S(_1288_),
    .X(_1290_));
 sky130_fd_sc_hd__clkbuf_1 _2852_ (.A(_1290_),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _2853_ (.A0(_1216_),
    .A1(\tms1x00.RAM[101][2] ),
    .S(_1288_),
    .X(_1291_));
 sky130_fd_sc_hd__clkbuf_1 _2854_ (.A(_1291_),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _2855_ (.A0(_1218_),
    .A1(\tms1x00.RAM[101][3] ),
    .S(_1288_),
    .X(_1292_));
 sky130_fd_sc_hd__clkbuf_1 _2856_ (.A(_1292_),
    .X(_0110_));
 sky130_fd_sc_hd__or3_4 _2857_ (.A(_0617_),
    .B(_0625_),
    .C(_1253_),
    .X(_1293_));
 sky130_fd_sc_hd__or2_2 _2858_ (.A(_0823_),
    .B(_1293_),
    .X(_1294_));
 sky130_fd_sc_hd__mux2_1 _2859_ (.A0(_1210_),
    .A1(\tms1x00.RAM[100][0] ),
    .S(_1294_),
    .X(_1295_));
 sky130_fd_sc_hd__clkbuf_1 _2860_ (.A(_1295_),
    .X(_0111_));
 sky130_fd_sc_hd__mux2_1 _2861_ (.A0(_1214_),
    .A1(\tms1x00.RAM[100][1] ),
    .S(_1294_),
    .X(_1296_));
 sky130_fd_sc_hd__clkbuf_1 _2862_ (.A(_1296_),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _2863_ (.A0(_1216_),
    .A1(\tms1x00.RAM[100][2] ),
    .S(_1294_),
    .X(_1297_));
 sky130_fd_sc_hd__clkbuf_1 _2864_ (.A(_1297_),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _2865_ (.A0(_1218_),
    .A1(\tms1x00.RAM[100][3] ),
    .S(_1294_),
    .X(_1298_));
 sky130_fd_sc_hd__clkbuf_1 _2866_ (.A(_1298_),
    .X(_0114_));
 sky130_fd_sc_hd__or3_4 _2867_ (.A(_0617_),
    .B(_0625_),
    .C(_0826_),
    .X(_1299_));
 sky130_fd_sc_hd__or2_2 _2868_ (.A(_1233_),
    .B(_1299_),
    .X(_1300_));
 sky130_fd_sc_hd__mux2_1 _2869_ (.A0(_1210_),
    .A1(\tms1x00.RAM[0][0] ),
    .S(_1300_),
    .X(_1301_));
 sky130_fd_sc_hd__clkbuf_1 _2870_ (.A(_1301_),
    .X(_0115_));
 sky130_fd_sc_hd__mux2_1 _2871_ (.A0(_1214_),
    .A1(\tms1x00.RAM[0][1] ),
    .S(_1300_),
    .X(_1302_));
 sky130_fd_sc_hd__clkbuf_1 _2872_ (.A(_1302_),
    .X(_0116_));
 sky130_fd_sc_hd__mux2_1 _2873_ (.A0(_1216_),
    .A1(\tms1x00.RAM[0][2] ),
    .S(_1300_),
    .X(_1303_));
 sky130_fd_sc_hd__clkbuf_1 _2874_ (.A(_1303_),
    .X(_0117_));
 sky130_fd_sc_hd__mux2_1 _2875_ (.A0(_1218_),
    .A1(\tms1x00.RAM[0][3] ),
    .S(_1300_),
    .X(_1304_));
 sky130_fd_sc_hd__clkbuf_1 _2876_ (.A(_1304_),
    .X(_0118_));
 sky130_fd_sc_hd__or3b_4 _2877_ (.A(_0826_),
    .B(_0617_),
    .C_N(_0625_),
    .X(_1305_));
 sky130_fd_sc_hd__or2_2 _2878_ (.A(_0822_),
    .B(_1305_),
    .X(_1306_));
 sky130_fd_sc_hd__mux2_1 _2879_ (.A0(_1210_),
    .A1(\tms1x00.RAM[98][0] ),
    .S(_1306_),
    .X(_1307_));
 sky130_fd_sc_hd__clkbuf_1 _2880_ (.A(_1307_),
    .X(_0119_));
 sky130_fd_sc_hd__mux2_1 _2881_ (.A0(_1214_),
    .A1(\tms1x00.RAM[98][1] ),
    .S(_1306_),
    .X(_1308_));
 sky130_fd_sc_hd__clkbuf_1 _2882_ (.A(_1308_),
    .X(_0120_));
 sky130_fd_sc_hd__mux2_1 _2883_ (.A0(_1216_),
    .A1(\tms1x00.RAM[98][2] ),
    .S(_1306_),
    .X(_1309_));
 sky130_fd_sc_hd__clkbuf_1 _2884_ (.A(_1309_),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _2885_ (.A0(_1218_),
    .A1(\tms1x00.RAM[98][3] ),
    .S(_1306_),
    .X(_1310_));
 sky130_fd_sc_hd__clkbuf_1 _2886_ (.A(_1310_),
    .X(_0122_));
 sky130_fd_sc_hd__or2_2 _2887_ (.A(_0822_),
    .B(_1182_),
    .X(_1311_));
 sky130_fd_sc_hd__mux2_1 _2888_ (.A0(_1210_),
    .A1(\tms1x00.RAM[97][0] ),
    .S(_1311_),
    .X(_1312_));
 sky130_fd_sc_hd__clkbuf_1 _2889_ (.A(_1312_),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _2890_ (.A0(_1214_),
    .A1(\tms1x00.RAM[97][1] ),
    .S(_1311_),
    .X(_1313_));
 sky130_fd_sc_hd__clkbuf_1 _2891_ (.A(_1313_),
    .X(_0124_));
 sky130_fd_sc_hd__mux2_1 _2892_ (.A0(_1216_),
    .A1(\tms1x00.RAM[97][2] ),
    .S(_1311_),
    .X(_1314_));
 sky130_fd_sc_hd__clkbuf_1 _2893_ (.A(_1314_),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_1 _2894_ (.A0(_1218_),
    .A1(\tms1x00.RAM[97][3] ),
    .S(_1311_),
    .X(_1315_));
 sky130_fd_sc_hd__clkbuf_1 _2895_ (.A(_1315_),
    .X(_0126_));
 sky130_fd_sc_hd__or2_2 _2896_ (.A(_0822_),
    .B(_1299_),
    .X(_1316_));
 sky130_fd_sc_hd__mux2_1 _2897_ (.A0(_1210_),
    .A1(\tms1x00.RAM[96][0] ),
    .S(_1316_),
    .X(_1317_));
 sky130_fd_sc_hd__clkbuf_1 _2898_ (.A(_1317_),
    .X(_0127_));
 sky130_fd_sc_hd__mux2_1 _2899_ (.A0(_1214_),
    .A1(\tms1x00.RAM[96][1] ),
    .S(_1316_),
    .X(_1318_));
 sky130_fd_sc_hd__clkbuf_1 _2900_ (.A(_1318_),
    .X(_0128_));
 sky130_fd_sc_hd__mux2_1 _2901_ (.A0(_1216_),
    .A1(\tms1x00.RAM[96][2] ),
    .S(_1316_),
    .X(_1319_));
 sky130_fd_sc_hd__clkbuf_1 _2902_ (.A(_1319_),
    .X(_0129_));
 sky130_fd_sc_hd__mux2_1 _2903_ (.A0(_1218_),
    .A1(\tms1x00.RAM[96][3] ),
    .S(_1316_),
    .X(_1320_));
 sky130_fd_sc_hd__clkbuf_1 _2904_ (.A(_1320_),
    .X(_0130_));
 sky130_fd_sc_hd__or2_2 _2905_ (.A(_0827_),
    .B(_1176_),
    .X(_1321_));
 sky130_fd_sc_hd__mux2_1 _2906_ (.A0(_1210_),
    .A1(\tms1x00.RAM[115][0] ),
    .S(_1321_),
    .X(_1322_));
 sky130_fd_sc_hd__clkbuf_1 _2907_ (.A(_1322_),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_1 _2908_ (.A0(_1214_),
    .A1(\tms1x00.RAM[115][1] ),
    .S(_1321_),
    .X(_1323_));
 sky130_fd_sc_hd__clkbuf_1 _2909_ (.A(_1323_),
    .X(_0132_));
 sky130_fd_sc_hd__mux2_1 _2910_ (.A0(_1216_),
    .A1(\tms1x00.RAM[115][2] ),
    .S(_1321_),
    .X(_1324_));
 sky130_fd_sc_hd__clkbuf_1 _2911_ (.A(_1324_),
    .X(_0133_));
 sky130_fd_sc_hd__mux2_1 _2912_ (.A0(_1218_),
    .A1(\tms1x00.RAM[115][3] ),
    .S(_1321_),
    .X(_1325_));
 sky130_fd_sc_hd__clkbuf_1 _2913_ (.A(_1325_),
    .X(_0134_));
 sky130_fd_sc_hd__clkbuf_4 _2914_ (.A(_0820_),
    .X(_1326_));
 sky130_fd_sc_hd__or2_2 _2915_ (.A(_1176_),
    .B(_1305_),
    .X(_1327_));
 sky130_fd_sc_hd__mux2_1 _2916_ (.A0(_1326_),
    .A1(\tms1x00.RAM[114][0] ),
    .S(_1327_),
    .X(_1328_));
 sky130_fd_sc_hd__clkbuf_1 _2917_ (.A(_1328_),
    .X(_0135_));
 sky130_fd_sc_hd__buf_2 _2918_ (.A(_0929_),
    .X(_1329_));
 sky130_fd_sc_hd__mux2_1 _2919_ (.A0(_1329_),
    .A1(\tms1x00.RAM[114][1] ),
    .S(_1327_),
    .X(_1330_));
 sky130_fd_sc_hd__clkbuf_1 _2920_ (.A(_1330_),
    .X(_0136_));
 sky130_fd_sc_hd__buf_2 _2921_ (.A(_1029_),
    .X(_1331_));
 sky130_fd_sc_hd__mux2_1 _2922_ (.A0(_1331_),
    .A1(\tms1x00.RAM[114][2] ),
    .S(_1327_),
    .X(_1332_));
 sky130_fd_sc_hd__clkbuf_1 _2923_ (.A(_1332_),
    .X(_0137_));
 sky130_fd_sc_hd__buf_2 _2924_ (.A(_1127_),
    .X(_1333_));
 sky130_fd_sc_hd__mux2_1 _2925_ (.A0(_1333_),
    .A1(\tms1x00.RAM[114][3] ),
    .S(_1327_),
    .X(_1334_));
 sky130_fd_sc_hd__clkbuf_1 _2926_ (.A(_1334_),
    .X(_0138_));
 sky130_fd_sc_hd__or2_2 _2927_ (.A(_1176_),
    .B(_1182_),
    .X(_1335_));
 sky130_fd_sc_hd__mux2_1 _2928_ (.A0(_1326_),
    .A1(\tms1x00.RAM[113][0] ),
    .S(_1335_),
    .X(_1336_));
 sky130_fd_sc_hd__clkbuf_1 _2929_ (.A(_1336_),
    .X(_0139_));
 sky130_fd_sc_hd__mux2_1 _2930_ (.A0(_1329_),
    .A1(\tms1x00.RAM[113][1] ),
    .S(_1335_),
    .X(_1337_));
 sky130_fd_sc_hd__clkbuf_1 _2931_ (.A(_1337_),
    .X(_0140_));
 sky130_fd_sc_hd__mux2_1 _2932_ (.A0(_1331_),
    .A1(\tms1x00.RAM[113][2] ),
    .S(_1335_),
    .X(_1338_));
 sky130_fd_sc_hd__clkbuf_1 _2933_ (.A(_1338_),
    .X(_0141_));
 sky130_fd_sc_hd__mux2_1 _2934_ (.A0(_1333_),
    .A1(\tms1x00.RAM[113][3] ),
    .S(_1335_),
    .X(_1339_));
 sky130_fd_sc_hd__clkbuf_1 _2935_ (.A(_1339_),
    .X(_0142_));
 sky130_fd_sc_hd__or2_2 _2936_ (.A(_1176_),
    .B(_1299_),
    .X(_1340_));
 sky130_fd_sc_hd__mux2_1 _2937_ (.A0(_1326_),
    .A1(\tms1x00.RAM[112][0] ),
    .S(_1340_),
    .X(_1341_));
 sky130_fd_sc_hd__clkbuf_1 _2938_ (.A(_1341_),
    .X(_0143_));
 sky130_fd_sc_hd__mux2_1 _2939_ (.A0(_1329_),
    .A1(\tms1x00.RAM[112][1] ),
    .S(_1340_),
    .X(_1342_));
 sky130_fd_sc_hd__clkbuf_1 _2940_ (.A(_1342_),
    .X(_0144_));
 sky130_fd_sc_hd__mux2_1 _2941_ (.A0(_1331_),
    .A1(\tms1x00.RAM[112][2] ),
    .S(_1340_),
    .X(_1343_));
 sky130_fd_sc_hd__clkbuf_1 _2942_ (.A(_1343_),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _2943_ (.A0(_1333_),
    .A1(\tms1x00.RAM[112][3] ),
    .S(_1340_),
    .X(_1344_));
 sky130_fd_sc_hd__clkbuf_1 _2944_ (.A(_1344_),
    .X(_0146_));
 sky130_fd_sc_hd__or2_2 _2945_ (.A(_0822_),
    .B(_1169_),
    .X(_1345_));
 sky130_fd_sc_hd__mux2_1 _2946_ (.A0(_1326_),
    .A1(\tms1x00.RAM[111][0] ),
    .S(_1345_),
    .X(_1346_));
 sky130_fd_sc_hd__clkbuf_1 _2947_ (.A(_1346_),
    .X(_0147_));
 sky130_fd_sc_hd__mux2_1 _2948_ (.A0(_1329_),
    .A1(\tms1x00.RAM[111][1] ),
    .S(_1345_),
    .X(_1347_));
 sky130_fd_sc_hd__clkbuf_1 _2949_ (.A(_1347_),
    .X(_0148_));
 sky130_fd_sc_hd__mux2_1 _2950_ (.A0(_1331_),
    .A1(\tms1x00.RAM[111][2] ),
    .S(_1345_),
    .X(_1348_));
 sky130_fd_sc_hd__clkbuf_1 _2951_ (.A(_1348_),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_1 _2952_ (.A0(_1333_),
    .A1(\tms1x00.RAM[111][3] ),
    .S(_1345_),
    .X(_1349_));
 sky130_fd_sc_hd__clkbuf_1 _2953_ (.A(_1349_),
    .X(_0150_));
 sky130_fd_sc_hd__or2_2 _2954_ (.A(_0822_),
    .B(_1199_),
    .X(_1350_));
 sky130_fd_sc_hd__mux2_1 _2955_ (.A0(_1326_),
    .A1(\tms1x00.RAM[110][0] ),
    .S(_1350_),
    .X(_1351_));
 sky130_fd_sc_hd__clkbuf_1 _2956_ (.A(_1351_),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _2957_ (.A0(_1329_),
    .A1(\tms1x00.RAM[110][1] ),
    .S(_1350_),
    .X(_1352_));
 sky130_fd_sc_hd__clkbuf_1 _2958_ (.A(_1352_),
    .X(_0152_));
 sky130_fd_sc_hd__mux2_1 _2959_ (.A0(_1331_),
    .A1(\tms1x00.RAM[110][2] ),
    .S(_1350_),
    .X(_1353_));
 sky130_fd_sc_hd__clkbuf_1 _2960_ (.A(_1353_),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _2961_ (.A0(_1333_),
    .A1(\tms1x00.RAM[110][3] ),
    .S(_1350_),
    .X(_1354_));
 sky130_fd_sc_hd__clkbuf_1 _2962_ (.A(_1354_),
    .X(_0154_));
 sky130_fd_sc_hd__nor2_2 _2963_ (.A(_1226_),
    .B(_1233_),
    .Y(_1355_));
 sky130_fd_sc_hd__mux2_1 _2964_ (.A0(\tms1x00.RAM[10][0] ),
    .A1(_1266_),
    .S(_1355_),
    .X(_1356_));
 sky130_fd_sc_hd__clkbuf_1 _2965_ (.A(_1356_),
    .X(_0155_));
 sky130_fd_sc_hd__mux2_1 _2966_ (.A0(\tms1x00.RAM[10][1] ),
    .A1(_1270_),
    .S(_1355_),
    .X(_1357_));
 sky130_fd_sc_hd__clkbuf_1 _2967_ (.A(_1357_),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _2968_ (.A0(\tms1x00.RAM[10][2] ),
    .A1(_1273_),
    .S(_1355_),
    .X(_1358_));
 sky130_fd_sc_hd__clkbuf_1 _2969_ (.A(_1358_),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_1 _2970_ (.A0(\tms1x00.RAM[10][3] ),
    .A1(_1276_),
    .S(_1355_),
    .X(_1359_));
 sky130_fd_sc_hd__clkbuf_1 _2971_ (.A(_1359_),
    .X(_0158_));
 sky130_fd_sc_hd__or2_2 _2972_ (.A(_0822_),
    .B(_1211_),
    .X(_1360_));
 sky130_fd_sc_hd__mux2_1 _2973_ (.A0(_1326_),
    .A1(\tms1x00.RAM[108][0] ),
    .S(_1360_),
    .X(_1361_));
 sky130_fd_sc_hd__clkbuf_1 _2974_ (.A(_1361_),
    .X(_0159_));
 sky130_fd_sc_hd__mux2_1 _2975_ (.A0(_1329_),
    .A1(\tms1x00.RAM[108][1] ),
    .S(_1360_),
    .X(_1362_));
 sky130_fd_sc_hd__clkbuf_1 _2976_ (.A(_1362_),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _2977_ (.A0(_1331_),
    .A1(\tms1x00.RAM[108][2] ),
    .S(_1360_),
    .X(_1363_));
 sky130_fd_sc_hd__clkbuf_1 _2978_ (.A(_1363_),
    .X(_0161_));
 sky130_fd_sc_hd__mux2_1 _2979_ (.A0(_1333_),
    .A1(\tms1x00.RAM[108][3] ),
    .S(_1360_),
    .X(_1364_));
 sky130_fd_sc_hd__clkbuf_1 _2980_ (.A(_1364_),
    .X(_0162_));
 sky130_fd_sc_hd__nor2_2 _2981_ (.A(_0823_),
    .B(_1147_),
    .Y(_1365_));
 sky130_fd_sc_hd__mux2_1 _2982_ (.A0(\tms1x00.RAM[107][0] ),
    .A1(_1266_),
    .S(_1365_),
    .X(_1366_));
 sky130_fd_sc_hd__clkbuf_1 _2983_ (.A(_1366_),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _2984_ (.A0(\tms1x00.RAM[107][1] ),
    .A1(_1270_),
    .S(_1365_),
    .X(_1367_));
 sky130_fd_sc_hd__clkbuf_1 _2985_ (.A(_1367_),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_1 _2986_ (.A0(\tms1x00.RAM[107][2] ),
    .A1(_1273_),
    .S(_1365_),
    .X(_1368_));
 sky130_fd_sc_hd__clkbuf_1 _2987_ (.A(_1368_),
    .X(_0165_));
 sky130_fd_sc_hd__mux2_1 _2988_ (.A0(\tms1x00.RAM[107][3] ),
    .A1(_1276_),
    .S(_1365_),
    .X(_1369_));
 sky130_fd_sc_hd__clkbuf_1 _2989_ (.A(_1369_),
    .X(_0166_));
 sky130_fd_sc_hd__nor2_2 _2990_ (.A(_0823_),
    .B(_1226_),
    .Y(_1370_));
 sky130_fd_sc_hd__mux2_1 _2991_ (.A0(\tms1x00.RAM[106][0] ),
    .A1(_1266_),
    .S(_1370_),
    .X(_1371_));
 sky130_fd_sc_hd__clkbuf_1 _2992_ (.A(_1371_),
    .X(_0167_));
 sky130_fd_sc_hd__mux2_1 _2993_ (.A0(\tms1x00.RAM[106][1] ),
    .A1(_1270_),
    .S(_1370_),
    .X(_1372_));
 sky130_fd_sc_hd__clkbuf_1 _2994_ (.A(_1372_),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _2995_ (.A0(\tms1x00.RAM[106][2] ),
    .A1(_1273_),
    .S(_1370_),
    .X(_1373_));
 sky130_fd_sc_hd__clkbuf_1 _2996_ (.A(_1373_),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_1 _2997_ (.A0(\tms1x00.RAM[106][3] ),
    .A1(_1276_),
    .S(_1370_),
    .X(_1374_));
 sky130_fd_sc_hd__clkbuf_1 _2998_ (.A(_1374_),
    .X(_0170_));
 sky130_fd_sc_hd__or2_2 _2999_ (.A(_1154_),
    .B(_1175_),
    .X(_1375_));
 sky130_fd_sc_hd__mux2_1 _3000_ (.A0(_1326_),
    .A1(\tms1x00.RAM[125][0] ),
    .S(_1375_),
    .X(_1376_));
 sky130_fd_sc_hd__clkbuf_1 _3001_ (.A(_1376_),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _3002_ (.A0(_1329_),
    .A1(\tms1x00.RAM[125][1] ),
    .S(_1375_),
    .X(_1377_));
 sky130_fd_sc_hd__clkbuf_1 _3003_ (.A(_1377_),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_1 _3004_ (.A0(_1331_),
    .A1(\tms1x00.RAM[125][2] ),
    .S(_1375_),
    .X(_1378_));
 sky130_fd_sc_hd__clkbuf_1 _3005_ (.A(_1378_),
    .X(_0173_));
 sky130_fd_sc_hd__mux2_1 _3006_ (.A0(_1333_),
    .A1(\tms1x00.RAM[125][3] ),
    .S(_1375_),
    .X(_1379_));
 sky130_fd_sc_hd__clkbuf_1 _3007_ (.A(_1379_),
    .X(_0174_));
 sky130_fd_sc_hd__or2_2 _3008_ (.A(_1176_),
    .B(_1211_),
    .X(_1380_));
 sky130_fd_sc_hd__mux2_1 _3009_ (.A0(_1326_),
    .A1(\tms1x00.RAM[124][0] ),
    .S(_1380_),
    .X(_1381_));
 sky130_fd_sc_hd__clkbuf_1 _3010_ (.A(_1381_),
    .X(_0175_));
 sky130_fd_sc_hd__mux2_1 _3011_ (.A0(_1329_),
    .A1(\tms1x00.RAM[124][1] ),
    .S(_1380_),
    .X(_1382_));
 sky130_fd_sc_hd__clkbuf_1 _3012_ (.A(_1382_),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _3013_ (.A0(_1331_),
    .A1(\tms1x00.RAM[124][2] ),
    .S(_1380_),
    .X(_1383_));
 sky130_fd_sc_hd__clkbuf_1 _3014_ (.A(_1383_),
    .X(_0177_));
 sky130_fd_sc_hd__mux2_1 _3015_ (.A0(_1333_),
    .A1(\tms1x00.RAM[124][3] ),
    .S(_1380_),
    .X(_1384_));
 sky130_fd_sc_hd__clkbuf_1 _3016_ (.A(_1384_),
    .X(_0178_));
 sky130_fd_sc_hd__or2_2 _3017_ (.A(_1147_),
    .B(_1175_),
    .X(_1385_));
 sky130_fd_sc_hd__mux2_1 _3018_ (.A0(_1326_),
    .A1(\tms1x00.RAM[123][0] ),
    .S(_1385_),
    .X(_1386_));
 sky130_fd_sc_hd__clkbuf_1 _3019_ (.A(_1386_),
    .X(_0179_));
 sky130_fd_sc_hd__mux2_1 _3020_ (.A0(_1329_),
    .A1(\tms1x00.RAM[123][1] ),
    .S(_1385_),
    .X(_1387_));
 sky130_fd_sc_hd__clkbuf_1 _3021_ (.A(_1387_),
    .X(_0180_));
 sky130_fd_sc_hd__mux2_1 _3022_ (.A0(_1331_),
    .A1(\tms1x00.RAM[123][2] ),
    .S(_1385_),
    .X(_1388_));
 sky130_fd_sc_hd__clkbuf_1 _3023_ (.A(_1388_),
    .X(_0181_));
 sky130_fd_sc_hd__mux2_1 _3024_ (.A0(_1333_),
    .A1(\tms1x00.RAM[123][3] ),
    .S(_1385_),
    .X(_1389_));
 sky130_fd_sc_hd__clkbuf_1 _3025_ (.A(_1389_),
    .X(_0182_));
 sky130_fd_sc_hd__or4bb_1 _3026_ (.A(\tms1x00.ram_addr_buff[0] ),
    .B(\tms1x00.ram_addr_buff[2] ),
    .C_N(\tms1x00.ram_addr_buff[3] ),
    .D_N(\tms1x00.ram_addr_buff[1] ),
    .X(_1390_));
 sky130_fd_sc_hd__or3_4 _3027_ (.A(_0825_),
    .B(_1175_),
    .C(_1390_),
    .X(_1391_));
 sky130_fd_sc_hd__mux2_1 _3028_ (.A0(_1326_),
    .A1(\tms1x00.RAM[122][0] ),
    .S(_1391_),
    .X(_1392_));
 sky130_fd_sc_hd__clkbuf_1 _3029_ (.A(_1392_),
    .X(_0183_));
 sky130_fd_sc_hd__mux2_1 _3030_ (.A0(_1329_),
    .A1(\tms1x00.RAM[122][1] ),
    .S(_1391_),
    .X(_1393_));
 sky130_fd_sc_hd__clkbuf_1 _3031_ (.A(_1393_),
    .X(_0184_));
 sky130_fd_sc_hd__mux2_1 _3032_ (.A0(_1331_),
    .A1(\tms1x00.RAM[122][2] ),
    .S(_1391_),
    .X(_1394_));
 sky130_fd_sc_hd__clkbuf_1 _3033_ (.A(_1394_),
    .X(_0185_));
 sky130_fd_sc_hd__mux2_1 _3034_ (.A0(_1333_),
    .A1(\tms1x00.RAM[122][3] ),
    .S(_1391_),
    .X(_1395_));
 sky130_fd_sc_hd__clkbuf_1 _3035_ (.A(_1395_),
    .X(_0186_));
 sky130_fd_sc_hd__clkbuf_4 _3036_ (.A(_0820_),
    .X(_1396_));
 sky130_fd_sc_hd__or4bb_1 _3037_ (.A(\tms1x00.ram_addr_buff[1] ),
    .B(\tms1x00.ram_addr_buff[2] ),
    .C_N(\tms1x00.ram_addr_buff[3] ),
    .D_N(\tms1x00.ram_addr_buff[0] ),
    .X(_1397_));
 sky130_fd_sc_hd__or3_4 _3038_ (.A(_0825_),
    .B(_1397_),
    .C(_1175_),
    .X(_1398_));
 sky130_fd_sc_hd__mux2_1 _3039_ (.A0(_1396_),
    .A1(\tms1x00.RAM[121][0] ),
    .S(_1398_),
    .X(_1399_));
 sky130_fd_sc_hd__clkbuf_1 _3040_ (.A(_1399_),
    .X(_0187_));
 sky130_fd_sc_hd__clkbuf_4 _3041_ (.A(_0929_),
    .X(_1400_));
 sky130_fd_sc_hd__mux2_1 _3042_ (.A0(_1400_),
    .A1(\tms1x00.RAM[121][1] ),
    .S(_1398_),
    .X(_1401_));
 sky130_fd_sc_hd__clkbuf_1 _3043_ (.A(_1401_),
    .X(_0188_));
 sky130_fd_sc_hd__clkbuf_4 _3044_ (.A(_1029_),
    .X(_1402_));
 sky130_fd_sc_hd__mux2_1 _3045_ (.A0(_1402_),
    .A1(\tms1x00.RAM[121][2] ),
    .S(_1398_),
    .X(_1403_));
 sky130_fd_sc_hd__clkbuf_1 _3046_ (.A(_1403_),
    .X(_0189_));
 sky130_fd_sc_hd__clkbuf_4 _3047_ (.A(_1127_),
    .X(_1404_));
 sky130_fd_sc_hd__mux2_1 _3048_ (.A0(_1404_),
    .A1(\tms1x00.RAM[121][3] ),
    .S(_1398_),
    .X(_1405_));
 sky130_fd_sc_hd__clkbuf_1 _3049_ (.A(_1405_),
    .X(_0190_));
 sky130_fd_sc_hd__or4b_1 _3050_ (.A(\tms1x00.ram_addr_buff[0] ),
    .B(\tms1x00.ram_addr_buff[1] ),
    .C(\tms1x00.ram_addr_buff[2] ),
    .D_N(\tms1x00.ram_addr_buff[3] ),
    .X(_1406_));
 sky130_fd_sc_hd__or3_4 _3051_ (.A(_0825_),
    .B(_1175_),
    .C(_1406_),
    .X(_1407_));
 sky130_fd_sc_hd__mux2_1 _3052_ (.A0(_1396_),
    .A1(\tms1x00.RAM[120][0] ),
    .S(_1407_),
    .X(_1408_));
 sky130_fd_sc_hd__clkbuf_1 _3053_ (.A(_1408_),
    .X(_0191_));
 sky130_fd_sc_hd__mux2_1 _3054_ (.A0(_1400_),
    .A1(\tms1x00.RAM[120][1] ),
    .S(_1407_),
    .X(_1409_));
 sky130_fd_sc_hd__clkbuf_1 _3055_ (.A(_1409_),
    .X(_0192_));
 sky130_fd_sc_hd__mux2_1 _3056_ (.A0(_1402_),
    .A1(\tms1x00.RAM[120][2] ),
    .S(_1407_),
    .X(_1410_));
 sky130_fd_sc_hd__clkbuf_1 _3057_ (.A(_1410_),
    .X(_0193_));
 sky130_fd_sc_hd__mux2_1 _3058_ (.A0(_1404_),
    .A1(\tms1x00.RAM[120][3] ),
    .S(_1407_),
    .X(_1411_));
 sky130_fd_sc_hd__clkbuf_1 _3059_ (.A(_1411_),
    .X(_0194_));
 sky130_fd_sc_hd__nor2_2 _3060_ (.A(_1147_),
    .B(_1233_),
    .Y(_1412_));
 sky130_fd_sc_hd__mux2_1 _3061_ (.A0(\tms1x00.RAM[11][0] ),
    .A1(_1266_),
    .S(_1412_),
    .X(_1413_));
 sky130_fd_sc_hd__clkbuf_1 _3062_ (.A(_1413_),
    .X(_0195_));
 sky130_fd_sc_hd__mux2_1 _3063_ (.A0(\tms1x00.RAM[11][1] ),
    .A1(_1270_),
    .S(_1412_),
    .X(_1414_));
 sky130_fd_sc_hd__clkbuf_1 _3064_ (.A(_1414_),
    .X(_0196_));
 sky130_fd_sc_hd__mux2_1 _3065_ (.A0(\tms1x00.RAM[11][2] ),
    .A1(_1273_),
    .S(_1412_),
    .X(_1415_));
 sky130_fd_sc_hd__clkbuf_1 _3066_ (.A(_1415_),
    .X(_0197_));
 sky130_fd_sc_hd__mux2_1 _3067_ (.A0(\tms1x00.RAM[11][3] ),
    .A1(_1276_),
    .S(_1412_),
    .X(_1416_));
 sky130_fd_sc_hd__clkbuf_1 _3068_ (.A(_1416_),
    .X(_0198_));
 sky130_fd_sc_hd__or2_2 _3069_ (.A(_1176_),
    .B(_1254_),
    .X(_1417_));
 sky130_fd_sc_hd__mux2_1 _3070_ (.A0(_1396_),
    .A1(\tms1x00.RAM[118][0] ),
    .S(_1417_),
    .X(_1418_));
 sky130_fd_sc_hd__clkbuf_1 _3071_ (.A(_1418_),
    .X(_0199_));
 sky130_fd_sc_hd__mux2_1 _3072_ (.A0(_1400_),
    .A1(\tms1x00.RAM[118][1] ),
    .S(_1417_),
    .X(_1419_));
 sky130_fd_sc_hd__clkbuf_1 _3073_ (.A(_1419_),
    .X(_0200_));
 sky130_fd_sc_hd__mux2_1 _3074_ (.A0(_1402_),
    .A1(\tms1x00.RAM[118][2] ),
    .S(_1417_),
    .X(_1420_));
 sky130_fd_sc_hd__clkbuf_1 _3075_ (.A(_1420_),
    .X(_0201_));
 sky130_fd_sc_hd__mux2_1 _3076_ (.A0(_1404_),
    .A1(\tms1x00.RAM[118][3] ),
    .S(_1417_),
    .X(_1421_));
 sky130_fd_sc_hd__clkbuf_1 _3077_ (.A(_1421_),
    .X(_0202_));
 sky130_fd_sc_hd__or2_2 _3078_ (.A(_1163_),
    .B(_1175_),
    .X(_1422_));
 sky130_fd_sc_hd__mux2_1 _3079_ (.A0(_1396_),
    .A1(\tms1x00.RAM[117][0] ),
    .S(_1422_),
    .X(_1423_));
 sky130_fd_sc_hd__clkbuf_1 _3080_ (.A(_1423_),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_1 _3081_ (.A0(_1400_),
    .A1(\tms1x00.RAM[117][1] ),
    .S(_1422_),
    .X(_1424_));
 sky130_fd_sc_hd__clkbuf_1 _3082_ (.A(_1424_),
    .X(_0204_));
 sky130_fd_sc_hd__mux2_1 _3083_ (.A0(_1402_),
    .A1(\tms1x00.RAM[117][2] ),
    .S(_1422_),
    .X(_1425_));
 sky130_fd_sc_hd__clkbuf_1 _3084_ (.A(_1425_),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _3085_ (.A0(_1404_),
    .A1(\tms1x00.RAM[117][3] ),
    .S(_1422_),
    .X(_1426_));
 sky130_fd_sc_hd__clkbuf_1 _3086_ (.A(_1426_),
    .X(_0206_));
 sky130_fd_sc_hd__or2_2 _3087_ (.A(_1176_),
    .B(_1293_),
    .X(_1427_));
 sky130_fd_sc_hd__mux2_1 _3088_ (.A0(_1396_),
    .A1(\tms1x00.RAM[116][0] ),
    .S(_1427_),
    .X(_1428_));
 sky130_fd_sc_hd__clkbuf_1 _3089_ (.A(_1428_),
    .X(_0207_));
 sky130_fd_sc_hd__mux2_1 _3090_ (.A0(_1400_),
    .A1(\tms1x00.RAM[116][1] ),
    .S(_1427_),
    .X(_1429_));
 sky130_fd_sc_hd__clkbuf_1 _3091_ (.A(_1429_),
    .X(_0208_));
 sky130_fd_sc_hd__mux2_1 _3092_ (.A0(_1402_),
    .A1(\tms1x00.RAM[116][2] ),
    .S(_1427_),
    .X(_1430_));
 sky130_fd_sc_hd__clkbuf_1 _3093_ (.A(_1430_),
    .X(_0209_));
 sky130_fd_sc_hd__mux2_1 _3094_ (.A0(_1404_),
    .A1(\tms1x00.RAM[116][3] ),
    .S(_1427_),
    .X(_1431_));
 sky130_fd_sc_hd__clkbuf_1 _3095_ (.A(_1431_),
    .X(_0210_));
 sky130_fd_sc_hd__or2_2 _3096_ (.A(_1176_),
    .B(_1199_),
    .X(_1432_));
 sky130_fd_sc_hd__mux2_1 _3097_ (.A0(_1396_),
    .A1(\tms1x00.RAM[126][0] ),
    .S(_1432_),
    .X(_1433_));
 sky130_fd_sc_hd__clkbuf_1 _3098_ (.A(_1433_),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_1 _3099_ (.A0(_1400_),
    .A1(\tms1x00.RAM[126][1] ),
    .S(_1432_),
    .X(_1434_));
 sky130_fd_sc_hd__clkbuf_1 _3100_ (.A(_1434_),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_1 _3101_ (.A0(_1402_),
    .A1(\tms1x00.RAM[126][2] ),
    .S(_1432_),
    .X(_1435_));
 sky130_fd_sc_hd__clkbuf_1 _3102_ (.A(_1435_),
    .X(_0213_));
 sky130_fd_sc_hd__mux2_1 _3103_ (.A0(_1404_),
    .A1(\tms1x00.RAM[126][3] ),
    .S(_1432_),
    .X(_1436_));
 sky130_fd_sc_hd__clkbuf_1 _3104_ (.A(_1436_),
    .X(_0214_));
 sky130_fd_sc_hd__or2_2 _3105_ (.A(_1182_),
    .B(_1233_),
    .X(_1437_));
 sky130_fd_sc_hd__mux2_1 _3106_ (.A0(_1396_),
    .A1(\tms1x00.RAM[1][0] ),
    .S(_1437_),
    .X(_1438_));
 sky130_fd_sc_hd__clkbuf_1 _3107_ (.A(_1438_),
    .X(_0215_));
 sky130_fd_sc_hd__mux2_1 _3108_ (.A0(_1400_),
    .A1(\tms1x00.RAM[1][1] ),
    .S(_1437_),
    .X(_1439_));
 sky130_fd_sc_hd__clkbuf_1 _3109_ (.A(_1439_),
    .X(_0216_));
 sky130_fd_sc_hd__mux2_1 _3110_ (.A0(_1402_),
    .A1(\tms1x00.RAM[1][2] ),
    .S(_1437_),
    .X(_1440_));
 sky130_fd_sc_hd__clkbuf_1 _3111_ (.A(_1440_),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _3112_ (.A0(_1404_),
    .A1(\tms1x00.RAM[1][3] ),
    .S(_1437_),
    .X(_1441_));
 sky130_fd_sc_hd__clkbuf_1 _3113_ (.A(_1441_),
    .X(_0218_));
 sky130_fd_sc_hd__buf_4 _3114_ (.A(_1188_),
    .X(_1442_));
 sky130_fd_sc_hd__nor2_2 _3115_ (.A(_1442_),
    .B(_1247_),
    .Y(_1443_));
 sky130_fd_sc_hd__mux2_1 _3116_ (.A0(\tms1x00.RAM[23][0] ),
    .A1(_1266_),
    .S(_1443_),
    .X(_1444_));
 sky130_fd_sc_hd__clkbuf_1 _3117_ (.A(_1444_),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _3118_ (.A0(\tms1x00.RAM[23][1] ),
    .A1(_1270_),
    .S(_1443_),
    .X(_1445_));
 sky130_fd_sc_hd__clkbuf_1 _3119_ (.A(_1445_),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _3120_ (.A0(\tms1x00.RAM[23][2] ),
    .A1(_1273_),
    .S(_1443_),
    .X(_1446_));
 sky130_fd_sc_hd__clkbuf_1 _3121_ (.A(_1446_),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _3122_ (.A0(\tms1x00.RAM[23][3] ),
    .A1(_1276_),
    .S(_1443_),
    .X(_1447_));
 sky130_fd_sc_hd__clkbuf_1 _3123_ (.A(_1447_),
    .X(_0222_));
 sky130_fd_sc_hd__or2_2 _3124_ (.A(_1442_),
    .B(_1254_),
    .X(_1448_));
 sky130_fd_sc_hd__mux2_1 _3125_ (.A0(_1396_),
    .A1(\tms1x00.RAM[22][0] ),
    .S(_1448_),
    .X(_1449_));
 sky130_fd_sc_hd__clkbuf_1 _3126_ (.A(_1449_),
    .X(_0223_));
 sky130_fd_sc_hd__mux2_1 _3127_ (.A0(_1400_),
    .A1(\tms1x00.RAM[22][1] ),
    .S(_1448_),
    .X(_1450_));
 sky130_fd_sc_hd__clkbuf_1 _3128_ (.A(_1450_),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_1 _3129_ (.A0(_1402_),
    .A1(\tms1x00.RAM[22][2] ),
    .S(_1448_),
    .X(_1451_));
 sky130_fd_sc_hd__clkbuf_1 _3130_ (.A(_1451_),
    .X(_0225_));
 sky130_fd_sc_hd__mux2_1 _3131_ (.A0(_1404_),
    .A1(\tms1x00.RAM[22][3] ),
    .S(_1448_),
    .X(_1452_));
 sky130_fd_sc_hd__clkbuf_1 _3132_ (.A(_1452_),
    .X(_0226_));
 sky130_fd_sc_hd__or2_2 _3133_ (.A(_1163_),
    .B(_1188_),
    .X(_1453_));
 sky130_fd_sc_hd__mux2_1 _3134_ (.A0(_1396_),
    .A1(\tms1x00.RAM[21][0] ),
    .S(_1453_),
    .X(_1454_));
 sky130_fd_sc_hd__clkbuf_1 _3135_ (.A(_1454_),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_1 _3136_ (.A0(_1400_),
    .A1(\tms1x00.RAM[21][1] ),
    .S(_1453_),
    .X(_1455_));
 sky130_fd_sc_hd__clkbuf_1 _3137_ (.A(_1455_),
    .X(_0228_));
 sky130_fd_sc_hd__mux2_1 _3138_ (.A0(_1402_),
    .A1(\tms1x00.RAM[21][2] ),
    .S(_1453_),
    .X(_1456_));
 sky130_fd_sc_hd__clkbuf_1 _3139_ (.A(_1456_),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_1 _3140_ (.A0(_1404_),
    .A1(\tms1x00.RAM[21][3] ),
    .S(_1453_),
    .X(_1457_));
 sky130_fd_sc_hd__clkbuf_1 _3141_ (.A(_1457_),
    .X(_0230_));
 sky130_fd_sc_hd__or2_2 _3142_ (.A(_1442_),
    .B(_1293_),
    .X(_1458_));
 sky130_fd_sc_hd__mux2_1 _3143_ (.A0(_1396_),
    .A1(\tms1x00.RAM[20][0] ),
    .S(_1458_),
    .X(_1459_));
 sky130_fd_sc_hd__clkbuf_1 _3144_ (.A(_1459_),
    .X(_0231_));
 sky130_fd_sc_hd__mux2_1 _3145_ (.A0(_1400_),
    .A1(\tms1x00.RAM[20][1] ),
    .S(_1458_),
    .X(_1460_));
 sky130_fd_sc_hd__clkbuf_1 _3146_ (.A(_1460_),
    .X(_0232_));
 sky130_fd_sc_hd__mux2_1 _3147_ (.A0(_1402_),
    .A1(\tms1x00.RAM[20][2] ),
    .S(_1458_),
    .X(_1461_));
 sky130_fd_sc_hd__clkbuf_1 _3148_ (.A(_1461_),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_1 _3149_ (.A0(_1404_),
    .A1(\tms1x00.RAM[20][3] ),
    .S(_1458_),
    .X(_1462_));
 sky130_fd_sc_hd__clkbuf_1 _3150_ (.A(_1462_),
    .X(_0234_));
 sky130_fd_sc_hd__buf_2 _3151_ (.A(_0820_),
    .X(_1463_));
 sky130_fd_sc_hd__or2_2 _3152_ (.A(_1442_),
    .B(_1211_),
    .X(_1464_));
 sky130_fd_sc_hd__mux2_1 _3153_ (.A0(_1463_),
    .A1(\tms1x00.RAM[28][0] ),
    .S(_1464_),
    .X(_1465_));
 sky130_fd_sc_hd__clkbuf_1 _3154_ (.A(_1465_),
    .X(_0235_));
 sky130_fd_sc_hd__clkbuf_4 _3155_ (.A(_0929_),
    .X(_1466_));
 sky130_fd_sc_hd__mux2_1 _3156_ (.A0(_1466_),
    .A1(\tms1x00.RAM[28][1] ),
    .S(_1464_),
    .X(_1467_));
 sky130_fd_sc_hd__clkbuf_1 _3157_ (.A(_1467_),
    .X(_0236_));
 sky130_fd_sc_hd__buf_2 _3158_ (.A(_1029_),
    .X(_1468_));
 sky130_fd_sc_hd__mux2_1 _3159_ (.A0(_1468_),
    .A1(\tms1x00.RAM[28][2] ),
    .S(_1464_),
    .X(_1469_));
 sky130_fd_sc_hd__clkbuf_1 _3160_ (.A(_1469_),
    .X(_0237_));
 sky130_fd_sc_hd__buf_2 _3161_ (.A(_1127_),
    .X(_1470_));
 sky130_fd_sc_hd__mux2_1 _3162_ (.A0(_1470_),
    .A1(\tms1x00.RAM[28][3] ),
    .S(_1464_),
    .X(_1471_));
 sky130_fd_sc_hd__clkbuf_1 _3163_ (.A(_1471_),
    .X(_0238_));
 sky130_fd_sc_hd__nor2_2 _3164_ (.A(_1147_),
    .B(_1442_),
    .Y(_1472_));
 sky130_fd_sc_hd__mux2_1 _3165_ (.A0(\tms1x00.RAM[27][0] ),
    .A1(_1266_),
    .S(_1472_),
    .X(_1473_));
 sky130_fd_sc_hd__clkbuf_1 _3166_ (.A(_1473_),
    .X(_0239_));
 sky130_fd_sc_hd__mux2_1 _3167_ (.A0(\tms1x00.RAM[27][1] ),
    .A1(_1270_),
    .S(_1472_),
    .X(_1474_));
 sky130_fd_sc_hd__clkbuf_1 _3168_ (.A(_1474_),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _3169_ (.A0(\tms1x00.RAM[27][2] ),
    .A1(_1273_),
    .S(_1472_),
    .X(_1475_));
 sky130_fd_sc_hd__clkbuf_1 _3170_ (.A(_1475_),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_1 _3171_ (.A0(\tms1x00.RAM[27][3] ),
    .A1(_1276_),
    .S(_1472_),
    .X(_1476_));
 sky130_fd_sc_hd__clkbuf_1 _3172_ (.A(_1476_),
    .X(_0242_));
 sky130_fd_sc_hd__nor2_2 _3173_ (.A(_1442_),
    .B(_1226_),
    .Y(_1477_));
 sky130_fd_sc_hd__mux2_1 _3174_ (.A0(\tms1x00.RAM[26][0] ),
    .A1(_1266_),
    .S(_1477_),
    .X(_1478_));
 sky130_fd_sc_hd__clkbuf_1 _3175_ (.A(_1478_),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _3176_ (.A0(\tms1x00.RAM[26][1] ),
    .A1(_1270_),
    .S(_1477_),
    .X(_1479_));
 sky130_fd_sc_hd__clkbuf_1 _3177_ (.A(_1479_),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _3178_ (.A0(\tms1x00.RAM[26][2] ),
    .A1(_1273_),
    .S(_1477_),
    .X(_1480_));
 sky130_fd_sc_hd__clkbuf_1 _3179_ (.A(_1480_),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _3180_ (.A0(\tms1x00.RAM[26][3] ),
    .A1(_1276_),
    .S(_1477_),
    .X(_1481_));
 sky130_fd_sc_hd__clkbuf_1 _3181_ (.A(_1481_),
    .X(_0246_));
 sky130_fd_sc_hd__nor2_2 _3182_ (.A(_1135_),
    .B(_1442_),
    .Y(_1482_));
 sky130_fd_sc_hd__mux2_1 _3183_ (.A0(\tms1x00.RAM[25][0] ),
    .A1(_1266_),
    .S(_1482_),
    .X(_1483_));
 sky130_fd_sc_hd__clkbuf_1 _3184_ (.A(_1483_),
    .X(_0247_));
 sky130_fd_sc_hd__mux2_1 _3185_ (.A0(\tms1x00.RAM[25][1] ),
    .A1(_1270_),
    .S(_1482_),
    .X(_1484_));
 sky130_fd_sc_hd__clkbuf_1 _3186_ (.A(_1484_),
    .X(_0248_));
 sky130_fd_sc_hd__mux2_1 _3187_ (.A0(\tms1x00.RAM[25][2] ),
    .A1(_1273_),
    .S(_1482_),
    .X(_1485_));
 sky130_fd_sc_hd__clkbuf_1 _3188_ (.A(_1485_),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _3189_ (.A0(\tms1x00.RAM[25][3] ),
    .A1(_1276_),
    .S(_1482_),
    .X(_1486_));
 sky130_fd_sc_hd__clkbuf_1 _3190_ (.A(_1486_),
    .X(_0250_));
 sky130_fd_sc_hd__clkbuf_4 _3191_ (.A(_1265_),
    .X(_1487_));
 sky130_fd_sc_hd__nor2_2 _3192_ (.A(_1442_),
    .B(_1235_),
    .Y(_1488_));
 sky130_fd_sc_hd__mux2_1 _3193_ (.A0(\tms1x00.RAM[24][0] ),
    .A1(_1487_),
    .S(_1488_),
    .X(_1489_));
 sky130_fd_sc_hd__clkbuf_1 _3194_ (.A(_1489_),
    .X(_0251_));
 sky130_fd_sc_hd__clkbuf_4 _3195_ (.A(_1269_),
    .X(_1490_));
 sky130_fd_sc_hd__mux2_1 _3196_ (.A0(\tms1x00.RAM[24][1] ),
    .A1(_1490_),
    .S(_1488_),
    .X(_1491_));
 sky130_fd_sc_hd__clkbuf_1 _3197_ (.A(_1491_),
    .X(_0252_));
 sky130_fd_sc_hd__clkbuf_4 _3198_ (.A(_1272_),
    .X(_1492_));
 sky130_fd_sc_hd__mux2_1 _3199_ (.A0(\tms1x00.RAM[24][2] ),
    .A1(_1492_),
    .S(_1488_),
    .X(_1493_));
 sky130_fd_sc_hd__clkbuf_1 _3200_ (.A(_1493_),
    .X(_0253_));
 sky130_fd_sc_hd__clkbuf_4 _3201_ (.A(_1275_),
    .X(_1494_));
 sky130_fd_sc_hd__mux2_1 _3202_ (.A0(\tms1x00.RAM[24][3] ),
    .A1(_1494_),
    .S(_1488_),
    .X(_1495_));
 sky130_fd_sc_hd__clkbuf_1 _3203_ (.A(_1495_),
    .X(_0254_));
 sky130_fd_sc_hd__or3b_2 _3204_ (.A(\tms1x00.ram_addr_buff[4] ),
    .B(\tms1x00.ram_addr_buff[6] ),
    .C_N(\tms1x00.ram_addr_buff[5] ),
    .X(_1496_));
 sky130_fd_sc_hd__buf_4 _3205_ (.A(_1496_),
    .X(_1497_));
 sky130_fd_sc_hd__or2_2 _3206_ (.A(_1299_),
    .B(_1497_),
    .X(_1498_));
 sky130_fd_sc_hd__mux2_1 _3207_ (.A0(_1463_),
    .A1(\tms1x00.RAM[32][0] ),
    .S(_1498_),
    .X(_1499_));
 sky130_fd_sc_hd__clkbuf_1 _3208_ (.A(_1499_),
    .X(_0255_));
 sky130_fd_sc_hd__mux2_1 _3209_ (.A0(_1466_),
    .A1(\tms1x00.RAM[32][1] ),
    .S(_1498_),
    .X(_1500_));
 sky130_fd_sc_hd__clkbuf_1 _3210_ (.A(_1500_),
    .X(_0256_));
 sky130_fd_sc_hd__mux2_1 _3211_ (.A0(_1468_),
    .A1(\tms1x00.RAM[32][2] ),
    .S(_1498_),
    .X(_1501_));
 sky130_fd_sc_hd__clkbuf_1 _3212_ (.A(_1501_),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _3213_ (.A0(_1470_),
    .A1(\tms1x00.RAM[32][3] ),
    .S(_1498_),
    .X(_1502_));
 sky130_fd_sc_hd__clkbuf_1 _3214_ (.A(_1502_),
    .X(_0258_));
 sky130_fd_sc_hd__or2_2 _3215_ (.A(_1169_),
    .B(_1188_),
    .X(_1503_));
 sky130_fd_sc_hd__mux2_1 _3216_ (.A0(_1463_),
    .A1(\tms1x00.RAM[31][0] ),
    .S(_1503_),
    .X(_1504_));
 sky130_fd_sc_hd__clkbuf_1 _3217_ (.A(_1504_),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _3218_ (.A0(_1466_),
    .A1(\tms1x00.RAM[31][1] ),
    .S(_1503_),
    .X(_1505_));
 sky130_fd_sc_hd__clkbuf_1 _3219_ (.A(_1505_),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_1 _3220_ (.A0(_1468_),
    .A1(\tms1x00.RAM[31][2] ),
    .S(_1503_),
    .X(_1506_));
 sky130_fd_sc_hd__clkbuf_1 _3221_ (.A(_1506_),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _3222_ (.A0(_1470_),
    .A1(\tms1x00.RAM[31][3] ),
    .S(_1503_),
    .X(_1507_));
 sky130_fd_sc_hd__clkbuf_1 _3223_ (.A(_1507_),
    .X(_0262_));
 sky130_fd_sc_hd__or2_2 _3224_ (.A(_1442_),
    .B(_1199_),
    .X(_1508_));
 sky130_fd_sc_hd__mux2_1 _3225_ (.A0(_1463_),
    .A1(\tms1x00.RAM[30][0] ),
    .S(_1508_),
    .X(_1509_));
 sky130_fd_sc_hd__clkbuf_1 _3226_ (.A(_1509_),
    .X(_0263_));
 sky130_fd_sc_hd__mux2_1 _3227_ (.A0(_1466_),
    .A1(\tms1x00.RAM[30][1] ),
    .S(_1508_),
    .X(_1510_));
 sky130_fd_sc_hd__clkbuf_1 _3228_ (.A(_1510_),
    .X(_0264_));
 sky130_fd_sc_hd__mux2_1 _3229_ (.A0(_1468_),
    .A1(\tms1x00.RAM[30][2] ),
    .S(_1508_),
    .X(_1511_));
 sky130_fd_sc_hd__clkbuf_1 _3230_ (.A(_1511_),
    .X(_0265_));
 sky130_fd_sc_hd__mux2_1 _3231_ (.A0(_1470_),
    .A1(\tms1x00.RAM[30][3] ),
    .S(_1508_),
    .X(_1512_));
 sky130_fd_sc_hd__clkbuf_1 _3232_ (.A(_1512_),
    .X(_0266_));
 sky130_fd_sc_hd__or2_2 _3233_ (.A(_1233_),
    .B(_1305_),
    .X(_1513_));
 sky130_fd_sc_hd__mux2_1 _3234_ (.A0(_1463_),
    .A1(\tms1x00.RAM[2][0] ),
    .S(_1513_),
    .X(_1514_));
 sky130_fd_sc_hd__clkbuf_1 _3235_ (.A(_1514_),
    .X(_0267_));
 sky130_fd_sc_hd__mux2_1 _3236_ (.A0(_1466_),
    .A1(\tms1x00.RAM[2][1] ),
    .S(_1513_),
    .X(_1515_));
 sky130_fd_sc_hd__clkbuf_1 _3237_ (.A(_1515_),
    .X(_0268_));
 sky130_fd_sc_hd__mux2_1 _3238_ (.A0(_1468_),
    .A1(\tms1x00.RAM[2][2] ),
    .S(_1513_),
    .X(_1516_));
 sky130_fd_sc_hd__clkbuf_1 _3239_ (.A(_1516_),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _3240_ (.A0(_1470_),
    .A1(\tms1x00.RAM[2][3] ),
    .S(_1513_),
    .X(_1517_));
 sky130_fd_sc_hd__clkbuf_1 _3241_ (.A(_1517_),
    .X(_0270_));
 sky130_fd_sc_hd__or2_2 _3242_ (.A(_1293_),
    .B(_1497_),
    .X(_1518_));
 sky130_fd_sc_hd__mux2_1 _3243_ (.A0(_1463_),
    .A1(\tms1x00.RAM[36][0] ),
    .S(_1518_),
    .X(_1519_));
 sky130_fd_sc_hd__clkbuf_1 _3244_ (.A(_1519_),
    .X(_0271_));
 sky130_fd_sc_hd__mux2_1 _3245_ (.A0(_1466_),
    .A1(\tms1x00.RAM[36][1] ),
    .S(_1518_),
    .X(_1520_));
 sky130_fd_sc_hd__clkbuf_1 _3246_ (.A(_1520_),
    .X(_0272_));
 sky130_fd_sc_hd__mux2_1 _3247_ (.A0(_1468_),
    .A1(\tms1x00.RAM[36][2] ),
    .S(_1518_),
    .X(_1521_));
 sky130_fd_sc_hd__clkbuf_1 _3248_ (.A(_1521_),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _3249_ (.A0(_1470_),
    .A1(\tms1x00.RAM[36][3] ),
    .S(_1518_),
    .X(_1522_));
 sky130_fd_sc_hd__clkbuf_1 _3250_ (.A(_1522_),
    .X(_0274_));
 sky130_fd_sc_hd__or2_2 _3251_ (.A(_0827_),
    .B(_1497_),
    .X(_1523_));
 sky130_fd_sc_hd__mux2_1 _3252_ (.A0(_1463_),
    .A1(\tms1x00.RAM[35][0] ),
    .S(_1523_),
    .X(_1524_));
 sky130_fd_sc_hd__clkbuf_1 _3253_ (.A(_1524_),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_1 _3254_ (.A0(_1466_),
    .A1(\tms1x00.RAM[35][1] ),
    .S(_1523_),
    .X(_1525_));
 sky130_fd_sc_hd__clkbuf_1 _3255_ (.A(_1525_),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_1 _3256_ (.A0(_1468_),
    .A1(\tms1x00.RAM[35][2] ),
    .S(_1523_),
    .X(_1526_));
 sky130_fd_sc_hd__clkbuf_1 _3257_ (.A(_1526_),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_1 _3258_ (.A0(_1470_),
    .A1(\tms1x00.RAM[35][3] ),
    .S(_1523_),
    .X(_1527_));
 sky130_fd_sc_hd__clkbuf_1 _3259_ (.A(_1527_),
    .X(_0278_));
 sky130_fd_sc_hd__or2_2 _3260_ (.A(_1305_),
    .B(_1497_),
    .X(_1528_));
 sky130_fd_sc_hd__mux2_1 _3261_ (.A0(_1463_),
    .A1(\tms1x00.RAM[34][0] ),
    .S(_1528_),
    .X(_1529_));
 sky130_fd_sc_hd__clkbuf_1 _3262_ (.A(_1529_),
    .X(_0279_));
 sky130_fd_sc_hd__mux2_1 _3263_ (.A0(_1466_),
    .A1(\tms1x00.RAM[34][1] ),
    .S(_1528_),
    .X(_1530_));
 sky130_fd_sc_hd__clkbuf_1 _3264_ (.A(_1530_),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_1 _3265_ (.A0(_1468_),
    .A1(\tms1x00.RAM[34][2] ),
    .S(_1528_),
    .X(_1531_));
 sky130_fd_sc_hd__clkbuf_1 _3266_ (.A(_1531_),
    .X(_0281_));
 sky130_fd_sc_hd__mux2_1 _3267_ (.A0(_1470_),
    .A1(\tms1x00.RAM[34][3] ),
    .S(_1528_),
    .X(_1532_));
 sky130_fd_sc_hd__clkbuf_1 _3268_ (.A(_1532_),
    .X(_0282_));
 sky130_fd_sc_hd__or2_2 _3269_ (.A(_1182_),
    .B(_1497_),
    .X(_1533_));
 sky130_fd_sc_hd__mux2_1 _3270_ (.A0(_1463_),
    .A1(\tms1x00.RAM[33][0] ),
    .S(_1533_),
    .X(_1534_));
 sky130_fd_sc_hd__clkbuf_1 _3271_ (.A(_1534_),
    .X(_0283_));
 sky130_fd_sc_hd__mux2_1 _3272_ (.A0(_1466_),
    .A1(\tms1x00.RAM[33][1] ),
    .S(_1533_),
    .X(_1535_));
 sky130_fd_sc_hd__clkbuf_1 _3273_ (.A(_1535_),
    .X(_0284_));
 sky130_fd_sc_hd__mux2_1 _3274_ (.A0(_1468_),
    .A1(\tms1x00.RAM[33][2] ),
    .S(_1533_),
    .X(_1536_));
 sky130_fd_sc_hd__clkbuf_1 _3275_ (.A(_1536_),
    .X(_0285_));
 sky130_fd_sc_hd__mux2_1 _3276_ (.A0(_1470_),
    .A1(\tms1x00.RAM[33][3] ),
    .S(_1533_),
    .X(_1537_));
 sky130_fd_sc_hd__clkbuf_1 _3277_ (.A(_1537_),
    .X(_0286_));
 sky130_fd_sc_hd__nor2_2 _3278_ (.A(_1135_),
    .B(_1497_),
    .Y(_1538_));
 sky130_fd_sc_hd__mux2_1 _3279_ (.A0(\tms1x00.RAM[41][0] ),
    .A1(_1487_),
    .S(_1538_),
    .X(_1539_));
 sky130_fd_sc_hd__clkbuf_1 _3280_ (.A(_1539_),
    .X(_0287_));
 sky130_fd_sc_hd__mux2_1 _3281_ (.A0(\tms1x00.RAM[41][1] ),
    .A1(_1490_),
    .S(_1538_),
    .X(_1540_));
 sky130_fd_sc_hd__clkbuf_1 _3282_ (.A(_1540_),
    .X(_0288_));
 sky130_fd_sc_hd__mux2_1 _3283_ (.A0(\tms1x00.RAM[41][2] ),
    .A1(_1492_),
    .S(_1538_),
    .X(_1541_));
 sky130_fd_sc_hd__clkbuf_1 _3284_ (.A(_1541_),
    .X(_0289_));
 sky130_fd_sc_hd__mux2_1 _3285_ (.A0(\tms1x00.RAM[41][3] ),
    .A1(_1494_),
    .S(_1538_),
    .X(_1542_));
 sky130_fd_sc_hd__clkbuf_1 _3286_ (.A(_1542_),
    .X(_0290_));
 sky130_fd_sc_hd__nor2_2 _3287_ (.A(_1235_),
    .B(_1497_),
    .Y(_1543_));
 sky130_fd_sc_hd__mux2_1 _3288_ (.A0(\tms1x00.RAM[40][0] ),
    .A1(_1487_),
    .S(_1543_),
    .X(_1544_));
 sky130_fd_sc_hd__clkbuf_1 _3289_ (.A(_1544_),
    .X(_0291_));
 sky130_fd_sc_hd__mux2_1 _3290_ (.A0(\tms1x00.RAM[40][1] ),
    .A1(_1490_),
    .S(_1543_),
    .X(_1545_));
 sky130_fd_sc_hd__clkbuf_1 _3291_ (.A(_1545_),
    .X(_0292_));
 sky130_fd_sc_hd__mux2_1 _3292_ (.A0(\tms1x00.RAM[40][2] ),
    .A1(_1492_),
    .S(_1543_),
    .X(_1546_));
 sky130_fd_sc_hd__clkbuf_1 _3293_ (.A(_1546_),
    .X(_0293_));
 sky130_fd_sc_hd__mux2_1 _3294_ (.A0(\tms1x00.RAM[40][3] ),
    .A1(_1494_),
    .S(_1543_),
    .X(_1547_));
 sky130_fd_sc_hd__clkbuf_1 _3295_ (.A(_1547_),
    .X(_0294_));
 sky130_fd_sc_hd__or2_2 _3296_ (.A(_0827_),
    .B(_1232_),
    .X(_1548_));
 sky130_fd_sc_hd__mux2_1 _3297_ (.A0(_1463_),
    .A1(\tms1x00.RAM[3][0] ),
    .S(_1548_),
    .X(_1549_));
 sky130_fd_sc_hd__clkbuf_1 _3298_ (.A(_1549_),
    .X(_0295_));
 sky130_fd_sc_hd__mux2_1 _3299_ (.A0(_1466_),
    .A1(\tms1x00.RAM[3][1] ),
    .S(_1548_),
    .X(_1550_));
 sky130_fd_sc_hd__clkbuf_1 _3300_ (.A(_1550_),
    .X(_0296_));
 sky130_fd_sc_hd__mux2_1 _3301_ (.A0(_1468_),
    .A1(\tms1x00.RAM[3][2] ),
    .S(_1548_),
    .X(_1551_));
 sky130_fd_sc_hd__clkbuf_1 _3302_ (.A(_1551_),
    .X(_0297_));
 sky130_fd_sc_hd__mux2_1 _3303_ (.A0(_1470_),
    .A1(\tms1x00.RAM[3][3] ),
    .S(_1548_),
    .X(_1552_));
 sky130_fd_sc_hd__clkbuf_1 _3304_ (.A(_1552_),
    .X(_0298_));
 sky130_fd_sc_hd__buf_2 _3305_ (.A(_0820_),
    .X(_1553_));
 sky130_fd_sc_hd__or2_2 _3306_ (.A(_1254_),
    .B(_1496_),
    .X(_1554_));
 sky130_fd_sc_hd__mux2_1 _3307_ (.A0(_1553_),
    .A1(\tms1x00.RAM[38][0] ),
    .S(_1554_),
    .X(_1555_));
 sky130_fd_sc_hd__clkbuf_1 _3308_ (.A(_1555_),
    .X(_0299_));
 sky130_fd_sc_hd__clkbuf_4 _3309_ (.A(_0929_),
    .X(_1556_));
 sky130_fd_sc_hd__mux2_1 _3310_ (.A0(_1556_),
    .A1(\tms1x00.RAM[38][1] ),
    .S(_1554_),
    .X(_1557_));
 sky130_fd_sc_hd__clkbuf_1 _3311_ (.A(_1557_),
    .X(_0300_));
 sky130_fd_sc_hd__buf_2 _3312_ (.A(_1029_),
    .X(_1558_));
 sky130_fd_sc_hd__mux2_1 _3313_ (.A0(_1558_),
    .A1(\tms1x00.RAM[38][2] ),
    .S(_1554_),
    .X(_1559_));
 sky130_fd_sc_hd__clkbuf_1 _3314_ (.A(_1559_),
    .X(_0301_));
 sky130_fd_sc_hd__buf_2 _3315_ (.A(_1127_),
    .X(_1560_));
 sky130_fd_sc_hd__mux2_1 _3316_ (.A0(_1560_),
    .A1(\tms1x00.RAM[38][3] ),
    .S(_1554_),
    .X(_1561_));
 sky130_fd_sc_hd__clkbuf_1 _3317_ (.A(_1561_),
    .X(_0302_));
 sky130_fd_sc_hd__or2_2 _3318_ (.A(_1163_),
    .B(_1496_),
    .X(_1562_));
 sky130_fd_sc_hd__mux2_1 _3319_ (.A0(_1553_),
    .A1(\tms1x00.RAM[37][0] ),
    .S(_1562_),
    .X(_1563_));
 sky130_fd_sc_hd__clkbuf_1 _3320_ (.A(_1563_),
    .X(_0303_));
 sky130_fd_sc_hd__mux2_1 _3321_ (.A0(_1556_),
    .A1(\tms1x00.RAM[37][1] ),
    .S(_1562_),
    .X(_1564_));
 sky130_fd_sc_hd__clkbuf_1 _3322_ (.A(_1564_),
    .X(_0304_));
 sky130_fd_sc_hd__mux2_1 _3323_ (.A0(_1558_),
    .A1(\tms1x00.RAM[37][2] ),
    .S(_1562_),
    .X(_1565_));
 sky130_fd_sc_hd__clkbuf_1 _3324_ (.A(_1565_),
    .X(_0305_));
 sky130_fd_sc_hd__mux2_1 _3325_ (.A0(_1560_),
    .A1(\tms1x00.RAM[37][3] ),
    .S(_1562_),
    .X(_1566_));
 sky130_fd_sc_hd__clkbuf_1 _3326_ (.A(_1566_),
    .X(_0306_));
 sky130_fd_sc_hd__or2_2 _3327_ (.A(_1154_),
    .B(_1496_),
    .X(_1567_));
 sky130_fd_sc_hd__mux2_1 _3328_ (.A0(_1553_),
    .A1(\tms1x00.RAM[45][0] ),
    .S(_1567_),
    .X(_1568_));
 sky130_fd_sc_hd__clkbuf_1 _3329_ (.A(_1568_),
    .X(_0307_));
 sky130_fd_sc_hd__mux2_1 _3330_ (.A0(_1556_),
    .A1(\tms1x00.RAM[45][1] ),
    .S(_1567_),
    .X(_1569_));
 sky130_fd_sc_hd__clkbuf_1 _3331_ (.A(_1569_),
    .X(_0308_));
 sky130_fd_sc_hd__mux2_1 _3332_ (.A0(_1558_),
    .A1(\tms1x00.RAM[45][2] ),
    .S(_1567_),
    .X(_1570_));
 sky130_fd_sc_hd__clkbuf_1 _3333_ (.A(_1570_),
    .X(_0309_));
 sky130_fd_sc_hd__mux2_1 _3334_ (.A0(_1560_),
    .A1(\tms1x00.RAM[45][3] ),
    .S(_1567_),
    .X(_1571_));
 sky130_fd_sc_hd__clkbuf_1 _3335_ (.A(_1571_),
    .X(_0310_));
 sky130_fd_sc_hd__or2_2 _3336_ (.A(_1211_),
    .B(_1496_),
    .X(_1572_));
 sky130_fd_sc_hd__mux2_1 _3337_ (.A0(_1553_),
    .A1(\tms1x00.RAM[44][0] ),
    .S(_1572_),
    .X(_1573_));
 sky130_fd_sc_hd__clkbuf_1 _3338_ (.A(_1573_),
    .X(_0311_));
 sky130_fd_sc_hd__mux2_1 _3339_ (.A0(_1556_),
    .A1(\tms1x00.RAM[44][1] ),
    .S(_1572_),
    .X(_1574_));
 sky130_fd_sc_hd__clkbuf_1 _3340_ (.A(_1574_),
    .X(_0312_));
 sky130_fd_sc_hd__mux2_1 _3341_ (.A0(_1558_),
    .A1(\tms1x00.RAM[44][2] ),
    .S(_1572_),
    .X(_1575_));
 sky130_fd_sc_hd__clkbuf_1 _3342_ (.A(_1575_),
    .X(_0313_));
 sky130_fd_sc_hd__mux2_1 _3343_ (.A0(_1560_),
    .A1(\tms1x00.RAM[44][3] ),
    .S(_1572_),
    .X(_1576_));
 sky130_fd_sc_hd__clkbuf_1 _3344_ (.A(_1576_),
    .X(_0314_));
 sky130_fd_sc_hd__nor2_2 _3345_ (.A(_1147_),
    .B(_1497_),
    .Y(_1577_));
 sky130_fd_sc_hd__mux2_1 _3346_ (.A0(\tms1x00.RAM[43][0] ),
    .A1(_1487_),
    .S(_1577_),
    .X(_1578_));
 sky130_fd_sc_hd__clkbuf_1 _3347_ (.A(_1578_),
    .X(_0315_));
 sky130_fd_sc_hd__mux2_1 _3348_ (.A0(\tms1x00.RAM[43][1] ),
    .A1(_1490_),
    .S(_1577_),
    .X(_1579_));
 sky130_fd_sc_hd__clkbuf_1 _3349_ (.A(_1579_),
    .X(_0316_));
 sky130_fd_sc_hd__mux2_1 _3350_ (.A0(\tms1x00.RAM[43][2] ),
    .A1(_1492_),
    .S(_1577_),
    .X(_1580_));
 sky130_fd_sc_hd__clkbuf_1 _3351_ (.A(_1580_),
    .X(_0317_));
 sky130_fd_sc_hd__mux2_1 _3352_ (.A0(\tms1x00.RAM[43][3] ),
    .A1(_1494_),
    .S(_1577_),
    .X(_1581_));
 sky130_fd_sc_hd__clkbuf_1 _3353_ (.A(_1581_),
    .X(_0318_));
 sky130_fd_sc_hd__nor2_2 _3354_ (.A(_1226_),
    .B(_1497_),
    .Y(_1582_));
 sky130_fd_sc_hd__mux2_1 _3355_ (.A0(\tms1x00.RAM[42][0] ),
    .A1(_1487_),
    .S(_1582_),
    .X(_1583_));
 sky130_fd_sc_hd__clkbuf_1 _3356_ (.A(_1583_),
    .X(_0319_));
 sky130_fd_sc_hd__mux2_1 _3357_ (.A0(\tms1x00.RAM[42][1] ),
    .A1(_1490_),
    .S(_1582_),
    .X(_1584_));
 sky130_fd_sc_hd__clkbuf_1 _3358_ (.A(_1584_),
    .X(_0320_));
 sky130_fd_sc_hd__mux2_1 _3359_ (.A0(\tms1x00.RAM[42][2] ),
    .A1(_1492_),
    .S(_1582_),
    .X(_1585_));
 sky130_fd_sc_hd__clkbuf_1 _3360_ (.A(_1585_),
    .X(_0321_));
 sky130_fd_sc_hd__mux2_1 _3361_ (.A0(\tms1x00.RAM[42][3] ),
    .A1(_1494_),
    .S(_1582_),
    .X(_1586_));
 sky130_fd_sc_hd__clkbuf_1 _3362_ (.A(_1586_),
    .X(_0322_));
 sky130_fd_sc_hd__or2_2 _3363_ (.A(_1145_),
    .B(_1305_),
    .X(_1587_));
 sky130_fd_sc_hd__mux2_1 _3364_ (.A0(_1553_),
    .A1(\tms1x00.RAM[50][0] ),
    .S(_1587_),
    .X(_1588_));
 sky130_fd_sc_hd__clkbuf_1 _3365_ (.A(_1588_),
    .X(_0323_));
 sky130_fd_sc_hd__mux2_1 _3366_ (.A0(_1556_),
    .A1(\tms1x00.RAM[50][1] ),
    .S(_1587_),
    .X(_1589_));
 sky130_fd_sc_hd__clkbuf_1 _3367_ (.A(_1589_),
    .X(_0324_));
 sky130_fd_sc_hd__mux2_1 _3368_ (.A0(_1558_),
    .A1(\tms1x00.RAM[50][2] ),
    .S(_1587_),
    .X(_1590_));
 sky130_fd_sc_hd__clkbuf_1 _3369_ (.A(_1590_),
    .X(_0325_));
 sky130_fd_sc_hd__mux2_1 _3370_ (.A0(_1560_),
    .A1(\tms1x00.RAM[50][3] ),
    .S(_1587_),
    .X(_1591_));
 sky130_fd_sc_hd__clkbuf_1 _3371_ (.A(_1591_),
    .X(_0326_));
 sky130_fd_sc_hd__or2_2 _3372_ (.A(_1233_),
    .B(_1293_),
    .X(_1592_));
 sky130_fd_sc_hd__mux2_1 _3373_ (.A0(_1553_),
    .A1(\tms1x00.RAM[4][0] ),
    .S(_1592_),
    .X(_1593_));
 sky130_fd_sc_hd__clkbuf_1 _3374_ (.A(_1593_),
    .X(_0327_));
 sky130_fd_sc_hd__mux2_1 _3375_ (.A0(_1556_),
    .A1(\tms1x00.RAM[4][1] ),
    .S(_1592_),
    .X(_1594_));
 sky130_fd_sc_hd__clkbuf_1 _3376_ (.A(_1594_),
    .X(_0328_));
 sky130_fd_sc_hd__mux2_1 _3377_ (.A0(_1558_),
    .A1(\tms1x00.RAM[4][2] ),
    .S(_1592_),
    .X(_1595_));
 sky130_fd_sc_hd__clkbuf_1 _3378_ (.A(_1595_),
    .X(_0329_));
 sky130_fd_sc_hd__mux2_1 _3379_ (.A0(_1560_),
    .A1(\tms1x00.RAM[4][3] ),
    .S(_1592_),
    .X(_1596_));
 sky130_fd_sc_hd__clkbuf_1 _3380_ (.A(_1596_),
    .X(_0330_));
 sky130_fd_sc_hd__or2_2 _3381_ (.A(_1145_),
    .B(_1299_),
    .X(_1597_));
 sky130_fd_sc_hd__mux2_1 _3382_ (.A0(_1553_),
    .A1(\tms1x00.RAM[48][0] ),
    .S(_1597_),
    .X(_1598_));
 sky130_fd_sc_hd__clkbuf_1 _3383_ (.A(_1598_),
    .X(_0331_));
 sky130_fd_sc_hd__mux2_1 _3384_ (.A0(_1556_),
    .A1(\tms1x00.RAM[48][1] ),
    .S(_1597_),
    .X(_1599_));
 sky130_fd_sc_hd__clkbuf_1 _3385_ (.A(_1599_),
    .X(_0332_));
 sky130_fd_sc_hd__mux2_1 _3386_ (.A0(_1558_),
    .A1(\tms1x00.RAM[48][2] ),
    .S(_1597_),
    .X(_1600_));
 sky130_fd_sc_hd__clkbuf_1 _3387_ (.A(_1600_),
    .X(_0333_));
 sky130_fd_sc_hd__mux2_1 _3388_ (.A0(_1560_),
    .A1(\tms1x00.RAM[48][3] ),
    .S(_1597_),
    .X(_1601_));
 sky130_fd_sc_hd__clkbuf_1 _3389_ (.A(_1601_),
    .X(_0334_));
 sky130_fd_sc_hd__or2_2 _3390_ (.A(_1169_),
    .B(_1496_),
    .X(_1602_));
 sky130_fd_sc_hd__mux2_1 _3391_ (.A0(_1553_),
    .A1(\tms1x00.RAM[47][0] ),
    .S(_1602_),
    .X(_1603_));
 sky130_fd_sc_hd__clkbuf_1 _3392_ (.A(_1603_),
    .X(_0335_));
 sky130_fd_sc_hd__mux2_1 _3393_ (.A0(_1556_),
    .A1(\tms1x00.RAM[47][1] ),
    .S(_1602_),
    .X(_1604_));
 sky130_fd_sc_hd__clkbuf_1 _3394_ (.A(_1604_),
    .X(_0336_));
 sky130_fd_sc_hd__mux2_1 _3395_ (.A0(_1558_),
    .A1(\tms1x00.RAM[47][2] ),
    .S(_1602_),
    .X(_1605_));
 sky130_fd_sc_hd__clkbuf_1 _3396_ (.A(_1605_),
    .X(_0337_));
 sky130_fd_sc_hd__mux2_1 _3397_ (.A0(_1560_),
    .A1(\tms1x00.RAM[47][3] ),
    .S(_1602_),
    .X(_1606_));
 sky130_fd_sc_hd__clkbuf_1 _3398_ (.A(_1606_),
    .X(_0338_));
 sky130_fd_sc_hd__or2_2 _3399_ (.A(_1199_),
    .B(_1496_),
    .X(_1607_));
 sky130_fd_sc_hd__mux2_1 _3400_ (.A0(_1553_),
    .A1(\tms1x00.RAM[46][0] ),
    .S(_1607_),
    .X(_1608_));
 sky130_fd_sc_hd__clkbuf_1 _3401_ (.A(_1608_),
    .X(_0339_));
 sky130_fd_sc_hd__mux2_1 _3402_ (.A0(_1556_),
    .A1(\tms1x00.RAM[46][1] ),
    .S(_1607_),
    .X(_1609_));
 sky130_fd_sc_hd__clkbuf_1 _3403_ (.A(_1609_),
    .X(_0340_));
 sky130_fd_sc_hd__mux2_1 _3404_ (.A0(_1558_),
    .A1(\tms1x00.RAM[46][2] ),
    .S(_1607_),
    .X(_1610_));
 sky130_fd_sc_hd__clkbuf_1 _3405_ (.A(_1610_),
    .X(_0341_));
 sky130_fd_sc_hd__mux2_1 _3406_ (.A0(_1560_),
    .A1(\tms1x00.RAM[46][3] ),
    .S(_1607_),
    .X(_1611_));
 sky130_fd_sc_hd__clkbuf_1 _3407_ (.A(_1611_),
    .X(_0342_));
 sky130_fd_sc_hd__or2_2 _3408_ (.A(_1145_),
    .B(_1254_),
    .X(_1612_));
 sky130_fd_sc_hd__mux2_1 _3409_ (.A0(_1553_),
    .A1(\tms1x00.RAM[54][0] ),
    .S(_1612_),
    .X(_1613_));
 sky130_fd_sc_hd__clkbuf_1 _3410_ (.A(_1613_),
    .X(_0343_));
 sky130_fd_sc_hd__mux2_1 _3411_ (.A0(_1556_),
    .A1(\tms1x00.RAM[54][1] ),
    .S(_1612_),
    .X(_1614_));
 sky130_fd_sc_hd__clkbuf_1 _3412_ (.A(_1614_),
    .X(_0344_));
 sky130_fd_sc_hd__mux2_1 _3413_ (.A0(_1558_),
    .A1(\tms1x00.RAM[54][2] ),
    .S(_1612_),
    .X(_1615_));
 sky130_fd_sc_hd__clkbuf_1 _3414_ (.A(_1615_),
    .X(_0345_));
 sky130_fd_sc_hd__mux2_1 _3415_ (.A0(_1560_),
    .A1(\tms1x00.RAM[54][3] ),
    .S(_1612_),
    .X(_1616_));
 sky130_fd_sc_hd__clkbuf_1 _3416_ (.A(_1616_),
    .X(_0346_));
 sky130_fd_sc_hd__buf_2 _3417_ (.A(_0820_),
    .X(_1617_));
 sky130_fd_sc_hd__or2_2 _3418_ (.A(_1145_),
    .B(_1163_),
    .X(_1618_));
 sky130_fd_sc_hd__mux2_1 _3419_ (.A0(_1617_),
    .A1(\tms1x00.RAM[53][0] ),
    .S(_1618_),
    .X(_1619_));
 sky130_fd_sc_hd__clkbuf_1 _3420_ (.A(_1619_),
    .X(_0347_));
 sky130_fd_sc_hd__buf_2 _3421_ (.A(_0929_),
    .X(_1620_));
 sky130_fd_sc_hd__mux2_1 _3422_ (.A0(_1620_),
    .A1(\tms1x00.RAM[53][1] ),
    .S(_1618_),
    .X(_1621_));
 sky130_fd_sc_hd__clkbuf_1 _3423_ (.A(_1621_),
    .X(_0348_));
 sky130_fd_sc_hd__buf_2 _3424_ (.A(_1029_),
    .X(_1622_));
 sky130_fd_sc_hd__mux2_1 _3425_ (.A0(_1622_),
    .A1(\tms1x00.RAM[53][2] ),
    .S(_1618_),
    .X(_1623_));
 sky130_fd_sc_hd__clkbuf_1 _3426_ (.A(_1623_),
    .X(_0349_));
 sky130_fd_sc_hd__buf_2 _3427_ (.A(_1127_),
    .X(_1624_));
 sky130_fd_sc_hd__mux2_1 _3428_ (.A0(_1624_),
    .A1(\tms1x00.RAM[53][3] ),
    .S(_1618_),
    .X(_1625_));
 sky130_fd_sc_hd__clkbuf_1 _3429_ (.A(_1625_),
    .X(_0350_));
 sky130_fd_sc_hd__or2_2 _3430_ (.A(_1144_),
    .B(_1293_),
    .X(_1626_));
 sky130_fd_sc_hd__mux2_1 _3431_ (.A0(_1617_),
    .A1(\tms1x00.RAM[52][0] ),
    .S(_1626_),
    .X(_1627_));
 sky130_fd_sc_hd__clkbuf_1 _3432_ (.A(_1627_),
    .X(_0351_));
 sky130_fd_sc_hd__mux2_1 _3433_ (.A0(_1620_),
    .A1(\tms1x00.RAM[52][1] ),
    .S(_1626_),
    .X(_1628_));
 sky130_fd_sc_hd__clkbuf_1 _3434_ (.A(_1628_),
    .X(_0352_));
 sky130_fd_sc_hd__mux2_1 _3435_ (.A0(_1622_),
    .A1(\tms1x00.RAM[52][2] ),
    .S(_1626_),
    .X(_1629_));
 sky130_fd_sc_hd__clkbuf_1 _3436_ (.A(_1629_),
    .X(_0353_));
 sky130_fd_sc_hd__mux2_1 _3437_ (.A0(_1624_),
    .A1(\tms1x00.RAM[52][3] ),
    .S(_1626_),
    .X(_1630_));
 sky130_fd_sc_hd__clkbuf_1 _3438_ (.A(_1630_),
    .X(_0354_));
 sky130_fd_sc_hd__or2_2 _3439_ (.A(_0827_),
    .B(_1144_),
    .X(_1631_));
 sky130_fd_sc_hd__mux2_1 _3440_ (.A0(_1617_),
    .A1(\tms1x00.RAM[51][0] ),
    .S(_1631_),
    .X(_1632_));
 sky130_fd_sc_hd__clkbuf_1 _3441_ (.A(_1632_),
    .X(_0355_));
 sky130_fd_sc_hd__mux2_1 _3442_ (.A0(_1620_),
    .A1(\tms1x00.RAM[51][1] ),
    .S(_1631_),
    .X(_1633_));
 sky130_fd_sc_hd__clkbuf_1 _3443_ (.A(_1633_),
    .X(_0356_));
 sky130_fd_sc_hd__mux2_1 _3444_ (.A0(_1622_),
    .A1(\tms1x00.RAM[51][2] ),
    .S(_1631_),
    .X(_1634_));
 sky130_fd_sc_hd__clkbuf_1 _3445_ (.A(_1634_),
    .X(_0357_));
 sky130_fd_sc_hd__mux2_1 _3446_ (.A0(_1624_),
    .A1(\tms1x00.RAM[51][3] ),
    .S(_1631_),
    .X(_1635_));
 sky130_fd_sc_hd__clkbuf_1 _3447_ (.A(_1635_),
    .X(_0358_));
 sky130_fd_sc_hd__nor2_2 _3448_ (.A(_1145_),
    .B(_1226_),
    .Y(_1636_));
 sky130_fd_sc_hd__mux2_1 _3449_ (.A0(\tms1x00.RAM[58][0] ),
    .A1(_1487_),
    .S(_1636_),
    .X(_1637_));
 sky130_fd_sc_hd__clkbuf_1 _3450_ (.A(_1637_),
    .X(_0359_));
 sky130_fd_sc_hd__mux2_1 _3451_ (.A0(\tms1x00.RAM[58][1] ),
    .A1(_1490_),
    .S(_1636_),
    .X(_1638_));
 sky130_fd_sc_hd__clkbuf_1 _3452_ (.A(_1638_),
    .X(_0360_));
 sky130_fd_sc_hd__mux2_1 _3453_ (.A0(\tms1x00.RAM[58][2] ),
    .A1(_1492_),
    .S(_1636_),
    .X(_1639_));
 sky130_fd_sc_hd__clkbuf_1 _3454_ (.A(_1639_),
    .X(_0361_));
 sky130_fd_sc_hd__mux2_1 _3455_ (.A0(\tms1x00.RAM[58][3] ),
    .A1(_1494_),
    .S(_1636_),
    .X(_1640_));
 sky130_fd_sc_hd__clkbuf_1 _3456_ (.A(_1640_),
    .X(_0362_));
 sky130_fd_sc_hd__nor2_2 _3457_ (.A(_1135_),
    .B(_1145_),
    .Y(_1641_));
 sky130_fd_sc_hd__mux2_1 _3458_ (.A0(\tms1x00.RAM[57][0] ),
    .A1(_1487_),
    .S(_1641_),
    .X(_1642_));
 sky130_fd_sc_hd__clkbuf_1 _3459_ (.A(_1642_),
    .X(_0363_));
 sky130_fd_sc_hd__mux2_1 _3460_ (.A0(\tms1x00.RAM[57][1] ),
    .A1(_1490_),
    .S(_1641_),
    .X(_1643_));
 sky130_fd_sc_hd__clkbuf_1 _3461_ (.A(_1643_),
    .X(_0364_));
 sky130_fd_sc_hd__mux2_1 _3462_ (.A0(\tms1x00.RAM[57][2] ),
    .A1(_1492_),
    .S(_1641_),
    .X(_1644_));
 sky130_fd_sc_hd__clkbuf_1 _3463_ (.A(_1644_),
    .X(_0365_));
 sky130_fd_sc_hd__mux2_1 _3464_ (.A0(\tms1x00.RAM[57][3] ),
    .A1(_1494_),
    .S(_1641_),
    .X(_1645_));
 sky130_fd_sc_hd__clkbuf_1 _3465_ (.A(_1645_),
    .X(_0366_));
 sky130_fd_sc_hd__nor2_2 _3466_ (.A(_1145_),
    .B(_1235_),
    .Y(_1646_));
 sky130_fd_sc_hd__mux2_1 _3467_ (.A0(\tms1x00.RAM[56][0] ),
    .A1(_1487_),
    .S(_1646_),
    .X(_1647_));
 sky130_fd_sc_hd__clkbuf_1 _3468_ (.A(_1647_),
    .X(_0367_));
 sky130_fd_sc_hd__mux2_1 _3469_ (.A0(\tms1x00.RAM[56][1] ),
    .A1(_1490_),
    .S(_1646_),
    .X(_1648_));
 sky130_fd_sc_hd__clkbuf_1 _3470_ (.A(_1648_),
    .X(_0368_));
 sky130_fd_sc_hd__mux2_1 _3471_ (.A0(\tms1x00.RAM[56][2] ),
    .A1(_1492_),
    .S(_1646_),
    .X(_1649_));
 sky130_fd_sc_hd__clkbuf_1 _3472_ (.A(_1649_),
    .X(_0369_));
 sky130_fd_sc_hd__mux2_1 _3473_ (.A0(\tms1x00.RAM[56][3] ),
    .A1(_1494_),
    .S(_1646_),
    .X(_1650_));
 sky130_fd_sc_hd__clkbuf_1 _3474_ (.A(_1650_),
    .X(_0370_));
 sky130_fd_sc_hd__nor2_2 _3475_ (.A(_1145_),
    .B(_1247_),
    .Y(_1651_));
 sky130_fd_sc_hd__mux2_1 _3476_ (.A0(\tms1x00.RAM[55][0] ),
    .A1(_1487_),
    .S(_1651_),
    .X(_1652_));
 sky130_fd_sc_hd__clkbuf_1 _3477_ (.A(_1652_),
    .X(_0371_));
 sky130_fd_sc_hd__mux2_1 _3478_ (.A0(\tms1x00.RAM[55][1] ),
    .A1(_1490_),
    .S(_1651_),
    .X(_1653_));
 sky130_fd_sc_hd__clkbuf_1 _3479_ (.A(_1653_),
    .X(_0372_));
 sky130_fd_sc_hd__mux2_1 _3480_ (.A0(\tms1x00.RAM[55][2] ),
    .A1(_1492_),
    .S(_1651_),
    .X(_1654_));
 sky130_fd_sc_hd__clkbuf_1 _3481_ (.A(_1654_),
    .X(_0373_));
 sky130_fd_sc_hd__mux2_1 _3482_ (.A0(\tms1x00.RAM[55][3] ),
    .A1(_1494_),
    .S(_1651_),
    .X(_1655_));
 sky130_fd_sc_hd__clkbuf_1 _3483_ (.A(_1655_),
    .X(_0374_));
 sky130_fd_sc_hd__or2_2 _3484_ (.A(_1144_),
    .B(_1169_),
    .X(_1656_));
 sky130_fd_sc_hd__mux2_1 _3485_ (.A0(_1617_),
    .A1(\tms1x00.RAM[63][0] ),
    .S(_1656_),
    .X(_1657_));
 sky130_fd_sc_hd__clkbuf_1 _3486_ (.A(_1657_),
    .X(_0375_));
 sky130_fd_sc_hd__mux2_1 _3487_ (.A0(_1620_),
    .A1(\tms1x00.RAM[63][1] ),
    .S(_1656_),
    .X(_1658_));
 sky130_fd_sc_hd__clkbuf_1 _3488_ (.A(_1658_),
    .X(_0376_));
 sky130_fd_sc_hd__mux2_1 _3489_ (.A0(_1622_),
    .A1(\tms1x00.RAM[63][2] ),
    .S(_1656_),
    .X(_1659_));
 sky130_fd_sc_hd__clkbuf_1 _3490_ (.A(_1659_),
    .X(_0377_));
 sky130_fd_sc_hd__mux2_1 _3491_ (.A0(_1624_),
    .A1(\tms1x00.RAM[63][3] ),
    .S(_1656_),
    .X(_1660_));
 sky130_fd_sc_hd__clkbuf_1 _3492_ (.A(_1660_),
    .X(_0378_));
 sky130_fd_sc_hd__or2_2 _3493_ (.A(_1144_),
    .B(_1199_),
    .X(_1661_));
 sky130_fd_sc_hd__mux2_1 _3494_ (.A0(_1617_),
    .A1(\tms1x00.RAM[62][0] ),
    .S(_1661_),
    .X(_1662_));
 sky130_fd_sc_hd__clkbuf_1 _3495_ (.A(_1662_),
    .X(_0379_));
 sky130_fd_sc_hd__mux2_1 _3496_ (.A0(_1620_),
    .A1(\tms1x00.RAM[62][1] ),
    .S(_1661_),
    .X(_1663_));
 sky130_fd_sc_hd__clkbuf_1 _3497_ (.A(_1663_),
    .X(_0380_));
 sky130_fd_sc_hd__mux2_1 _3498_ (.A0(_1622_),
    .A1(\tms1x00.RAM[62][2] ),
    .S(_1661_),
    .X(_1664_));
 sky130_fd_sc_hd__clkbuf_1 _3499_ (.A(_1664_),
    .X(_0381_));
 sky130_fd_sc_hd__mux2_1 _3500_ (.A0(_1624_),
    .A1(\tms1x00.RAM[62][3] ),
    .S(_1661_),
    .X(_1665_));
 sky130_fd_sc_hd__clkbuf_1 _3501_ (.A(_1665_),
    .X(_0382_));
 sky130_fd_sc_hd__or2_2 _3502_ (.A(_1144_),
    .B(_1154_),
    .X(_1666_));
 sky130_fd_sc_hd__mux2_1 _3503_ (.A0(_1617_),
    .A1(\tms1x00.RAM[61][0] ),
    .S(_1666_),
    .X(_1667_));
 sky130_fd_sc_hd__clkbuf_1 _3504_ (.A(_1667_),
    .X(_0383_));
 sky130_fd_sc_hd__mux2_1 _3505_ (.A0(_1620_),
    .A1(\tms1x00.RAM[61][1] ),
    .S(_1666_),
    .X(_1668_));
 sky130_fd_sc_hd__clkbuf_1 _3506_ (.A(_1668_),
    .X(_0384_));
 sky130_fd_sc_hd__mux2_1 _3507_ (.A0(_1622_),
    .A1(\tms1x00.RAM[61][2] ),
    .S(_1666_),
    .X(_1669_));
 sky130_fd_sc_hd__clkbuf_1 _3508_ (.A(_1669_),
    .X(_0385_));
 sky130_fd_sc_hd__mux2_1 _3509_ (.A0(_1624_),
    .A1(\tms1x00.RAM[61][3] ),
    .S(_1666_),
    .X(_1670_));
 sky130_fd_sc_hd__clkbuf_1 _3510_ (.A(_1670_),
    .X(_0386_));
 sky130_fd_sc_hd__or2_2 _3511_ (.A(_1144_),
    .B(_1211_),
    .X(_1671_));
 sky130_fd_sc_hd__mux2_1 _3512_ (.A0(_1617_),
    .A1(\tms1x00.RAM[60][0] ),
    .S(_1671_),
    .X(_1672_));
 sky130_fd_sc_hd__clkbuf_1 _3513_ (.A(_1672_),
    .X(_0387_));
 sky130_fd_sc_hd__mux2_1 _3514_ (.A0(_1620_),
    .A1(\tms1x00.RAM[60][1] ),
    .S(_1671_),
    .X(_1673_));
 sky130_fd_sc_hd__clkbuf_1 _3515_ (.A(_1673_),
    .X(_0388_));
 sky130_fd_sc_hd__mux2_1 _3516_ (.A0(_1622_),
    .A1(\tms1x00.RAM[60][2] ),
    .S(_1671_),
    .X(_1674_));
 sky130_fd_sc_hd__clkbuf_1 _3517_ (.A(_1674_),
    .X(_0389_));
 sky130_fd_sc_hd__mux2_1 _3518_ (.A0(_1624_),
    .A1(\tms1x00.RAM[60][3] ),
    .S(_1671_),
    .X(_1675_));
 sky130_fd_sc_hd__clkbuf_1 _3519_ (.A(_1675_),
    .X(_0390_));
 sky130_fd_sc_hd__or2_2 _3520_ (.A(_1163_),
    .B(_1232_),
    .X(_1676_));
 sky130_fd_sc_hd__mux2_1 _3521_ (.A0(_1617_),
    .A1(\tms1x00.RAM[5][0] ),
    .S(_1676_),
    .X(_1677_));
 sky130_fd_sc_hd__clkbuf_1 _3522_ (.A(_1677_),
    .X(_0391_));
 sky130_fd_sc_hd__mux2_1 _3523_ (.A0(_1620_),
    .A1(\tms1x00.RAM[5][1] ),
    .S(_1676_),
    .X(_1678_));
 sky130_fd_sc_hd__clkbuf_1 _3524_ (.A(_1678_),
    .X(_0392_));
 sky130_fd_sc_hd__mux2_1 _3525_ (.A0(_1622_),
    .A1(\tms1x00.RAM[5][2] ),
    .S(_1676_),
    .X(_1679_));
 sky130_fd_sc_hd__clkbuf_1 _3526_ (.A(_1679_),
    .X(_0393_));
 sky130_fd_sc_hd__mux2_1 _3527_ (.A0(_1624_),
    .A1(\tms1x00.RAM[5][3] ),
    .S(_1676_),
    .X(_1680_));
 sky130_fd_sc_hd__clkbuf_1 _3528_ (.A(_1680_),
    .X(_0394_));
 sky130_fd_sc_hd__or2_2 _3529_ (.A(_0827_),
    .B(_1160_),
    .X(_1681_));
 sky130_fd_sc_hd__mux2_1 _3530_ (.A0(_1617_),
    .A1(\tms1x00.RAM[67][0] ),
    .S(_1681_),
    .X(_1682_));
 sky130_fd_sc_hd__clkbuf_1 _3531_ (.A(_1682_),
    .X(_0395_));
 sky130_fd_sc_hd__mux2_1 _3532_ (.A0(_1620_),
    .A1(\tms1x00.RAM[67][1] ),
    .S(_1681_),
    .X(_1683_));
 sky130_fd_sc_hd__clkbuf_1 _3533_ (.A(_1683_),
    .X(_0396_));
 sky130_fd_sc_hd__mux2_1 _3534_ (.A0(_1622_),
    .A1(\tms1x00.RAM[67][2] ),
    .S(_1681_),
    .X(_1684_));
 sky130_fd_sc_hd__clkbuf_1 _3535_ (.A(_1684_),
    .X(_0397_));
 sky130_fd_sc_hd__mux2_1 _3536_ (.A0(_1624_),
    .A1(\tms1x00.RAM[67][3] ),
    .S(_1681_),
    .X(_1685_));
 sky130_fd_sc_hd__clkbuf_1 _3537_ (.A(_1685_),
    .X(_0398_));
 sky130_fd_sc_hd__or2_2 _3538_ (.A(_1161_),
    .B(_1305_),
    .X(_1686_));
 sky130_fd_sc_hd__mux2_1 _3539_ (.A0(_1617_),
    .A1(\tms1x00.RAM[66][0] ),
    .S(_1686_),
    .X(_1687_));
 sky130_fd_sc_hd__clkbuf_1 _3540_ (.A(_1687_),
    .X(_0399_));
 sky130_fd_sc_hd__mux2_1 _3541_ (.A0(_1620_),
    .A1(\tms1x00.RAM[66][1] ),
    .S(_1686_),
    .X(_1688_));
 sky130_fd_sc_hd__clkbuf_1 _3542_ (.A(_1688_),
    .X(_0400_));
 sky130_fd_sc_hd__mux2_1 _3543_ (.A0(_1622_),
    .A1(\tms1x00.RAM[66][2] ),
    .S(_1686_),
    .X(_1689_));
 sky130_fd_sc_hd__clkbuf_1 _3544_ (.A(_1689_),
    .X(_0401_));
 sky130_fd_sc_hd__mux2_1 _3545_ (.A0(_1624_),
    .A1(\tms1x00.RAM[66][3] ),
    .S(_1686_),
    .X(_1690_));
 sky130_fd_sc_hd__clkbuf_1 _3546_ (.A(_1690_),
    .X(_0402_));
 sky130_fd_sc_hd__clkbuf_4 _3547_ (.A(_0820_),
    .X(_1691_));
 sky130_fd_sc_hd__or2_2 _3548_ (.A(_1161_),
    .B(_1182_),
    .X(_1692_));
 sky130_fd_sc_hd__mux2_1 _3549_ (.A0(_1691_),
    .A1(\tms1x00.RAM[65][0] ),
    .S(_1692_),
    .X(_1693_));
 sky130_fd_sc_hd__clkbuf_1 _3550_ (.A(_1693_),
    .X(_0403_));
 sky130_fd_sc_hd__buf_2 _3551_ (.A(_0929_),
    .X(_1694_));
 sky130_fd_sc_hd__mux2_1 _3552_ (.A0(_1694_),
    .A1(\tms1x00.RAM[65][1] ),
    .S(_1692_),
    .X(_1695_));
 sky130_fd_sc_hd__clkbuf_1 _3553_ (.A(_1695_),
    .X(_0404_));
 sky130_fd_sc_hd__clkbuf_4 _3554_ (.A(_1029_),
    .X(_1696_));
 sky130_fd_sc_hd__mux2_1 _3555_ (.A0(_1696_),
    .A1(\tms1x00.RAM[65][2] ),
    .S(_1692_),
    .X(_1697_));
 sky130_fd_sc_hd__clkbuf_1 _3556_ (.A(_1697_),
    .X(_0405_));
 sky130_fd_sc_hd__clkbuf_4 _3557_ (.A(_1127_),
    .X(_1698_));
 sky130_fd_sc_hd__mux2_1 _3558_ (.A0(_1698_),
    .A1(\tms1x00.RAM[65][3] ),
    .S(_1692_),
    .X(_1699_));
 sky130_fd_sc_hd__clkbuf_1 _3559_ (.A(_1699_),
    .X(_0406_));
 sky130_fd_sc_hd__or2_2 _3560_ (.A(_1161_),
    .B(_1299_),
    .X(_1700_));
 sky130_fd_sc_hd__mux2_1 _3561_ (.A0(_1691_),
    .A1(\tms1x00.RAM[64][0] ),
    .S(_1700_),
    .X(_1701_));
 sky130_fd_sc_hd__clkbuf_1 _3562_ (.A(_1701_),
    .X(_0407_));
 sky130_fd_sc_hd__mux2_1 _3563_ (.A0(_1694_),
    .A1(\tms1x00.RAM[64][1] ),
    .S(_1700_),
    .X(_1702_));
 sky130_fd_sc_hd__clkbuf_1 _3564_ (.A(_1702_),
    .X(_0408_));
 sky130_fd_sc_hd__mux2_1 _3565_ (.A0(_1696_),
    .A1(\tms1x00.RAM[64][2] ),
    .S(_1700_),
    .X(_1703_));
 sky130_fd_sc_hd__clkbuf_1 _3566_ (.A(_1703_),
    .X(_0409_));
 sky130_fd_sc_hd__mux2_1 _3567_ (.A0(_1698_),
    .A1(\tms1x00.RAM[64][3] ),
    .S(_1700_),
    .X(_1704_));
 sky130_fd_sc_hd__clkbuf_1 _3568_ (.A(_1704_),
    .X(_0410_));
 sky130_fd_sc_hd__nor2_2 _3569_ (.A(_1161_),
    .B(_1247_),
    .Y(_1705_));
 sky130_fd_sc_hd__mux2_1 _3570_ (.A0(\tms1x00.RAM[71][0] ),
    .A1(_1487_),
    .S(_1705_),
    .X(_1706_));
 sky130_fd_sc_hd__clkbuf_1 _3571_ (.A(_1706_),
    .X(_0411_));
 sky130_fd_sc_hd__mux2_1 _3572_ (.A0(\tms1x00.RAM[71][1] ),
    .A1(_1490_),
    .S(_1705_),
    .X(_1707_));
 sky130_fd_sc_hd__clkbuf_1 _3573_ (.A(_1707_),
    .X(_0412_));
 sky130_fd_sc_hd__mux2_1 _3574_ (.A0(\tms1x00.RAM[71][2] ),
    .A1(_1492_),
    .S(_1705_),
    .X(_1708_));
 sky130_fd_sc_hd__clkbuf_1 _3575_ (.A(_1708_),
    .X(_0413_));
 sky130_fd_sc_hd__mux2_1 _3576_ (.A0(\tms1x00.RAM[71][3] ),
    .A1(_1494_),
    .S(_1705_),
    .X(_1709_));
 sky130_fd_sc_hd__clkbuf_1 _3577_ (.A(_1709_),
    .X(_0414_));
 sky130_fd_sc_hd__or2_2 _3578_ (.A(_1160_),
    .B(_1254_),
    .X(_1710_));
 sky130_fd_sc_hd__mux2_1 _3579_ (.A0(_1691_),
    .A1(\tms1x00.RAM[70][0] ),
    .S(_1710_),
    .X(_1711_));
 sky130_fd_sc_hd__clkbuf_1 _3580_ (.A(_1711_),
    .X(_0415_));
 sky130_fd_sc_hd__mux2_1 _3581_ (.A0(_1694_),
    .A1(\tms1x00.RAM[70][1] ),
    .S(_1710_),
    .X(_1712_));
 sky130_fd_sc_hd__clkbuf_1 _3582_ (.A(_1712_),
    .X(_0416_));
 sky130_fd_sc_hd__mux2_1 _3583_ (.A0(_1696_),
    .A1(\tms1x00.RAM[70][2] ),
    .S(_1710_),
    .X(_1713_));
 sky130_fd_sc_hd__clkbuf_1 _3584_ (.A(_1713_),
    .X(_0417_));
 sky130_fd_sc_hd__mux2_1 _3585_ (.A0(_1698_),
    .A1(\tms1x00.RAM[70][3] ),
    .S(_1710_),
    .X(_1714_));
 sky130_fd_sc_hd__clkbuf_1 _3586_ (.A(_1714_),
    .X(_0418_));
 sky130_fd_sc_hd__or2_2 _3587_ (.A(_1233_),
    .B(_1254_),
    .X(_1715_));
 sky130_fd_sc_hd__mux2_1 _3588_ (.A0(_1691_),
    .A1(\tms1x00.RAM[6][0] ),
    .S(_1715_),
    .X(_1716_));
 sky130_fd_sc_hd__clkbuf_1 _3589_ (.A(_1716_),
    .X(_0419_));
 sky130_fd_sc_hd__mux2_1 _3590_ (.A0(_1694_),
    .A1(\tms1x00.RAM[6][1] ),
    .S(_1715_),
    .X(_1717_));
 sky130_fd_sc_hd__clkbuf_1 _3591_ (.A(_1717_),
    .X(_0420_));
 sky130_fd_sc_hd__mux2_1 _3592_ (.A0(_1696_),
    .A1(\tms1x00.RAM[6][2] ),
    .S(_1715_),
    .X(_1718_));
 sky130_fd_sc_hd__clkbuf_1 _3593_ (.A(_1718_),
    .X(_0421_));
 sky130_fd_sc_hd__mux2_1 _3594_ (.A0(_1698_),
    .A1(\tms1x00.RAM[6][3] ),
    .S(_1715_),
    .X(_1719_));
 sky130_fd_sc_hd__clkbuf_1 _3595_ (.A(_1719_),
    .X(_0422_));
 sky130_fd_sc_hd__or2_2 _3596_ (.A(_1160_),
    .B(_1293_),
    .X(_1720_));
 sky130_fd_sc_hd__mux2_1 _3597_ (.A0(_1691_),
    .A1(\tms1x00.RAM[68][0] ),
    .S(_1720_),
    .X(_1721_));
 sky130_fd_sc_hd__clkbuf_1 _3598_ (.A(_1721_),
    .X(_0423_));
 sky130_fd_sc_hd__mux2_1 _3599_ (.A0(_1694_),
    .A1(\tms1x00.RAM[68][1] ),
    .S(_1720_),
    .X(_1722_));
 sky130_fd_sc_hd__clkbuf_1 _3600_ (.A(_1722_),
    .X(_0424_));
 sky130_fd_sc_hd__mux2_1 _3601_ (.A0(_1696_),
    .A1(\tms1x00.RAM[68][2] ),
    .S(_1720_),
    .X(_1723_));
 sky130_fd_sc_hd__clkbuf_1 _3602_ (.A(_1723_),
    .X(_0425_));
 sky130_fd_sc_hd__mux2_1 _3603_ (.A0(_1698_),
    .A1(\tms1x00.RAM[68][3] ),
    .S(_1720_),
    .X(_1724_));
 sky130_fd_sc_hd__clkbuf_1 _3604_ (.A(_1724_),
    .X(_0426_));
 sky130_fd_sc_hd__or2_2 _3605_ (.A(_1160_),
    .B(_1211_),
    .X(_1725_));
 sky130_fd_sc_hd__mux2_1 _3606_ (.A0(_1691_),
    .A1(\tms1x00.RAM[76][0] ),
    .S(_1725_),
    .X(_1726_));
 sky130_fd_sc_hd__clkbuf_1 _3607_ (.A(_1726_),
    .X(_0427_));
 sky130_fd_sc_hd__mux2_1 _3608_ (.A0(_1694_),
    .A1(\tms1x00.RAM[76][1] ),
    .S(_1725_),
    .X(_1727_));
 sky130_fd_sc_hd__clkbuf_1 _3609_ (.A(_1727_),
    .X(_0428_));
 sky130_fd_sc_hd__mux2_1 _3610_ (.A0(_1696_),
    .A1(\tms1x00.RAM[76][2] ),
    .S(_1725_),
    .X(_1728_));
 sky130_fd_sc_hd__clkbuf_1 _3611_ (.A(_1728_),
    .X(_0429_));
 sky130_fd_sc_hd__mux2_1 _3612_ (.A0(_1698_),
    .A1(\tms1x00.RAM[76][3] ),
    .S(_1725_),
    .X(_1729_));
 sky130_fd_sc_hd__clkbuf_1 _3613_ (.A(_1729_),
    .X(_0430_));
 sky130_fd_sc_hd__nor2_2 _3614_ (.A(_1147_),
    .B(_1161_),
    .Y(_1730_));
 sky130_fd_sc_hd__mux2_1 _3615_ (.A0(\tms1x00.RAM[75][0] ),
    .A1(_1265_),
    .S(_1730_),
    .X(_1731_));
 sky130_fd_sc_hd__clkbuf_1 _3616_ (.A(_1731_),
    .X(_0431_));
 sky130_fd_sc_hd__mux2_1 _3617_ (.A0(\tms1x00.RAM[75][1] ),
    .A1(_1269_),
    .S(_1730_),
    .X(_1732_));
 sky130_fd_sc_hd__clkbuf_1 _3618_ (.A(_1732_),
    .X(_0432_));
 sky130_fd_sc_hd__mux2_1 _3619_ (.A0(\tms1x00.RAM[75][2] ),
    .A1(_1272_),
    .S(_1730_),
    .X(_1733_));
 sky130_fd_sc_hd__clkbuf_1 _3620_ (.A(_1733_),
    .X(_0433_));
 sky130_fd_sc_hd__mux2_1 _3621_ (.A0(\tms1x00.RAM[75][3] ),
    .A1(_1275_),
    .S(_1730_),
    .X(_1734_));
 sky130_fd_sc_hd__clkbuf_1 _3622_ (.A(_1734_),
    .X(_0434_));
 sky130_fd_sc_hd__nor2_2 _3623_ (.A(_1161_),
    .B(_1226_),
    .Y(_1735_));
 sky130_fd_sc_hd__mux2_1 _3624_ (.A0(\tms1x00.RAM[74][0] ),
    .A1(_1265_),
    .S(_1735_),
    .X(_1736_));
 sky130_fd_sc_hd__clkbuf_1 _3625_ (.A(_1736_),
    .X(_0435_));
 sky130_fd_sc_hd__mux2_1 _3626_ (.A0(\tms1x00.RAM[74][1] ),
    .A1(_1269_),
    .S(_1735_),
    .X(_1737_));
 sky130_fd_sc_hd__clkbuf_1 _3627_ (.A(_1737_),
    .X(_0436_));
 sky130_fd_sc_hd__mux2_1 _3628_ (.A0(\tms1x00.RAM[74][2] ),
    .A1(_1272_),
    .S(_1735_),
    .X(_1738_));
 sky130_fd_sc_hd__clkbuf_1 _3629_ (.A(_1738_),
    .X(_0437_));
 sky130_fd_sc_hd__mux2_1 _3630_ (.A0(\tms1x00.RAM[74][3] ),
    .A1(_1275_),
    .S(_1735_),
    .X(_1739_));
 sky130_fd_sc_hd__clkbuf_1 _3631_ (.A(_1739_),
    .X(_0438_));
 sky130_fd_sc_hd__nor2_2 _3632_ (.A(_1135_),
    .B(_1161_),
    .Y(_1740_));
 sky130_fd_sc_hd__mux2_1 _3633_ (.A0(\tms1x00.RAM[73][0] ),
    .A1(_1265_),
    .S(_1740_),
    .X(_1741_));
 sky130_fd_sc_hd__clkbuf_1 _3634_ (.A(_1741_),
    .X(_0439_));
 sky130_fd_sc_hd__mux2_1 _3635_ (.A0(\tms1x00.RAM[73][1] ),
    .A1(_1269_),
    .S(_1740_),
    .X(_1742_));
 sky130_fd_sc_hd__clkbuf_1 _3636_ (.A(_1742_),
    .X(_0440_));
 sky130_fd_sc_hd__mux2_1 _3637_ (.A0(\tms1x00.RAM[73][2] ),
    .A1(_1272_),
    .S(_1740_),
    .X(_1743_));
 sky130_fd_sc_hd__clkbuf_1 _3638_ (.A(_1743_),
    .X(_0441_));
 sky130_fd_sc_hd__mux2_1 _3639_ (.A0(\tms1x00.RAM[73][3] ),
    .A1(_1275_),
    .S(_1740_),
    .X(_1744_));
 sky130_fd_sc_hd__clkbuf_1 _3640_ (.A(_1744_),
    .X(_0442_));
 sky130_fd_sc_hd__nor2_2 _3641_ (.A(_1161_),
    .B(_1235_),
    .Y(_1745_));
 sky130_fd_sc_hd__mux2_1 _3642_ (.A0(\tms1x00.RAM[72][0] ),
    .A1(_1265_),
    .S(_1745_),
    .X(_1746_));
 sky130_fd_sc_hd__clkbuf_1 _3643_ (.A(_1746_),
    .X(_0443_));
 sky130_fd_sc_hd__mux2_1 _3644_ (.A0(\tms1x00.RAM[72][1] ),
    .A1(_1269_),
    .S(_1745_),
    .X(_1747_));
 sky130_fd_sc_hd__clkbuf_1 _3645_ (.A(_1747_),
    .X(_0444_));
 sky130_fd_sc_hd__mux2_1 _3646_ (.A0(\tms1x00.RAM[72][2] ),
    .A1(_1272_),
    .S(_1745_),
    .X(_1748_));
 sky130_fd_sc_hd__clkbuf_1 _3647_ (.A(_1748_),
    .X(_0445_));
 sky130_fd_sc_hd__mux2_1 _3648_ (.A0(\tms1x00.RAM[72][3] ),
    .A1(_1275_),
    .S(_1745_),
    .X(_1749_));
 sky130_fd_sc_hd__clkbuf_1 _3649_ (.A(_1749_),
    .X(_0446_));
 sky130_fd_sc_hd__or2_2 _3650_ (.A(_1154_),
    .B(_1160_),
    .X(_1750_));
 sky130_fd_sc_hd__mux2_1 _3651_ (.A0(_1691_),
    .A1(\tms1x00.RAM[77][0] ),
    .S(_1750_),
    .X(_1751_));
 sky130_fd_sc_hd__clkbuf_1 _3652_ (.A(_1751_),
    .X(_0447_));
 sky130_fd_sc_hd__mux2_1 _3653_ (.A0(_1694_),
    .A1(\tms1x00.RAM[77][1] ),
    .S(_1750_),
    .X(_1752_));
 sky130_fd_sc_hd__clkbuf_1 _3654_ (.A(_1752_),
    .X(_0448_));
 sky130_fd_sc_hd__mux2_1 _3655_ (.A0(_1696_),
    .A1(\tms1x00.RAM[77][2] ),
    .S(_1750_),
    .X(_1753_));
 sky130_fd_sc_hd__clkbuf_1 _3656_ (.A(_1753_),
    .X(_0449_));
 sky130_fd_sc_hd__mux2_1 _3657_ (.A0(_1698_),
    .A1(\tms1x00.RAM[77][3] ),
    .S(_1750_),
    .X(_1754_));
 sky130_fd_sc_hd__clkbuf_1 _3658_ (.A(_1754_),
    .X(_0450_));
 sky130_fd_sc_hd__or2_2 _3659_ (.A(_1131_),
    .B(_1299_),
    .X(_1755_));
 sky130_fd_sc_hd__mux2_1 _3660_ (.A0(_1691_),
    .A1(\tms1x00.RAM[80][0] ),
    .S(_1755_),
    .X(_1756_));
 sky130_fd_sc_hd__clkbuf_1 _3661_ (.A(_1756_),
    .X(_0451_));
 sky130_fd_sc_hd__mux2_1 _3662_ (.A0(_1694_),
    .A1(\tms1x00.RAM[80][1] ),
    .S(_1755_),
    .X(_1757_));
 sky130_fd_sc_hd__clkbuf_1 _3663_ (.A(_1757_),
    .X(_0452_));
 sky130_fd_sc_hd__mux2_1 _3664_ (.A0(_1696_),
    .A1(\tms1x00.RAM[80][2] ),
    .S(_1755_),
    .X(_1758_));
 sky130_fd_sc_hd__clkbuf_1 _3665_ (.A(_1758_),
    .X(_0453_));
 sky130_fd_sc_hd__mux2_1 _3666_ (.A0(_1698_),
    .A1(\tms1x00.RAM[80][3] ),
    .S(_1755_),
    .X(_1759_));
 sky130_fd_sc_hd__clkbuf_1 _3667_ (.A(_1759_),
    .X(_0454_));
 sky130_fd_sc_hd__nor2_2 _3668_ (.A(_1233_),
    .B(_1247_),
    .Y(_1760_));
 sky130_fd_sc_hd__mux2_1 _3669_ (.A0(\tms1x00.RAM[7][0] ),
    .A1(_1265_),
    .S(_1760_),
    .X(_1761_));
 sky130_fd_sc_hd__clkbuf_1 _3670_ (.A(_1761_),
    .X(_0455_));
 sky130_fd_sc_hd__mux2_1 _3671_ (.A0(\tms1x00.RAM[7][1] ),
    .A1(_1269_),
    .S(_1760_),
    .X(_1762_));
 sky130_fd_sc_hd__clkbuf_1 _3672_ (.A(_1762_),
    .X(_0456_));
 sky130_fd_sc_hd__mux2_1 _3673_ (.A0(\tms1x00.RAM[7][2] ),
    .A1(_1272_),
    .S(_1760_),
    .X(_1763_));
 sky130_fd_sc_hd__clkbuf_1 _3674_ (.A(_1763_),
    .X(_0457_));
 sky130_fd_sc_hd__mux2_1 _3675_ (.A0(\tms1x00.RAM[7][3] ),
    .A1(_1275_),
    .S(_1760_),
    .X(_1764_));
 sky130_fd_sc_hd__clkbuf_1 _3676_ (.A(_1764_),
    .X(_0458_));
 sky130_fd_sc_hd__or2_2 _3677_ (.A(_1160_),
    .B(_1199_),
    .X(_1765_));
 sky130_fd_sc_hd__mux2_1 _3678_ (.A0(_1691_),
    .A1(\tms1x00.RAM[78][0] ),
    .S(_1765_),
    .X(_1766_));
 sky130_fd_sc_hd__clkbuf_1 _3679_ (.A(_1766_),
    .X(_0459_));
 sky130_fd_sc_hd__mux2_1 _3680_ (.A0(_1694_),
    .A1(\tms1x00.RAM[78][1] ),
    .S(_1765_),
    .X(_1767_));
 sky130_fd_sc_hd__clkbuf_1 _3681_ (.A(_1767_),
    .X(_0460_));
 sky130_fd_sc_hd__mux2_1 _3682_ (.A0(_1696_),
    .A1(\tms1x00.RAM[78][2] ),
    .S(_1765_),
    .X(_1768_));
 sky130_fd_sc_hd__clkbuf_1 _3683_ (.A(_1768_),
    .X(_0461_));
 sky130_fd_sc_hd__mux2_1 _3684_ (.A0(_1698_),
    .A1(\tms1x00.RAM[78][3] ),
    .S(_1765_),
    .X(_1769_));
 sky130_fd_sc_hd__clkbuf_1 _3685_ (.A(_1769_),
    .X(_0462_));
 sky130_fd_sc_hd__or2_2 _3686_ (.A(_1131_),
    .B(_1163_),
    .X(_1770_));
 sky130_fd_sc_hd__mux2_1 _3687_ (.A0(_1691_),
    .A1(\tms1x00.RAM[85][0] ),
    .S(_1770_),
    .X(_1771_));
 sky130_fd_sc_hd__clkbuf_1 _3688_ (.A(_1771_),
    .X(_0463_));
 sky130_fd_sc_hd__mux2_1 _3689_ (.A0(_1694_),
    .A1(\tms1x00.RAM[85][1] ),
    .S(_1770_),
    .X(_1772_));
 sky130_fd_sc_hd__clkbuf_1 _3690_ (.A(_1772_),
    .X(_0464_));
 sky130_fd_sc_hd__mux2_1 _3691_ (.A0(_1696_),
    .A1(\tms1x00.RAM[85][2] ),
    .S(_1770_),
    .X(_1773_));
 sky130_fd_sc_hd__clkbuf_1 _3692_ (.A(_1773_),
    .X(_0465_));
 sky130_fd_sc_hd__mux2_1 _3693_ (.A0(_1698_),
    .A1(\tms1x00.RAM[85][3] ),
    .S(_1770_),
    .X(_1774_));
 sky130_fd_sc_hd__clkbuf_1 _3694_ (.A(_1774_),
    .X(_0466_));
 sky130_fd_sc_hd__buf_2 _3695_ (.A(_0820_),
    .X(_1775_));
 sky130_fd_sc_hd__or2_2 _3696_ (.A(_1131_),
    .B(_1293_),
    .X(_1776_));
 sky130_fd_sc_hd__mux2_1 _3697_ (.A0(_1775_),
    .A1(\tms1x00.RAM[84][0] ),
    .S(_1776_),
    .X(_1777_));
 sky130_fd_sc_hd__clkbuf_1 _3698_ (.A(_1777_),
    .X(_0467_));
 sky130_fd_sc_hd__buf_2 _3699_ (.A(_0929_),
    .X(_1778_));
 sky130_fd_sc_hd__mux2_1 _3700_ (.A0(_1778_),
    .A1(\tms1x00.RAM[84][1] ),
    .S(_1776_),
    .X(_1779_));
 sky130_fd_sc_hd__clkbuf_1 _3701_ (.A(_1779_),
    .X(_0468_));
 sky130_fd_sc_hd__buf_2 _3702_ (.A(_1029_),
    .X(_1780_));
 sky130_fd_sc_hd__mux2_1 _3703_ (.A0(_1780_),
    .A1(\tms1x00.RAM[84][2] ),
    .S(_1776_),
    .X(_1781_));
 sky130_fd_sc_hd__clkbuf_1 _3704_ (.A(_1781_),
    .X(_0469_));
 sky130_fd_sc_hd__buf_2 _3705_ (.A(_1127_),
    .X(_1782_));
 sky130_fd_sc_hd__mux2_1 _3706_ (.A0(_1782_),
    .A1(\tms1x00.RAM[84][3] ),
    .S(_1776_),
    .X(_1783_));
 sky130_fd_sc_hd__clkbuf_1 _3707_ (.A(_1783_),
    .X(_0470_));
 sky130_fd_sc_hd__or2_2 _3708_ (.A(_0827_),
    .B(_1131_),
    .X(_1784_));
 sky130_fd_sc_hd__mux2_1 _3709_ (.A0(_1775_),
    .A1(\tms1x00.RAM[83][0] ),
    .S(_1784_),
    .X(_1785_));
 sky130_fd_sc_hd__clkbuf_1 _3710_ (.A(_1785_),
    .X(_0471_));
 sky130_fd_sc_hd__mux2_1 _3711_ (.A0(_1778_),
    .A1(\tms1x00.RAM[83][1] ),
    .S(_1784_),
    .X(_1786_));
 sky130_fd_sc_hd__clkbuf_1 _3712_ (.A(_1786_),
    .X(_0472_));
 sky130_fd_sc_hd__mux2_1 _3713_ (.A0(_1780_),
    .A1(\tms1x00.RAM[83][2] ),
    .S(_1784_),
    .X(_1787_));
 sky130_fd_sc_hd__clkbuf_1 _3714_ (.A(_1787_),
    .X(_0473_));
 sky130_fd_sc_hd__mux2_1 _3715_ (.A0(_1782_),
    .A1(\tms1x00.RAM[83][3] ),
    .S(_1784_),
    .X(_1788_));
 sky130_fd_sc_hd__clkbuf_1 _3716_ (.A(_1788_),
    .X(_0474_));
 sky130_fd_sc_hd__or2_2 _3717_ (.A(_1131_),
    .B(_1305_),
    .X(_1789_));
 sky130_fd_sc_hd__mux2_1 _3718_ (.A0(_1775_),
    .A1(\tms1x00.RAM[82][0] ),
    .S(_1789_),
    .X(_1790_));
 sky130_fd_sc_hd__clkbuf_1 _3719_ (.A(_1790_),
    .X(_0475_));
 sky130_fd_sc_hd__mux2_1 _3720_ (.A0(_1778_),
    .A1(\tms1x00.RAM[82][1] ),
    .S(_1789_),
    .X(_1791_));
 sky130_fd_sc_hd__clkbuf_1 _3721_ (.A(_1791_),
    .X(_0476_));
 sky130_fd_sc_hd__mux2_1 _3722_ (.A0(_1780_),
    .A1(\tms1x00.RAM[82][2] ),
    .S(_1789_),
    .X(_1792_));
 sky130_fd_sc_hd__clkbuf_1 _3723_ (.A(_1792_),
    .X(_0477_));
 sky130_fd_sc_hd__mux2_1 _3724_ (.A0(_1782_),
    .A1(\tms1x00.RAM[82][3] ),
    .S(_1789_),
    .X(_1793_));
 sky130_fd_sc_hd__clkbuf_1 _3725_ (.A(_1793_),
    .X(_0478_));
 sky130_fd_sc_hd__or2_2 _3726_ (.A(_1131_),
    .B(_1182_),
    .X(_1794_));
 sky130_fd_sc_hd__mux2_1 _3727_ (.A0(_1775_),
    .A1(\tms1x00.RAM[81][0] ),
    .S(_1794_),
    .X(_1795_));
 sky130_fd_sc_hd__clkbuf_1 _3728_ (.A(_1795_),
    .X(_0479_));
 sky130_fd_sc_hd__mux2_1 _3729_ (.A0(_1778_),
    .A1(\tms1x00.RAM[81][1] ),
    .S(_1794_),
    .X(_1796_));
 sky130_fd_sc_hd__clkbuf_1 _3730_ (.A(_1796_),
    .X(_0480_));
 sky130_fd_sc_hd__mux2_1 _3731_ (.A0(_1780_),
    .A1(\tms1x00.RAM[81][2] ),
    .S(_1794_),
    .X(_1797_));
 sky130_fd_sc_hd__clkbuf_1 _3732_ (.A(_1797_),
    .X(_0481_));
 sky130_fd_sc_hd__mux2_1 _3733_ (.A0(_1782_),
    .A1(\tms1x00.RAM[81][3] ),
    .S(_1794_),
    .X(_1798_));
 sky130_fd_sc_hd__clkbuf_1 _3734_ (.A(_1798_),
    .X(_0482_));
 sky130_fd_sc_hd__mux2_1 _3735_ (.A0(_0616_),
    .A1(_0617_),
    .S(_0622_),
    .X(_1799_));
 sky130_fd_sc_hd__clkbuf_1 _3736_ (.A(_1799_),
    .X(_0483_));
 sky130_fd_sc_hd__mux2_1 _3737_ (.A0(_0624_),
    .A1(_0625_),
    .S(_0622_),
    .X(_1800_));
 sky130_fd_sc_hd__clkbuf_1 _3738_ (.A(_1800_),
    .X(_0484_));
 sky130_fd_sc_hd__mux2_1 _3739_ (.A0(_0627_),
    .A1(\tms1x00.ram_addr_buff[2] ),
    .S(_0622_),
    .X(_1801_));
 sky130_fd_sc_hd__clkbuf_1 _3740_ (.A(_1801_),
    .X(_0485_));
 sky130_fd_sc_hd__mux2_1 _3741_ (.A0(_0630_),
    .A1(\tms1x00.ram_addr_buff[3] ),
    .S(_0621_),
    .X(_1802_));
 sky130_fd_sc_hd__clkbuf_1 _3742_ (.A(_1802_),
    .X(_0486_));
 sky130_fd_sc_hd__mux2_1 _3743_ (.A0(\tms1x00.X[2] ),
    .A1(\tms1x00.ram_addr_buff[4] ),
    .S(_0621_),
    .X(_1803_));
 sky130_fd_sc_hd__clkbuf_1 _3744_ (.A(_1803_),
    .X(_0487_));
 sky130_fd_sc_hd__mux2_1 _3745_ (.A0(\tms1x00.X[0] ),
    .A1(\tms1x00.ram_addr_buff[5] ),
    .S(_0621_),
    .X(_1804_));
 sky130_fd_sc_hd__clkbuf_1 _3746_ (.A(_1804_),
    .X(_0488_));
 sky130_fd_sc_hd__mux2_1 _3747_ (.A0(\tms1x00.X[1] ),
    .A1(\tms1x00.ram_addr_buff[6] ),
    .S(_0621_),
    .X(_1805_));
 sky130_fd_sc_hd__clkbuf_1 _3748_ (.A(_1805_),
    .X(_0489_));
 sky130_fd_sc_hd__buf_2 _3749_ (.A(net16),
    .X(_1806_));
 sky130_fd_sc_hd__buf_2 _3750_ (.A(_1806_),
    .X(_1807_));
 sky130_fd_sc_hd__nor2_1 _3751_ (.A(net33),
    .B(_1807_),
    .Y(_0490_));
 sky130_fd_sc_hd__xnor2_1 _3752_ (.A(net33),
    .B(net34),
    .Y(_1808_));
 sky130_fd_sc_hd__and3b_1 _3753_ (.A_N(net34),
    .B(net33),
    .C(net35),
    .X(_1809_));
 sky130_fd_sc_hd__nor3_1 _3754_ (.A(_1807_),
    .B(_1808_),
    .C(_1809_),
    .Y(_0491_));
 sky130_fd_sc_hd__a21oi_1 _3755_ (.A1(_0619_),
    .A2(_0641_),
    .B1(_1807_),
    .Y(_0492_));
 sky130_fd_sc_hd__buf_2 _3756_ (.A(\tms1x00.rom_addr[1] ),
    .X(_1810_));
 sky130_fd_sc_hd__mux4_1 _3757_ (.A0(net5),
    .A1(net7),
    .A2(net8),
    .A3(net9),
    .S0(\tms1x00.rom_addr[0] ),
    .S1(_1810_),
    .X(_1811_));
 sky130_fd_sc_hd__mux2_1 _3758_ (.A0(\tms1x00.ins_in[0] ),
    .A1(_1811_),
    .S(_0620_),
    .X(_1812_));
 sky130_fd_sc_hd__or2_1 _3759_ (.A(_1807_),
    .B(_1812_),
    .X(_1813_));
 sky130_fd_sc_hd__clkbuf_1 _3760_ (.A(_1813_),
    .X(_0493_));
 sky130_fd_sc_hd__mux4_1 _3761_ (.A0(net7),
    .A1(net8),
    .A2(net9),
    .A3(net10),
    .S0(\tms1x00.rom_addr[0] ),
    .S1(_1810_),
    .X(_1814_));
 sky130_fd_sc_hd__mux2_1 _3762_ (.A0(\tms1x00.ins_in[1] ),
    .A1(_1814_),
    .S(_0620_),
    .X(_1815_));
 sky130_fd_sc_hd__or2_1 _3763_ (.A(_1807_),
    .B(_1815_),
    .X(_1816_));
 sky130_fd_sc_hd__clkbuf_1 _3764_ (.A(_1816_),
    .X(_0494_));
 sky130_fd_sc_hd__or2_1 _3765_ (.A(net34),
    .B(_0619_),
    .X(_1817_));
 sky130_fd_sc_hd__nor2_1 _3766_ (.A(_1806_),
    .B(_1817_),
    .Y(_1818_));
 sky130_fd_sc_hd__mux2_1 _3767_ (.A0(net8),
    .A1(net9),
    .S(\tms1x00.rom_addr[0] ),
    .X(_1819_));
 sky130_fd_sc_hd__or2_1 _3768_ (.A(_1810_),
    .B(_1819_),
    .X(_1820_));
 sky130_fd_sc_hd__mux2_1 _3769_ (.A0(net10),
    .A1(net11),
    .S(\tms1x00.rom_addr[0] ),
    .X(_1821_));
 sky130_fd_sc_hd__or2b_1 _3770_ (.A(_1821_),
    .B_N(_1810_),
    .X(_1822_));
 sky130_fd_sc_hd__nor2_2 _3771_ (.A(_1806_),
    .B(_0620_),
    .Y(_1823_));
 sky130_fd_sc_hd__a32o_1 _3772_ (.A1(_1818_),
    .A2(_1820_),
    .A3(_1822_),
    .B1(_1823_),
    .B2(\tms1x00.ins_in[2] ),
    .X(_0495_));
 sky130_fd_sc_hd__mux4_1 _3773_ (.A0(net9),
    .A1(net10),
    .A2(net11),
    .A3(net12),
    .S0(\tms1x00.rom_addr[0] ),
    .S1(_1810_),
    .X(_1824_));
 sky130_fd_sc_hd__or2_1 _3774_ (.A(_1817_),
    .B(_1824_),
    .X(_1825_));
 sky130_fd_sc_hd__clkbuf_4 _3775_ (.A(_0618_),
    .X(_1826_));
 sky130_fd_sc_hd__o211a_1 _3776_ (.A1(\tms1x00.ins_in[3] ),
    .A2(_0620_),
    .B1(_1825_),
    .C1(_1826_),
    .X(_0496_));
 sky130_fd_sc_hd__or2_1 _3777_ (.A(_1810_),
    .B(_1821_),
    .X(_1827_));
 sky130_fd_sc_hd__mux2_1 _3778_ (.A0(net12),
    .A1(net13),
    .S(\tms1x00.rom_addr[0] ),
    .X(_1828_));
 sky130_fd_sc_hd__or2b_1 _3779_ (.A(_1828_),
    .B_N(_1810_),
    .X(_1829_));
 sky130_fd_sc_hd__clkbuf_4 _3780_ (.A(\tms1x00.ins_in[4] ),
    .X(_1830_));
 sky130_fd_sc_hd__a32o_1 _3781_ (.A1(_1818_),
    .A2(_1827_),
    .A3(_1829_),
    .B1(_1823_),
    .B2(_1830_),
    .X(_0497_));
 sky130_fd_sc_hd__mux4_1 _3782_ (.A0(net11),
    .A1(net12),
    .A2(net13),
    .A3(net14),
    .S0(\tms1x00.rom_addr[0] ),
    .S1(\tms1x00.rom_addr[1] ),
    .X(_1831_));
 sky130_fd_sc_hd__mux2_1 _3783_ (.A0(_0926_),
    .A1(_1831_),
    .S(_0620_),
    .X(_1832_));
 sky130_fd_sc_hd__or2_1 _3784_ (.A(_1807_),
    .B(_1832_),
    .X(_1833_));
 sky130_fd_sc_hd__clkbuf_1 _3785_ (.A(_1833_),
    .X(_0498_));
 sky130_fd_sc_hd__mux4_1 _3786_ (.A0(net12),
    .A1(net13),
    .A2(net14),
    .A3(net15),
    .S0(\tms1x00.rom_addr[0] ),
    .S1(_1810_),
    .X(_1834_));
 sky130_fd_sc_hd__or2_1 _3787_ (.A(_1817_),
    .B(_1834_),
    .X(_1835_));
 sky130_fd_sc_hd__o211a_1 _3788_ (.A1(_0637_),
    .A2(_0620_),
    .B1(_1835_),
    .C1(_1826_),
    .X(_0499_));
 sky130_fd_sc_hd__mux4_1 _3789_ (.A0(net13),
    .A1(net14),
    .A2(net15),
    .A3(net6),
    .S0(\tms1x00.rom_addr[0] ),
    .S1(_1810_),
    .X(_1836_));
 sky130_fd_sc_hd__or2_1 _3790_ (.A(_1817_),
    .B(_1836_),
    .X(_1837_));
 sky130_fd_sc_hd__o211a_1 _3791_ (.A1(_0636_),
    .A2(_0620_),
    .B1(_1837_),
    .C1(_1826_),
    .X(_0500_));
 sky130_fd_sc_hd__or3b_1 _3792_ (.A(_0627_),
    .B(_0624_),
    .C_N(_0616_),
    .X(_1838_));
 sky130_fd_sc_hd__nor3b_1 _3793_ (.A(_0627_),
    .B(_0624_),
    .C_N(\tms1x00.Y[0] ),
    .Y(_1839_));
 sky130_fd_sc_hd__a31o_1 _3794_ (.A1(_0645_),
    .A2(_0650_),
    .A3(_1839_),
    .B1(net37),
    .X(_1840_));
 sky130_fd_sc_hd__o311a_1 _3795_ (.A1(_0630_),
    .A2(_0643_),
    .A3(_1838_),
    .B1(_1840_),
    .C1(_0652_),
    .X(_0501_));
 sky130_fd_sc_hd__or3b_1 _3796_ (.A(_0627_),
    .B(_0616_),
    .C_N(_0624_),
    .X(_1841_));
 sky130_fd_sc_hd__nor3b_1 _3797_ (.A(_0627_),
    .B(_0616_),
    .C_N(\tms1x00.Y[1] ),
    .Y(_1842_));
 sky130_fd_sc_hd__a31o_1 _3798_ (.A1(_0645_),
    .A2(_0650_),
    .A3(_1842_),
    .B1(net38),
    .X(_1843_));
 sky130_fd_sc_hd__buf_2 _3799_ (.A(_0618_),
    .X(_1844_));
 sky130_fd_sc_hd__o311a_1 _3800_ (.A1(_0630_),
    .A2(_0643_),
    .A3(_1841_),
    .B1(_1843_),
    .C1(_1844_),
    .X(_0502_));
 sky130_fd_sc_hd__and3b_1 _3801_ (.A_N(\tms1x00.Y[2] ),
    .B(\tms1x00.Y[1] ),
    .C(\tms1x00.Y[0] ),
    .X(_1845_));
 sky130_fd_sc_hd__a31o_1 _3802_ (.A1(_0645_),
    .A2(_0649_),
    .A3(_1845_),
    .B1(net39),
    .X(_1846_));
 sky130_fd_sc_hd__or3b_1 _3803_ (.A(\tms1x00.Y[3] ),
    .B(_0642_),
    .C_N(_1845_),
    .X(_1847_));
 sky130_fd_sc_hd__and3_1 _3804_ (.A(_1844_),
    .B(_1846_),
    .C(_1847_),
    .X(_1848_));
 sky130_fd_sc_hd__clkbuf_1 _3805_ (.A(_1848_),
    .X(_0503_));
 sky130_fd_sc_hd__or3b_1 _3806_ (.A(_0624_),
    .B(_0616_),
    .C_N(_0627_),
    .X(_1849_));
 sky130_fd_sc_hd__nor3b_1 _3807_ (.A(\tms1x00.Y[1] ),
    .B(\tms1x00.Y[0] ),
    .C_N(\tms1x00.Y[2] ),
    .Y(_1850_));
 sky130_fd_sc_hd__a31o_1 _3808_ (.A1(_0645_),
    .A2(_0650_),
    .A3(_1850_),
    .B1(net40),
    .X(_1851_));
 sky130_fd_sc_hd__o311a_1 _3809_ (.A1(_0630_),
    .A2(_0643_),
    .A3(_1849_),
    .B1(_1851_),
    .C1(_1844_),
    .X(_0504_));
 sky130_fd_sc_hd__and3b_1 _3810_ (.A_N(\tms1x00.Y[1] ),
    .B(\tms1x00.Y[0] ),
    .C(\tms1x00.Y[2] ),
    .X(_1852_));
 sky130_fd_sc_hd__a31o_1 _3811_ (.A1(_0645_),
    .A2(_0649_),
    .A3(_1852_),
    .B1(net41),
    .X(_1853_));
 sky130_fd_sc_hd__or3b_1 _3812_ (.A(\tms1x00.Y[3] ),
    .B(_0642_),
    .C_N(_1852_),
    .X(_1854_));
 sky130_fd_sc_hd__and3_1 _3813_ (.A(_1844_),
    .B(_1853_),
    .C(_1854_),
    .X(_1855_));
 sky130_fd_sc_hd__clkbuf_1 _3814_ (.A(_1855_),
    .X(_0505_));
 sky130_fd_sc_hd__and3b_1 _3815_ (.A_N(\tms1x00.Y[0] ),
    .B(\tms1x00.Y[1] ),
    .C(\tms1x00.Y[2] ),
    .X(_1856_));
 sky130_fd_sc_hd__a31o_1 _3816_ (.A1(_0644_),
    .A2(_0649_),
    .A3(_1856_),
    .B1(net42),
    .X(_1857_));
 sky130_fd_sc_hd__or3b_1 _3817_ (.A(\tms1x00.Y[3] ),
    .B(_0642_),
    .C_N(_1856_),
    .X(_1858_));
 sky130_fd_sc_hd__and3_1 _3818_ (.A(_1844_),
    .B(_1857_),
    .C(_1858_),
    .X(_1859_));
 sky130_fd_sc_hd__clkbuf_1 _3819_ (.A(_1859_),
    .X(_0506_));
 sky130_fd_sc_hd__and3_1 _3820_ (.A(\tms1x00.Y[2] ),
    .B(\tms1x00.Y[1] ),
    .C(\tms1x00.Y[0] ),
    .X(_1860_));
 sky130_fd_sc_hd__a31o_1 _3821_ (.A1(_0644_),
    .A2(_0649_),
    .A3(_1860_),
    .B1(net43),
    .X(_1861_));
 sky130_fd_sc_hd__or3b_1 _3822_ (.A(\tms1x00.Y[3] ),
    .B(_0642_),
    .C_N(_1860_),
    .X(_1862_));
 sky130_fd_sc_hd__and3_1 _3823_ (.A(_1844_),
    .B(_1861_),
    .C(_1862_),
    .X(_1863_));
 sky130_fd_sc_hd__clkbuf_1 _3824_ (.A(_1863_),
    .X(_0507_));
 sky130_fd_sc_hd__a31o_1 _3825_ (.A1(_0629_),
    .A2(_0646_),
    .A3(_0649_),
    .B1(net44),
    .X(_1864_));
 sky130_fd_sc_hd__o311a_1 _3826_ (.A1(_0645_),
    .A2(_0635_),
    .A3(_0643_),
    .B1(_1864_),
    .C1(_1844_),
    .X(_0508_));
 sky130_fd_sc_hd__a31o_1 _3827_ (.A1(_0629_),
    .A2(_0650_),
    .A3(_1839_),
    .B1(net45),
    .X(_1865_));
 sky130_fd_sc_hd__o311a_1 _3828_ (.A1(_0645_),
    .A2(_0643_),
    .A3(_1838_),
    .B1(_1865_),
    .C1(_1844_),
    .X(_0509_));
 sky130_fd_sc_hd__a31o_1 _3829_ (.A1(_0629_),
    .A2(_0650_),
    .A3(_1842_),
    .B1(net46),
    .X(_1866_));
 sky130_fd_sc_hd__o311a_1 _3830_ (.A1(_0645_),
    .A2(_0643_),
    .A3(_1841_),
    .B1(_1866_),
    .C1(_1844_),
    .X(_0510_));
 sky130_fd_sc_hd__a31o_1 _3831_ (.A1(_0629_),
    .A2(_0649_),
    .A3(_1845_),
    .B1(net47),
    .X(_1867_));
 sky130_fd_sc_hd__or3b_1 _3832_ (.A(_0644_),
    .B(_0642_),
    .C_N(_1845_),
    .X(_1868_));
 sky130_fd_sc_hd__and3_1 _3833_ (.A(_0618_),
    .B(_1867_),
    .C(_1868_),
    .X(_1869_));
 sky130_fd_sc_hd__clkbuf_1 _3834_ (.A(_1869_),
    .X(_0511_));
 sky130_fd_sc_hd__a31o_1 _3835_ (.A1(_0629_),
    .A2(_0650_),
    .A3(_1850_),
    .B1(net48),
    .X(_1870_));
 sky130_fd_sc_hd__o311a_1 _3836_ (.A1(_0645_),
    .A2(_0642_),
    .A3(_1849_),
    .B1(_1870_),
    .C1(_1844_),
    .X(_0512_));
 sky130_fd_sc_hd__nand2_1 _3837_ (.A(_0630_),
    .B(_1852_),
    .Y(_1871_));
 sky130_fd_sc_hd__a31o_1 _3838_ (.A1(_0629_),
    .A2(_0650_),
    .A3(_1852_),
    .B1(net49),
    .X(_1872_));
 sky130_fd_sc_hd__o211a_1 _3839_ (.A1(_0643_),
    .A2(_1871_),
    .B1(_1872_),
    .C1(_1826_),
    .X(_0513_));
 sky130_fd_sc_hd__nand2_1 _3840_ (.A(_0630_),
    .B(_1856_),
    .Y(_1873_));
 sky130_fd_sc_hd__a31o_1 _3841_ (.A1(_0629_),
    .A2(_0650_),
    .A3(_1856_),
    .B1(net50),
    .X(_1874_));
 sky130_fd_sc_hd__o211a_1 _3842_ (.A1(_0643_),
    .A2(_1873_),
    .B1(_1874_),
    .C1(_1826_),
    .X(_0514_));
 sky130_fd_sc_hd__nand2_1 _3843_ (.A(_0630_),
    .B(_1860_),
    .Y(_1875_));
 sky130_fd_sc_hd__a31o_1 _3844_ (.A1(_0629_),
    .A2(_0650_),
    .A3(_1860_),
    .B1(net51),
    .X(_1876_));
 sky130_fd_sc_hd__o211a_1 _3845_ (.A1(_0643_),
    .A2(_1875_),
    .B1(_1876_),
    .C1(_1826_),
    .X(_0515_));
 sky130_fd_sc_hd__nor2_1 _3846_ (.A(_0638_),
    .B(_0641_),
    .Y(_1877_));
 sky130_fd_sc_hd__and4b_1 _3847_ (.A_N(_0926_),
    .B(_1830_),
    .C(_1877_),
    .D(_0637_),
    .X(_1878_));
 sky130_fd_sc_hd__buf_2 _3848_ (.A(_1878_),
    .X(_1879_));
 sky130_fd_sc_hd__inv_2 _3849_ (.A(\tms1x00.A[0] ),
    .Y(_1880_));
 sky130_fd_sc_hd__o21ai_1 _3850_ (.A1(_0636_),
    .A2(_1880_),
    .B1(_1879_),
    .Y(_1881_));
 sky130_fd_sc_hd__o211a_1 _3851_ (.A1(net28),
    .A2(_1879_),
    .B1(_1881_),
    .C1(_1826_),
    .X(_0516_));
 sky130_fd_sc_hd__inv_2 _3852_ (.A(\tms1x00.A[1] ),
    .Y(_1882_));
 sky130_fd_sc_hd__o21ai_1 _3853_ (.A1(_0636_),
    .A2(_1882_),
    .B1(_1879_),
    .Y(_1883_));
 sky130_fd_sc_hd__o211a_1 _3854_ (.A1(net29),
    .A2(_1879_),
    .B1(_1883_),
    .C1(_1826_),
    .X(_0517_));
 sky130_fd_sc_hd__inv_2 _3855_ (.A(\tms1x00.A[2] ),
    .Y(_1884_));
 sky130_fd_sc_hd__o21ai_1 _3856_ (.A1(_0636_),
    .A2(_1884_),
    .B1(_1879_),
    .Y(_1885_));
 sky130_fd_sc_hd__o211a_1 _3857_ (.A1(net30),
    .A2(_1879_),
    .B1(_1885_),
    .C1(_1826_),
    .X(_0518_));
 sky130_fd_sc_hd__inv_2 _3858_ (.A(\tms1x00.A[3] ),
    .Y(_1886_));
 sky130_fd_sc_hd__o21ai_1 _3859_ (.A1(_0636_),
    .A2(_1886_),
    .B1(_1879_),
    .Y(_1887_));
 sky130_fd_sc_hd__o211a_1 _3860_ (.A1(net31),
    .A2(_1879_),
    .B1(_1887_),
    .C1(_1826_),
    .X(_0519_));
 sky130_fd_sc_hd__inv_2 _3861_ (.A(\tms1x00.status ),
    .Y(_1888_));
 sky130_fd_sc_hd__o21ai_1 _3862_ (.A1(_1888_),
    .A2(_0636_),
    .B1(_1879_),
    .Y(_1889_));
 sky130_fd_sc_hd__o211a_1 _3863_ (.A1(net32),
    .A2(_1879_),
    .B1(_1889_),
    .C1(_0652_),
    .X(_0520_));
 sky130_fd_sc_hd__inv_2 _3864_ (.A(\tms1x00.CL ),
    .Y(_1890_));
 sky130_fd_sc_hd__and3_1 _3865_ (.A(\tms1x00.status ),
    .B(\tms1x00.ins_in[0] ),
    .C(_1809_),
    .X(_1891_));
 sky130_fd_sc_hd__clkbuf_4 _3866_ (.A(_1891_),
    .X(_1892_));
 sky130_fd_sc_hd__nand2_2 _3867_ (.A(\tms1x00.ins_in[1] ),
    .B(_1892_),
    .Y(_1893_));
 sky130_fd_sc_hd__nor2_1 _3868_ (.A(_0640_),
    .B(_1124_),
    .Y(_1894_));
 sky130_fd_sc_hd__and3_1 _3869_ (.A(\tms1x00.CL ),
    .B(_1809_),
    .C(_1894_),
    .X(_1895_));
 sky130_fd_sc_hd__buf_2 _3870_ (.A(_1895_),
    .X(_1896_));
 sky130_fd_sc_hd__a211oi_1 _3871_ (.A1(_1890_),
    .A2(_1893_),
    .B1(_1896_),
    .C1(_1807_),
    .Y(_0521_));
 sky130_fd_sc_hd__or3_1 _3872_ (.A(\tms1x00.status ),
    .B(_1806_),
    .C(_1809_),
    .X(_1897_));
 sky130_fd_sc_hd__clkbuf_1 _3873_ (.A(_1897_),
    .X(_0522_));
 sky130_fd_sc_hd__mux2_1 _3874_ (.A0(\tms1x00.PA[0] ),
    .A1(\tms1x00.PB[0] ),
    .S(_1893_),
    .X(_1898_));
 sky130_fd_sc_hd__inv_2 _3875_ (.A(_0641_),
    .Y(_1899_));
 sky130_fd_sc_hd__and3b_1 _3876_ (.A_N(\tms1x00.ins_in[2] ),
    .B(_0813_),
    .C(\tms1x00.ins_in[3] ),
    .X(_1900_));
 sky130_fd_sc_hd__nand2_2 _3877_ (.A(_1899_),
    .B(_1900_),
    .Y(_1901_));
 sky130_fd_sc_hd__mux2_1 _3878_ (.A0(_1830_),
    .A1(_1898_),
    .S(_1901_),
    .X(_1902_));
 sky130_fd_sc_hd__or2_1 _3879_ (.A(_1807_),
    .B(_1902_),
    .X(_1903_));
 sky130_fd_sc_hd__clkbuf_1 _3880_ (.A(_1903_),
    .X(_0523_));
 sky130_fd_sc_hd__mux2_1 _3881_ (.A0(\tms1x00.PA[1] ),
    .A1(\tms1x00.PB[1] ),
    .S(_1893_),
    .X(_1904_));
 sky130_fd_sc_hd__mux2_1 _3882_ (.A0(_0926_),
    .A1(_1904_),
    .S(_1901_),
    .X(_1905_));
 sky130_fd_sc_hd__or2_1 _3883_ (.A(_1807_),
    .B(_1905_),
    .X(_1906_));
 sky130_fd_sc_hd__clkbuf_1 _3884_ (.A(_1906_),
    .X(_0524_));
 sky130_fd_sc_hd__mux2_1 _3885_ (.A0(\tms1x00.PA[2] ),
    .A1(\tms1x00.PB[2] ),
    .S(_1893_),
    .X(_1907_));
 sky130_fd_sc_hd__mux2_1 _3886_ (.A0(_0637_),
    .A1(_1907_),
    .S(_1901_),
    .X(_1908_));
 sky130_fd_sc_hd__or2_1 _3887_ (.A(_1806_),
    .B(_1908_),
    .X(_1909_));
 sky130_fd_sc_hd__clkbuf_1 _3888_ (.A(_1909_),
    .X(_0525_));
 sky130_fd_sc_hd__mux2_1 _3889_ (.A0(\tms1x00.PA[3] ),
    .A1(\tms1x00.PB[3] ),
    .S(_1893_),
    .X(_1910_));
 sky130_fd_sc_hd__mux2_1 _3890_ (.A0(_0636_),
    .A1(_1910_),
    .S(_1901_),
    .X(_1911_));
 sky130_fd_sc_hd__or2_1 _3891_ (.A(_1806_),
    .B(_1911_),
    .X(_1912_));
 sky130_fd_sc_hd__clkbuf_1 _3892_ (.A(_1912_),
    .X(_0526_));
 sky130_fd_sc_hd__and4_2 _3893_ (.A(_1890_),
    .B(\tms1x00.ins_in[1] ),
    .C(_0618_),
    .D(_1892_),
    .X(_1913_));
 sky130_fd_sc_hd__mux2_1 _3894_ (.A0(\tms1x00.SR[0] ),
    .A1(\tms1x00.PC[0] ),
    .S(_1913_),
    .X(_1914_));
 sky130_fd_sc_hd__clkbuf_1 _3895_ (.A(_1914_),
    .X(_0527_));
 sky130_fd_sc_hd__mux2_1 _3896_ (.A0(\tms1x00.SR[1] ),
    .A1(\tms1x00.PC[1] ),
    .S(_1913_),
    .X(_1915_));
 sky130_fd_sc_hd__clkbuf_1 _3897_ (.A(_1915_),
    .X(_0528_));
 sky130_fd_sc_hd__mux2_1 _3898_ (.A0(\tms1x00.SR[2] ),
    .A1(\tms1x00.PC[2] ),
    .S(_1913_),
    .X(_1916_));
 sky130_fd_sc_hd__clkbuf_1 _3899_ (.A(_1916_),
    .X(_0529_));
 sky130_fd_sc_hd__mux2_1 _3900_ (.A0(\tms1x00.SR[3] ),
    .A1(\tms1x00.PC[3] ),
    .S(_1913_),
    .X(_1917_));
 sky130_fd_sc_hd__clkbuf_1 _3901_ (.A(_1917_),
    .X(_0530_));
 sky130_fd_sc_hd__mux2_1 _3902_ (.A0(\tms1x00.SR[4] ),
    .A1(\tms1x00.PC[4] ),
    .S(_1913_),
    .X(_1918_));
 sky130_fd_sc_hd__clkbuf_1 _3903_ (.A(_1918_),
    .X(_0531_));
 sky130_fd_sc_hd__mux2_1 _3904_ (.A0(\tms1x00.SR[5] ),
    .A1(\tms1x00.PC[5] ),
    .S(_1913_),
    .X(_1919_));
 sky130_fd_sc_hd__clkbuf_1 _3905_ (.A(_1919_),
    .X(_0532_));
 sky130_fd_sc_hd__and3_1 _3906_ (.A(\tms1x00.status ),
    .B(_1890_),
    .C(\tms1x00.ins_in[0] ),
    .X(_1920_));
 sky130_fd_sc_hd__o21a_1 _3907_ (.A1(_1894_),
    .A2(_1920_),
    .B1(_1809_),
    .X(_1921_));
 sky130_fd_sc_hd__mux2_1 _3908_ (.A0(\tms1x00.PA[0] ),
    .A1(\tms1x00.PB[0] ),
    .S(_1921_),
    .X(_1922_));
 sky130_fd_sc_hd__or2_1 _3909_ (.A(_1806_),
    .B(_1922_),
    .X(_1923_));
 sky130_fd_sc_hd__clkbuf_1 _3910_ (.A(_1923_),
    .X(_0533_));
 sky130_fd_sc_hd__mux2_1 _3911_ (.A0(\tms1x00.PA[1] ),
    .A1(\tms1x00.PB[1] ),
    .S(_1921_),
    .X(_1924_));
 sky130_fd_sc_hd__or2_1 _3912_ (.A(_1806_),
    .B(_1924_),
    .X(_1925_));
 sky130_fd_sc_hd__clkbuf_1 _3913_ (.A(_1925_),
    .X(_0534_));
 sky130_fd_sc_hd__mux2_1 _3914_ (.A0(\tms1x00.PA[2] ),
    .A1(\tms1x00.PB[2] ),
    .S(_1921_),
    .X(_1926_));
 sky130_fd_sc_hd__or2_1 _3915_ (.A(_1806_),
    .B(_1926_),
    .X(_1927_));
 sky130_fd_sc_hd__clkbuf_1 _3916_ (.A(_1927_),
    .X(_0535_));
 sky130_fd_sc_hd__mux2_1 _3917_ (.A0(\tms1x00.PA[3] ),
    .A1(\tms1x00.PB[3] ),
    .S(_1921_),
    .X(_1928_));
 sky130_fd_sc_hd__or2_1 _3918_ (.A(_1806_),
    .B(_1928_),
    .X(_1929_));
 sky130_fd_sc_hd__clkbuf_1 _3919_ (.A(_1929_),
    .X(_0536_));
 sky130_fd_sc_hd__inv_2 _3920_ (.A(_1892_),
    .Y(_1930_));
 sky130_fd_sc_hd__inv_2 _3921_ (.A(_1896_),
    .Y(_1931_));
 sky130_fd_sc_hd__or3_1 _3922_ (.A(\tms1x00.PC[0] ),
    .B(_1892_),
    .C(_1896_),
    .X(_1932_));
 sky130_fd_sc_hd__o221a_1 _3923_ (.A1(\tms1x00.ins_in[2] ),
    .A2(_1930_),
    .B1(_1931_),
    .B2(\tms1x00.SR[0] ),
    .C1(_1932_),
    .X(_1933_));
 sky130_fd_sc_hd__a21oi_1 _3924_ (.A1(_0620_),
    .A2(_1933_),
    .B1(_1807_),
    .Y(_1934_));
 sky130_fd_sc_hd__o21a_1 _3925_ (.A1(_0620_),
    .A2(_1933_),
    .B1(_1934_),
    .X(_0537_));
 sky130_fd_sc_hd__nor2_1 _3926_ (.A(_1892_),
    .B(_1896_),
    .Y(_1935_));
 sky130_fd_sc_hd__and2_1 _3927_ (.A(\tms1x00.PC[1] ),
    .B(_1935_),
    .X(_1936_));
 sky130_fd_sc_hd__a22o_1 _3928_ (.A1(\tms1x00.ins_in[3] ),
    .A2(_1892_),
    .B1(_1896_),
    .B2(\tms1x00.SR[1] ),
    .X(_1937_));
 sky130_fd_sc_hd__o21a_1 _3929_ (.A1(_1936_),
    .A2(_1937_),
    .B1(_1823_),
    .X(_0538_));
 sky130_fd_sc_hd__a22o_1 _3930_ (.A1(_1830_),
    .A2(_1892_),
    .B1(_1896_),
    .B2(\tms1x00.SR[2] ),
    .X(_1938_));
 sky130_fd_sc_hd__a21o_1 _3931_ (.A1(\tms1x00.PC[2] ),
    .A2(_1935_),
    .B1(_1938_),
    .X(_1939_));
 sky130_fd_sc_hd__and2_1 _3932_ (.A(_1823_),
    .B(_1939_),
    .X(_1940_));
 sky130_fd_sc_hd__clkbuf_1 _3933_ (.A(_1940_),
    .X(_0539_));
 sky130_fd_sc_hd__and2_1 _3934_ (.A(\tms1x00.PC[3] ),
    .B(_1935_),
    .X(_1941_));
 sky130_fd_sc_hd__a22o_1 _3935_ (.A1(_0926_),
    .A2(_1892_),
    .B1(_1896_),
    .B2(\tms1x00.SR[3] ),
    .X(_1942_));
 sky130_fd_sc_hd__o21a_1 _3936_ (.A1(_1941_),
    .A2(_1942_),
    .B1(_1823_),
    .X(_0540_));
 sky130_fd_sc_hd__and2_1 _3937_ (.A(\tms1x00.PC[4] ),
    .B(_1935_),
    .X(_1943_));
 sky130_fd_sc_hd__a22o_1 _3938_ (.A1(_0637_),
    .A2(_1892_),
    .B1(_1896_),
    .B2(\tms1x00.SR[4] ),
    .X(_1944_));
 sky130_fd_sc_hd__o21a_1 _3939_ (.A1(_1943_),
    .A2(_1944_),
    .B1(_1823_),
    .X(_0541_));
 sky130_fd_sc_hd__and2_1 _3940_ (.A(\tms1x00.PC[5] ),
    .B(_1935_),
    .X(_1945_));
 sky130_fd_sc_hd__a22o_1 _3941_ (.A1(_0636_),
    .A2(_1892_),
    .B1(_1896_),
    .B2(\tms1x00.SR[5] ),
    .X(_1946_));
 sky130_fd_sc_hd__o21a_1 _3942_ (.A1(_1945_),
    .A2(_1946_),
    .B1(_1823_),
    .X(_0542_));
 sky130_fd_sc_hd__or3_1 _3943_ (.A(net35),
    .B(net34),
    .C(net16),
    .X(_1947_));
 sky130_fd_sc_hd__nor2_2 _3944_ (.A(net33),
    .B(_1947_),
    .Y(_1948_));
 sky130_fd_sc_hd__nor2_1 _3945_ (.A(_0757_),
    .B(_0811_),
    .Y(_1949_));
 sky130_fd_sc_hd__nand2_1 _3946_ (.A(_0653_),
    .B(_1900_),
    .Y(_1950_));
 sky130_fd_sc_hd__nand2_1 _3947_ (.A(\tms1x00.ins_in[1] ),
    .B(\tms1x00.ins_in[0] ),
    .Y(_1951_));
 sky130_fd_sc_hd__or2_1 _3948_ (.A(_0654_),
    .B(_1951_),
    .X(_1952_));
 sky130_fd_sc_hd__nor4_1 _3949_ (.A(\tms1x00.ins_in[7] ),
    .B(_0637_),
    .C(\tms1x00.ins_in[5] ),
    .D(_1830_),
    .Y(_1953_));
 sky130_fd_sc_hd__and2_1 _3950_ (.A(\tms1x00.ins_in[3] ),
    .B(_1953_),
    .X(_1954_));
 sky130_fd_sc_hd__or2_1 _3951_ (.A(net33),
    .B(_1947_),
    .X(_1955_));
 sky130_fd_sc_hd__a221o_1 _3952_ (.A1(_1830_),
    .A2(_0924_),
    .B1(_1954_),
    .B2(\tms1x00.K_latch[0] ),
    .C1(_1955_),
    .X(_1956_));
 sky130_fd_sc_hd__a21o_1 _3953_ (.A1(_0616_),
    .A2(_1952_),
    .B1(_1956_),
    .X(_1957_));
 sky130_fd_sc_hd__a21o_1 _3954_ (.A1(_1949_),
    .A2(_1950_),
    .B1(_1957_),
    .X(_1958_));
 sky130_fd_sc_hd__o21a_1 _3955_ (.A1(\tms1x00.P[0] ),
    .A2(_1948_),
    .B1(_1958_),
    .X(_0543_));
 sky130_fd_sc_hd__nor3b_1 _3956_ (.A(_0876_),
    .B(_0923_),
    .C_N(_1950_),
    .Y(_1959_));
 sky130_fd_sc_hd__a221o_1 _3957_ (.A1(_0926_),
    .A2(_0924_),
    .B1(_1954_),
    .B2(\tms1x00.K_latch[1] ),
    .C1(_1955_),
    .X(_1960_));
 sky130_fd_sc_hd__a21o_1 _3958_ (.A1(_0624_),
    .A2(_1952_),
    .B1(_1960_),
    .X(_1961_));
 sky130_fd_sc_hd__o22a_1 _3959_ (.A1(\tms1x00.P[1] ),
    .A2(_1948_),
    .B1(_1959_),
    .B2(_1961_),
    .X(_0544_));
 sky130_fd_sc_hd__nor2_1 _3960_ (.A(_0978_),
    .B(_1025_),
    .Y(_1962_));
 sky130_fd_sc_hd__a31o_1 _3961_ (.A1(\tms1x00.ins_in[3] ),
    .A2(\tms1x00.K_latch[2] ),
    .A3(_1953_),
    .B1(_0924_),
    .X(_1963_));
 sky130_fd_sc_hd__a221o_1 _3962_ (.A1(_1962_),
    .A2(_1950_),
    .B1(_1952_),
    .B2(\tms1x00.Y[2] ),
    .C1(_1963_),
    .X(_1964_));
 sky130_fd_sc_hd__mux2_1 _3963_ (.A0(\tms1x00.P[2] ),
    .A1(_1964_),
    .S(_1948_),
    .X(_1965_));
 sky130_fd_sc_hd__clkbuf_1 _3964_ (.A(_1965_),
    .X(_0545_));
 sky130_fd_sc_hd__and2_1 _3965_ (.A(_1123_),
    .B(_1950_),
    .X(_1966_));
 sky130_fd_sc_hd__a221o_1 _3966_ (.A1(_0629_),
    .A2(_1952_),
    .B1(_1954_),
    .B2(\tms1x00.K_latch[3] ),
    .C1(_1955_),
    .X(_1967_));
 sky130_fd_sc_hd__o22a_1 _3967_ (.A1(\tms1x00.P[3] ),
    .A2(_1948_),
    .B1(_1966_),
    .B2(_1967_),
    .X(_0546_));
 sky130_fd_sc_hd__nor3b_4 _3968_ (.A(_1830_),
    .B(_0648_),
    .C_N(_0926_),
    .Y(_1968_));
 sky130_fd_sc_hd__o31a_1 _3969_ (.A1(\tms1x00.ins_in[5] ),
    .A2(_1830_),
    .A3(_0647_),
    .B1(\tms1x00.N[0] ),
    .X(_1969_));
 sky130_fd_sc_hd__or4_1 _3970_ (.A(\tms1x00.ins_in[5] ),
    .B(\tms1x00.ins_in[4] ),
    .C(\tms1x00.N[0] ),
    .D(_0647_),
    .X(_1970_));
 sky130_fd_sc_hd__and2b_1 _3971_ (.A_N(_1969_),
    .B(_1970_),
    .X(_1971_));
 sky130_fd_sc_hd__xnor2_1 _3972_ (.A(\tms1x00.P[0] ),
    .B(_1971_),
    .Y(_1972_));
 sky130_fd_sc_hd__nand2_1 _3973_ (.A(_1968_),
    .B(_1972_),
    .Y(_1973_));
 sky130_fd_sc_hd__o211a_1 _3974_ (.A1(_0616_),
    .A2(_1968_),
    .B1(_1973_),
    .C1(_0652_),
    .X(_0547_));
 sky130_fd_sc_hd__nor2_1 _3975_ (.A(\tms1x00.P[1] ),
    .B(\tms1x00.N[1] ),
    .Y(_1974_));
 sky130_fd_sc_hd__and2_1 _3976_ (.A(\tms1x00.P[1] ),
    .B(\tms1x00.N[1] ),
    .X(_1975_));
 sky130_fd_sc_hd__or2_1 _3977_ (.A(_1974_),
    .B(_1975_),
    .X(_1976_));
 sky130_fd_sc_hd__a21oi_1 _3978_ (.A1(\tms1x00.P[0] ),
    .A2(_1970_),
    .B1(_1969_),
    .Y(_1977_));
 sky130_fd_sc_hd__xnor2_1 _3979_ (.A(_1976_),
    .B(_1977_),
    .Y(_1978_));
 sky130_fd_sc_hd__nand2_1 _3980_ (.A(_1968_),
    .B(_1978_),
    .Y(_1979_));
 sky130_fd_sc_hd__o211a_1 _3981_ (.A1(_0624_),
    .A2(_1968_),
    .B1(_1979_),
    .C1(_0652_),
    .X(_0548_));
 sky130_fd_sc_hd__or2_1 _3982_ (.A(\tms1x00.P[2] ),
    .B(\tms1x00.N[2] ),
    .X(_1980_));
 sky130_fd_sc_hd__nand2_1 _3983_ (.A(\tms1x00.P[2] ),
    .B(\tms1x00.N[2] ),
    .Y(_1981_));
 sky130_fd_sc_hd__nand2_1 _3984_ (.A(_1980_),
    .B(_1981_),
    .Y(_1982_));
 sky130_fd_sc_hd__o21ba_1 _3985_ (.A1(_1974_),
    .A2(_1977_),
    .B1_N(_1975_),
    .X(_1983_));
 sky130_fd_sc_hd__xnor2_1 _3986_ (.A(_1982_),
    .B(_1983_),
    .Y(_1984_));
 sky130_fd_sc_hd__nand2_1 _3987_ (.A(_1968_),
    .B(_1984_),
    .Y(_1985_));
 sky130_fd_sc_hd__o211a_1 _3988_ (.A1(_0627_),
    .A2(_1968_),
    .B1(_1985_),
    .C1(_0652_),
    .X(_0549_));
 sky130_fd_sc_hd__o21a_1 _3989_ (.A1(_1982_),
    .A2(_1983_),
    .B1(_1981_),
    .X(_1986_));
 sky130_fd_sc_hd__xnor2_1 _3990_ (.A(\tms1x00.P[3] ),
    .B(\tms1x00.N[3] ),
    .Y(_1987_));
 sky130_fd_sc_hd__xnor2_1 _3991_ (.A(_1986_),
    .B(_1987_),
    .Y(_1988_));
 sky130_fd_sc_hd__nand2_1 _3992_ (.A(_1968_),
    .B(_1988_),
    .Y(_1989_));
 sky130_fd_sc_hd__o211a_1 _3993_ (.A1(_0630_),
    .A2(_1968_),
    .B1(_1989_),
    .C1(_0652_),
    .X(_0550_));
 sky130_fd_sc_hd__and3_1 _3994_ (.A(_0926_),
    .B(_1830_),
    .C(_0814_),
    .X(_1990_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _3995_ (.A(_1990_),
    .X(_1991_));
 sky130_fd_sc_hd__a22o_1 _3996_ (.A1(_1877_),
    .A2(_1953_),
    .B1(_1991_),
    .B2(_1899_),
    .X(_1992_));
 sky130_fd_sc_hd__nand2_1 _3997_ (.A(_0637_),
    .B(_1991_),
    .Y(_1993_));
 sky130_fd_sc_hd__o211ai_1 _3998_ (.A1(\tms1x00.X[0] ),
    .A2(_1991_),
    .B1(_1992_),
    .C1(_1993_),
    .Y(_1994_));
 sky130_fd_sc_hd__o211a_1 _3999_ (.A1(\tms1x00.X[0] ),
    .A2(_1992_),
    .B1(_1994_),
    .C1(_0652_),
    .X(_0551_));
 sky130_fd_sc_hd__nand2_1 _4000_ (.A(_0636_),
    .B(_1991_),
    .Y(_1995_));
 sky130_fd_sc_hd__o211ai_1 _4001_ (.A1(\tms1x00.X[1] ),
    .A2(_1991_),
    .B1(_1992_),
    .C1(_1995_),
    .Y(_1996_));
 sky130_fd_sc_hd__o211a_1 _4002_ (.A1(\tms1x00.X[1] ),
    .A2(_1992_),
    .B1(_1996_),
    .C1(_0652_),
    .X(_0552_));
 sky130_fd_sc_hd__o21ai_1 _4003_ (.A1(\tms1x00.X[2] ),
    .A2(_0926_),
    .B1(_1992_),
    .Y(_1997_));
 sky130_fd_sc_hd__o211a_1 _4004_ (.A1(\tms1x00.X[2] ),
    .A2(_1992_),
    .B1(_1997_),
    .C1(_0652_),
    .X(_0553_));
 sky130_fd_sc_hd__or2_1 _4005_ (.A(\tms1x00.N[0] ),
    .B(_1948_),
    .X(_1998_));
 sky130_fd_sc_hd__clkbuf_1 _4006_ (.A(_1998_),
    .X(_0554_));
 sky130_fd_sc_hd__or2_1 _4007_ (.A(\tms1x00.N[1] ),
    .B(_1948_),
    .X(_1999_));
 sky130_fd_sc_hd__clkbuf_1 _4008_ (.A(_1999_),
    .X(_0555_));
 sky130_fd_sc_hd__or2_1 _4009_ (.A(\tms1x00.N[2] ),
    .B(_1948_),
    .X(_2000_));
 sky130_fd_sc_hd__clkbuf_1 _4010_ (.A(_2000_),
    .X(_0556_));
 sky130_fd_sc_hd__or2_1 _4011_ (.A(\tms1x00.N[3] ),
    .B(_1948_),
    .X(_2001_));
 sky130_fd_sc_hd__clkbuf_1 _4012_ (.A(_2001_),
    .X(_0557_));
 sky130_fd_sc_hd__or4b_1 _4013_ (.A(_0926_),
    .B(net16),
    .C(_0648_),
    .D_N(_1830_),
    .X(_2002_));
 sky130_fd_sc_hd__buf_2 _4014_ (.A(_2002_),
    .X(_2003_));
 sky130_fd_sc_hd__nand2_1 _4015_ (.A(\tms1x00.A[0] ),
    .B(_2003_),
    .Y(_2004_));
 sky130_fd_sc_hd__o21ai_1 _4016_ (.A1(_1972_),
    .A2(_2003_),
    .B1(_2004_),
    .Y(_0558_));
 sky130_fd_sc_hd__nand2_1 _4017_ (.A(\tms1x00.A[1] ),
    .B(_2003_),
    .Y(_2005_));
 sky130_fd_sc_hd__o21ai_1 _4018_ (.A1(_1978_),
    .A2(_2003_),
    .B1(_2005_),
    .Y(_0559_));
 sky130_fd_sc_hd__nand2_1 _4019_ (.A(\tms1x00.A[2] ),
    .B(_2003_),
    .Y(_2006_));
 sky130_fd_sc_hd__o21ai_1 _4020_ (.A1(_1984_),
    .A2(_2003_),
    .B1(_2006_),
    .Y(_0560_));
 sky130_fd_sc_hd__nand2_1 _4021_ (.A(\tms1x00.A[3] ),
    .B(_2003_),
    .Y(_2007_));
 sky130_fd_sc_hd__o21ai_1 _4022_ (.A1(_1988_),
    .A2(_2003_),
    .B1(_2007_),
    .Y(_0561_));
 sky130_fd_sc_hd__or2_2 _4023_ (.A(_1154_),
    .B(_1232_),
    .X(_2008_));
 sky130_fd_sc_hd__mux2_1 _4024_ (.A0(_1775_),
    .A1(\tms1x00.RAM[13][0] ),
    .S(_2008_),
    .X(_2009_));
 sky130_fd_sc_hd__clkbuf_1 _4025_ (.A(_2009_),
    .X(_0562_));
 sky130_fd_sc_hd__mux2_1 _4026_ (.A0(_1778_),
    .A1(\tms1x00.RAM[13][1] ),
    .S(_2008_),
    .X(_2010_));
 sky130_fd_sc_hd__clkbuf_1 _4027_ (.A(_2010_),
    .X(_0563_));
 sky130_fd_sc_hd__mux2_1 _4028_ (.A0(_1780_),
    .A1(\tms1x00.RAM[13][2] ),
    .S(_2008_),
    .X(_2011_));
 sky130_fd_sc_hd__clkbuf_1 _4029_ (.A(_2011_),
    .X(_0564_));
 sky130_fd_sc_hd__mux2_1 _4030_ (.A0(_1782_),
    .A1(\tms1x00.RAM[13][3] ),
    .S(_2008_),
    .X(_2012_));
 sky130_fd_sc_hd__clkbuf_1 _4031_ (.A(_2012_),
    .X(_0565_));
 sky130_fd_sc_hd__or2_2 _4032_ (.A(_1442_),
    .B(_1305_),
    .X(_2013_));
 sky130_fd_sc_hd__mux2_1 _4033_ (.A0(_1775_),
    .A1(\tms1x00.RAM[18][0] ),
    .S(_2013_),
    .X(_2014_));
 sky130_fd_sc_hd__clkbuf_1 _4034_ (.A(_2014_),
    .X(_0566_));
 sky130_fd_sc_hd__mux2_1 _4035_ (.A0(_1778_),
    .A1(\tms1x00.RAM[18][1] ),
    .S(_2013_),
    .X(_2015_));
 sky130_fd_sc_hd__clkbuf_1 _4036_ (.A(_2015_),
    .X(_0567_));
 sky130_fd_sc_hd__mux2_1 _4037_ (.A0(_1780_),
    .A1(\tms1x00.RAM[18][2] ),
    .S(_2013_),
    .X(_2016_));
 sky130_fd_sc_hd__clkbuf_1 _4038_ (.A(_2016_),
    .X(_0568_));
 sky130_fd_sc_hd__mux2_1 _4039_ (.A0(_1782_),
    .A1(\tms1x00.RAM[18][3] ),
    .S(_2013_),
    .X(_2017_));
 sky130_fd_sc_hd__clkbuf_1 _4040_ (.A(_2017_),
    .X(_0569_));
 sky130_fd_sc_hd__nor2_2 _4041_ (.A(_1247_),
    .B(_1497_),
    .Y(_2018_));
 sky130_fd_sc_hd__mux2_1 _4042_ (.A0(\tms1x00.RAM[39][0] ),
    .A1(_1265_),
    .S(_2018_),
    .X(_2019_));
 sky130_fd_sc_hd__clkbuf_1 _4043_ (.A(_2019_),
    .X(_0570_));
 sky130_fd_sc_hd__mux2_1 _4044_ (.A0(\tms1x00.RAM[39][1] ),
    .A1(_1269_),
    .S(_2018_),
    .X(_2020_));
 sky130_fd_sc_hd__clkbuf_1 _4045_ (.A(_2020_),
    .X(_0571_));
 sky130_fd_sc_hd__mux2_1 _4046_ (.A0(\tms1x00.RAM[39][2] ),
    .A1(_1272_),
    .S(_2018_),
    .X(_2021_));
 sky130_fd_sc_hd__clkbuf_1 _4047_ (.A(_2021_),
    .X(_0572_));
 sky130_fd_sc_hd__mux2_1 _4048_ (.A0(\tms1x00.RAM[39][3] ),
    .A1(_1275_),
    .S(_2018_),
    .X(_2022_));
 sky130_fd_sc_hd__clkbuf_1 _4049_ (.A(_2022_),
    .X(_0573_));
 sky130_fd_sc_hd__or2_2 _4050_ (.A(_1199_),
    .B(_1232_),
    .X(_2023_));
 sky130_fd_sc_hd__mux2_1 _4051_ (.A0(_1775_),
    .A1(\tms1x00.RAM[14][0] ),
    .S(_2023_),
    .X(_2024_));
 sky130_fd_sc_hd__clkbuf_1 _4052_ (.A(_2024_),
    .X(_0574_));
 sky130_fd_sc_hd__mux2_1 _4053_ (.A0(_1778_),
    .A1(\tms1x00.RAM[14][1] ),
    .S(_2023_),
    .X(_2025_));
 sky130_fd_sc_hd__clkbuf_1 _4054_ (.A(_2025_),
    .X(_0575_));
 sky130_fd_sc_hd__mux2_1 _4055_ (.A0(_1780_),
    .A1(\tms1x00.RAM[14][2] ),
    .S(_2023_),
    .X(_2026_));
 sky130_fd_sc_hd__clkbuf_1 _4056_ (.A(_2026_),
    .X(_0576_));
 sky130_fd_sc_hd__mux2_1 _4057_ (.A0(_1782_),
    .A1(\tms1x00.RAM[14][3] ),
    .S(_2023_),
    .X(_2027_));
 sky130_fd_sc_hd__clkbuf_1 _4058_ (.A(_2027_),
    .X(_0577_));
 sky130_fd_sc_hd__or2_2 _4059_ (.A(_1182_),
    .B(_1188_),
    .X(_2028_));
 sky130_fd_sc_hd__mux2_1 _4060_ (.A0(_1775_),
    .A1(\tms1x00.RAM[17][0] ),
    .S(_2028_),
    .X(_2029_));
 sky130_fd_sc_hd__clkbuf_1 _4061_ (.A(_2029_),
    .X(_0578_));
 sky130_fd_sc_hd__mux2_1 _4062_ (.A0(_1778_),
    .A1(\tms1x00.RAM[17][1] ),
    .S(_2028_),
    .X(_2030_));
 sky130_fd_sc_hd__clkbuf_1 _4063_ (.A(_2030_),
    .X(_0579_));
 sky130_fd_sc_hd__mux2_1 _4064_ (.A0(_1780_),
    .A1(\tms1x00.RAM[17][2] ),
    .S(_2028_),
    .X(_2031_));
 sky130_fd_sc_hd__clkbuf_1 _4065_ (.A(_2031_),
    .X(_0580_));
 sky130_fd_sc_hd__mux2_1 _4066_ (.A0(_1782_),
    .A1(\tms1x00.RAM[17][3] ),
    .S(_2028_),
    .X(_2032_));
 sky130_fd_sc_hd__clkbuf_1 _4067_ (.A(_2032_),
    .X(_0581_));
 sky130_fd_sc_hd__or2_2 _4068_ (.A(_1154_),
    .B(_1188_),
    .X(_2033_));
 sky130_fd_sc_hd__mux2_1 _4069_ (.A0(_1775_),
    .A1(\tms1x00.RAM[29][0] ),
    .S(_2033_),
    .X(_2034_));
 sky130_fd_sc_hd__clkbuf_1 _4070_ (.A(_2034_),
    .X(_0582_));
 sky130_fd_sc_hd__mux2_1 _4071_ (.A0(_1778_),
    .A1(\tms1x00.RAM[29][1] ),
    .S(_2033_),
    .X(_2035_));
 sky130_fd_sc_hd__clkbuf_1 _4072_ (.A(_2035_),
    .X(_0583_));
 sky130_fd_sc_hd__mux2_1 _4073_ (.A0(_1780_),
    .A1(\tms1x00.RAM[29][2] ),
    .S(_2033_),
    .X(_2036_));
 sky130_fd_sc_hd__clkbuf_1 _4074_ (.A(_2036_),
    .X(_0584_));
 sky130_fd_sc_hd__mux2_1 _4075_ (.A0(_1782_),
    .A1(\tms1x00.RAM[29][3] ),
    .S(_2033_),
    .X(_2037_));
 sky130_fd_sc_hd__clkbuf_1 _4076_ (.A(_2037_),
    .X(_0585_));
 sky130_fd_sc_hd__or2_2 _4077_ (.A(_1188_),
    .B(_1299_),
    .X(_2038_));
 sky130_fd_sc_hd__mux2_1 _4078_ (.A0(_1775_),
    .A1(\tms1x00.RAM[16][0] ),
    .S(_2038_),
    .X(_2039_));
 sky130_fd_sc_hd__clkbuf_1 _4079_ (.A(_2039_),
    .X(_0586_));
 sky130_fd_sc_hd__mux2_1 _4080_ (.A0(_1778_),
    .A1(\tms1x00.RAM[16][1] ),
    .S(_2038_),
    .X(_2040_));
 sky130_fd_sc_hd__clkbuf_1 _4081_ (.A(_2040_),
    .X(_0587_));
 sky130_fd_sc_hd__mux2_1 _4082_ (.A0(_1780_),
    .A1(\tms1x00.RAM[16][2] ),
    .S(_2038_),
    .X(_2041_));
 sky130_fd_sc_hd__clkbuf_1 _4083_ (.A(_2041_),
    .X(_0588_));
 sky130_fd_sc_hd__mux2_1 _4084_ (.A0(_1782_),
    .A1(\tms1x00.RAM[16][3] ),
    .S(_2038_),
    .X(_2042_));
 sky130_fd_sc_hd__clkbuf_1 _4085_ (.A(_2042_),
    .X(_0589_));
 sky130_fd_sc_hd__nor2_2 _4086_ (.A(_1176_),
    .B(_1247_),
    .Y(_2043_));
 sky130_fd_sc_hd__mux2_1 _4087_ (.A0(\tms1x00.RAM[119][0] ),
    .A1(_1265_),
    .S(_2043_),
    .X(_2044_));
 sky130_fd_sc_hd__clkbuf_1 _4088_ (.A(_2044_),
    .X(_0590_));
 sky130_fd_sc_hd__mux2_1 _4089_ (.A0(\tms1x00.RAM[119][1] ),
    .A1(_1269_),
    .S(_2043_),
    .X(_2045_));
 sky130_fd_sc_hd__clkbuf_1 _4090_ (.A(_2045_),
    .X(_0591_));
 sky130_fd_sc_hd__mux2_1 _4091_ (.A0(\tms1x00.RAM[119][2] ),
    .A1(_1272_),
    .S(_2043_),
    .X(_2046_));
 sky130_fd_sc_hd__clkbuf_1 _4092_ (.A(_2046_),
    .X(_0592_));
 sky130_fd_sc_hd__mux2_1 _4093_ (.A0(\tms1x00.RAM[119][3] ),
    .A1(_1275_),
    .S(_2043_),
    .X(_2047_));
 sky130_fd_sc_hd__clkbuf_1 _4094_ (.A(_2047_),
    .X(_0593_));
 sky130_fd_sc_hd__or2_2 _4095_ (.A(_1211_),
    .B(_1232_),
    .X(_2048_));
 sky130_fd_sc_hd__mux2_1 _4096_ (.A0(_1130_),
    .A1(\tms1x00.RAM[12][0] ),
    .S(_2048_),
    .X(_2049_));
 sky130_fd_sc_hd__clkbuf_1 _4097_ (.A(_2049_),
    .X(_0594_));
 sky130_fd_sc_hd__mux2_1 _4098_ (.A0(_1138_),
    .A1(\tms1x00.RAM[12][1] ),
    .S(_2048_),
    .X(_2050_));
 sky130_fd_sc_hd__clkbuf_1 _4099_ (.A(_2050_),
    .X(_0595_));
 sky130_fd_sc_hd__mux2_1 _4100_ (.A0(_1140_),
    .A1(\tms1x00.RAM[12][2] ),
    .S(_2048_),
    .X(_2051_));
 sky130_fd_sc_hd__clkbuf_1 _4101_ (.A(_2051_),
    .X(_0596_));
 sky130_fd_sc_hd__mux2_1 _4102_ (.A0(_1142_),
    .A1(\tms1x00.RAM[12][3] ),
    .S(_2048_),
    .X(_2052_));
 sky130_fd_sc_hd__clkbuf_1 _4103_ (.A(_2052_),
    .X(_0597_));
 sky130_fd_sc_hd__or2_2 _4104_ (.A(_1169_),
    .B(_1232_),
    .X(_2053_));
 sky130_fd_sc_hd__mux2_1 _4105_ (.A0(_1130_),
    .A1(\tms1x00.RAM[15][0] ),
    .S(_2053_),
    .X(_2054_));
 sky130_fd_sc_hd__clkbuf_1 _4106_ (.A(_2054_),
    .X(_0598_));
 sky130_fd_sc_hd__mux2_1 _4107_ (.A0(_1138_),
    .A1(\tms1x00.RAM[15][1] ),
    .S(_2053_),
    .X(_2055_));
 sky130_fd_sc_hd__clkbuf_1 _4108_ (.A(_2055_),
    .X(_0599_));
 sky130_fd_sc_hd__mux2_1 _4109_ (.A0(_1140_),
    .A1(\tms1x00.RAM[15][2] ),
    .S(_2053_),
    .X(_2056_));
 sky130_fd_sc_hd__clkbuf_1 _4110_ (.A(_2056_),
    .X(_0600_));
 sky130_fd_sc_hd__mux2_1 _4111_ (.A0(_1142_),
    .A1(\tms1x00.RAM[15][3] ),
    .S(_2053_),
    .X(_2057_));
 sky130_fd_sc_hd__clkbuf_1 _4112_ (.A(_2057_),
    .X(_0601_));
 sky130_fd_sc_hd__buf_4 _4113_ (.A(_1947_),
    .X(_2058_));
 sky130_fd_sc_hd__mux2_1 _4114_ (.A0(\tms1x00.PC[0] ),
    .A1(\tms1x00.rom_addr[0] ),
    .S(_2058_),
    .X(_2059_));
 sky130_fd_sc_hd__clkbuf_1 _4115_ (.A(_2059_),
    .X(_0602_));
 sky130_fd_sc_hd__mux2_1 _4116_ (.A0(\tms1x00.PC[1] ),
    .A1(_1810_),
    .S(_2058_),
    .X(_2060_));
 sky130_fd_sc_hd__clkbuf_1 _4117_ (.A(_2060_),
    .X(_0603_));
 sky130_fd_sc_hd__mux2_1 _4118_ (.A0(\tms1x00.PC[2] ),
    .A1(net52),
    .S(_2058_),
    .X(_2061_));
 sky130_fd_sc_hd__clkbuf_1 _4119_ (.A(_2061_),
    .X(_0604_));
 sky130_fd_sc_hd__mux2_1 _4120_ (.A0(\tms1x00.PC[3] ),
    .A1(net53),
    .S(_2058_),
    .X(_2062_));
 sky130_fd_sc_hd__clkbuf_1 _4121_ (.A(_2062_),
    .X(_0605_));
 sky130_fd_sc_hd__mux2_1 _4122_ (.A0(\tms1x00.PC[4] ),
    .A1(net54),
    .S(_2058_),
    .X(_2063_));
 sky130_fd_sc_hd__clkbuf_1 _4123_ (.A(_2063_),
    .X(_0606_));
 sky130_fd_sc_hd__mux2_1 _4124_ (.A0(\tms1x00.PC[5] ),
    .A1(net55),
    .S(_2058_),
    .X(_2064_));
 sky130_fd_sc_hd__clkbuf_1 _4125_ (.A(_2064_),
    .X(_0607_));
 sky130_fd_sc_hd__mux2_1 _4126_ (.A0(\tms1x00.PA[0] ),
    .A1(net56),
    .S(_2058_),
    .X(_2065_));
 sky130_fd_sc_hd__clkbuf_1 _4127_ (.A(_2065_),
    .X(_0608_));
 sky130_fd_sc_hd__mux2_1 _4128_ (.A0(\tms1x00.PA[1] ),
    .A1(net57),
    .S(_2058_),
    .X(_2066_));
 sky130_fd_sc_hd__clkbuf_1 _4129_ (.A(_2066_),
    .X(_0609_));
 sky130_fd_sc_hd__mux2_1 _4130_ (.A0(\tms1x00.PA[2] ),
    .A1(net58),
    .S(_2058_),
    .X(_2067_));
 sky130_fd_sc_hd__clkbuf_1 _4131_ (.A(_2067_),
    .X(_0610_));
 sky130_fd_sc_hd__mux2_1 _4132_ (.A0(\tms1x00.PA[3] ),
    .A1(net59),
    .S(_2058_),
    .X(_2068_));
 sky130_fd_sc_hd__clkbuf_1 _4133_ (.A(_2068_),
    .X(_0611_));
 sky130_fd_sc_hd__nor2_2 _4134_ (.A(_1135_),
    .B(_1233_),
    .Y(_2069_));
 sky130_fd_sc_hd__mux2_1 _4135_ (.A0(\tms1x00.RAM[9][0] ),
    .A1(_1265_),
    .S(_2069_),
    .X(_2070_));
 sky130_fd_sc_hd__clkbuf_1 _4136_ (.A(_2070_),
    .X(_0612_));
 sky130_fd_sc_hd__mux2_1 _4137_ (.A0(\tms1x00.RAM[9][1] ),
    .A1(_1269_),
    .S(_2069_),
    .X(_2071_));
 sky130_fd_sc_hd__clkbuf_1 _4138_ (.A(_2071_),
    .X(_0613_));
 sky130_fd_sc_hd__mux2_1 _4139_ (.A0(\tms1x00.RAM[9][2] ),
    .A1(_1272_),
    .S(_2069_),
    .X(_2072_));
 sky130_fd_sc_hd__clkbuf_1 _4140_ (.A(_2072_),
    .X(_0614_));
 sky130_fd_sc_hd__mux2_1 _4141_ (.A0(\tms1x00.RAM[9][3] ),
    .A1(_1275_),
    .S(_2069_),
    .X(_2073_));
 sky130_fd_sc_hd__clkbuf_1 _4142_ (.A(_2073_),
    .X(_0615_));
 sky130_fd_sc_hd__dfxtp_1 _4143_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0014_),
    .Q(net36));
 sky130_fd_sc_hd__dfxtp_1 _4144_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0015_),
    .Q(\tms1x00.RAM[99][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4145_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0016_),
    .Q(\tms1x00.RAM[99][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4146_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0017_),
    .Q(\tms1x00.RAM[99][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4147_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0018_),
    .Q(\tms1x00.RAM[99][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4148_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0019_),
    .Q(\tms1x00.RAM[89][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4149_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0020_),
    .Q(\tms1x00.RAM[89][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4150_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0021_),
    .Q(\tms1x00.RAM[89][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4151_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0022_),
    .Q(\tms1x00.RAM[89][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4152_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0023_),
    .Q(\tms1x00.RAM[59][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4153_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0024_),
    .Q(\tms1x00.RAM[59][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4154_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0025_),
    .Q(\tms1x00.RAM[59][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4155_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0026_),
    .Q(\tms1x00.RAM[59][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4156_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0027_),
    .Q(\tms1x00.RAM[109][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4157_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0028_),
    .Q(\tms1x00.RAM[109][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4158_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0029_),
    .Q(\tms1x00.RAM[109][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4159_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0030_),
    .Q(\tms1x00.RAM[109][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4160_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0031_),
    .Q(\tms1x00.RAM[69][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4161_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0032_),
    .Q(\tms1x00.RAM[69][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4162_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0033_),
    .Q(\tms1x00.RAM[69][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4163_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0034_),
    .Q(\tms1x00.RAM[69][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4164_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0035_),
    .Q(\tms1x00.RAM[79][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4165_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0036_),
    .Q(\tms1x00.RAM[79][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4166_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0037_),
    .Q(\tms1x00.RAM[79][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4167_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0038_),
    .Q(\tms1x00.RAM[79][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4168_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0039_),
    .Q(\tms1x00.RAM[127][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4169_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0040_),
    .Q(\tms1x00.RAM[127][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4170_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0041_),
    .Q(\tms1x00.RAM[127][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4171_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0042_),
    .Q(\tms1x00.RAM[127][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4172_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0043_),
    .Q(\tms1x00.RAM[49][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4173_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0044_),
    .Q(\tms1x00.RAM[49][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4174_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0045_),
    .Q(\tms1x00.RAM[49][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4175_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0046_),
    .Q(\tms1x00.RAM[49][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4176_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0047_),
    .Q(\tms1x00.RAM[19][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4177_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0048_),
    .Q(\tms1x00.RAM[19][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4178_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0049_),
    .Q(\tms1x00.RAM[19][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4179_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0050_),
    .Q(\tms1x00.RAM[19][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4180_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0051_),
    .Q(\tms1x00.RAM[95][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4181_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0052_),
    .Q(\tms1x00.RAM[95][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4182_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0053_),
    .Q(\tms1x00.RAM[95][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4183_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0054_),
    .Q(\tms1x00.RAM[95][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4184_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0055_),
    .Q(\tms1x00.RAM[94][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4185_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0056_),
    .Q(\tms1x00.RAM[94][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4186_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0057_),
    .Q(\tms1x00.RAM[94][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4187_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0058_),
    .Q(\tms1x00.RAM[94][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4188_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0059_),
    .Q(\tms1x00.RAM[93][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4189_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0060_),
    .Q(\tms1x00.RAM[93][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4190_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0061_),
    .Q(\tms1x00.RAM[93][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4191_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0062_),
    .Q(\tms1x00.RAM[93][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4192_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0063_),
    .Q(\tms1x00.RAM[92][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4193_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0064_),
    .Q(\tms1x00.RAM[92][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4194_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0065_),
    .Q(\tms1x00.RAM[92][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4195_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0066_),
    .Q(\tms1x00.RAM[92][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4196_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0067_),
    .Q(\tms1x00.RAM[91][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4197_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0068_),
    .Q(\tms1x00.RAM[91][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4198_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0069_),
    .Q(\tms1x00.RAM[91][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4199_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0070_),
    .Q(\tms1x00.RAM[91][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4200_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0071_),
    .Q(\tms1x00.RAM[90][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4201_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0072_),
    .Q(\tms1x00.RAM[90][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4202_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0073_),
    .Q(\tms1x00.RAM[90][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4203_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0074_),
    .Q(\tms1x00.RAM[90][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4204_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0075_),
    .Q(\tms1x00.RAM[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4205_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0076_),
    .Q(\tms1x00.RAM[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4206_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0077_),
    .Q(\tms1x00.RAM[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4207_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0078_),
    .Q(\tms1x00.RAM[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4208_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0079_),
    .Q(\tms1x00.RAM[88][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4209_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0080_),
    .Q(\tms1x00.RAM[88][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4210_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0081_),
    .Q(\tms1x00.RAM[88][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4211_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0082_),
    .Q(\tms1x00.RAM[88][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4212_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0083_),
    .Q(\tms1x00.RAM[87][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4213_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0084_),
    .Q(\tms1x00.RAM[87][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4214_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0085_),
    .Q(\tms1x00.RAM[87][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4215_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0086_),
    .Q(\tms1x00.RAM[87][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4216_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0087_),
    .Q(\tms1x00.RAM[86][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4217_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0088_),
    .Q(\tms1x00.RAM[86][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4218_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0089_),
    .Q(\tms1x00.RAM[86][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4219_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0090_),
    .Q(\tms1x00.RAM[86][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4220_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0091_),
    .Q(\tms1x00.RAM[105][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4221_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0092_),
    .Q(\tms1x00.RAM[105][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4222_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0093_),
    .Q(\tms1x00.RAM[105][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4223_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0094_),
    .Q(\tms1x00.RAM[105][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4224_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0095_),
    .Q(\tms1x00.RAM[104][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4225_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0096_),
    .Q(\tms1x00.RAM[104][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4226_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0097_),
    .Q(\tms1x00.RAM[104][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4227_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0098_),
    .Q(\tms1x00.RAM[104][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4228_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0099_),
    .Q(\tms1x00.RAM[103][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4229_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0100_),
    .Q(\tms1x00.RAM[103][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4230_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0101_),
    .Q(\tms1x00.RAM[103][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4231_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0102_),
    .Q(\tms1x00.RAM[103][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4232_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0103_),
    .Q(\tms1x00.RAM[102][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4233_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0104_),
    .Q(\tms1x00.RAM[102][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4234_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0105_),
    .Q(\tms1x00.RAM[102][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4235_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0106_),
    .Q(\tms1x00.RAM[102][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4236_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0107_),
    .Q(\tms1x00.RAM[101][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4237_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0108_),
    .Q(\tms1x00.RAM[101][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4238_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0109_),
    .Q(\tms1x00.RAM[101][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4239_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0110_),
    .Q(\tms1x00.RAM[101][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4240_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0111_),
    .Q(\tms1x00.RAM[100][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4241_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0112_),
    .Q(\tms1x00.RAM[100][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4242_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0113_),
    .Q(\tms1x00.RAM[100][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4243_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0114_),
    .Q(\tms1x00.RAM[100][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4244_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0115_),
    .Q(\tms1x00.RAM[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4245_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0116_),
    .Q(\tms1x00.RAM[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4246_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0117_),
    .Q(\tms1x00.RAM[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4247_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0118_),
    .Q(\tms1x00.RAM[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4248_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0119_),
    .Q(\tms1x00.RAM[98][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4249_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0120_),
    .Q(\tms1x00.RAM[98][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4250_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0121_),
    .Q(\tms1x00.RAM[98][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4251_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0122_),
    .Q(\tms1x00.RAM[98][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4252_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0123_),
    .Q(\tms1x00.RAM[97][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4253_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0124_),
    .Q(\tms1x00.RAM[97][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4254_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0125_),
    .Q(\tms1x00.RAM[97][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4255_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0126_),
    .Q(\tms1x00.RAM[97][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4256_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0127_),
    .Q(\tms1x00.RAM[96][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4257_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0128_),
    .Q(\tms1x00.RAM[96][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4258_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0129_),
    .Q(\tms1x00.RAM[96][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4259_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0130_),
    .Q(\tms1x00.RAM[96][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4260_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0131_),
    .Q(\tms1x00.RAM[115][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4261_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0132_),
    .Q(\tms1x00.RAM[115][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4262_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0133_),
    .Q(\tms1x00.RAM[115][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4263_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0134_),
    .Q(\tms1x00.RAM[115][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4264_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0135_),
    .Q(\tms1x00.RAM[114][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4265_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0136_),
    .Q(\tms1x00.RAM[114][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4266_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0137_),
    .Q(\tms1x00.RAM[114][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4267_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0138_),
    .Q(\tms1x00.RAM[114][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4268_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0139_),
    .Q(\tms1x00.RAM[113][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4269_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0140_),
    .Q(\tms1x00.RAM[113][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4270_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0141_),
    .Q(\tms1x00.RAM[113][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4271_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0142_),
    .Q(\tms1x00.RAM[113][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4272_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0143_),
    .Q(\tms1x00.RAM[112][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4273_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0144_),
    .Q(\tms1x00.RAM[112][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4274_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0145_),
    .Q(\tms1x00.RAM[112][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4275_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0146_),
    .Q(\tms1x00.RAM[112][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4276_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0147_),
    .Q(\tms1x00.RAM[111][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4277_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0148_),
    .Q(\tms1x00.RAM[111][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4278_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0149_),
    .Q(\tms1x00.RAM[111][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4279_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0150_),
    .Q(\tms1x00.RAM[111][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4280_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0151_),
    .Q(\tms1x00.RAM[110][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4281_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0152_),
    .Q(\tms1x00.RAM[110][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4282_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0153_),
    .Q(\tms1x00.RAM[110][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4283_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0154_),
    .Q(\tms1x00.RAM[110][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4284_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0155_),
    .Q(\tms1x00.RAM[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4285_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0156_),
    .Q(\tms1x00.RAM[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4286_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0157_),
    .Q(\tms1x00.RAM[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4287_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0158_),
    .Q(\tms1x00.RAM[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4288_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0159_),
    .Q(\tms1x00.RAM[108][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4289_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0160_),
    .Q(\tms1x00.RAM[108][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4290_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0161_),
    .Q(\tms1x00.RAM[108][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4291_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0162_),
    .Q(\tms1x00.RAM[108][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4292_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0163_),
    .Q(\tms1x00.RAM[107][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4293_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0164_),
    .Q(\tms1x00.RAM[107][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4294_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0165_),
    .Q(\tms1x00.RAM[107][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4295_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0166_),
    .Q(\tms1x00.RAM[107][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4296_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0167_),
    .Q(\tms1x00.RAM[106][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4297_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0168_),
    .Q(\tms1x00.RAM[106][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4298_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0169_),
    .Q(\tms1x00.RAM[106][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4299_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0170_),
    .Q(\tms1x00.RAM[106][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4300_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0171_),
    .Q(\tms1x00.RAM[125][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4301_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0172_),
    .Q(\tms1x00.RAM[125][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4302_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0173_),
    .Q(\tms1x00.RAM[125][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4303_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0174_),
    .Q(\tms1x00.RAM[125][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4304_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0175_),
    .Q(\tms1x00.RAM[124][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4305_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0176_),
    .Q(\tms1x00.RAM[124][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4306_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0177_),
    .Q(\tms1x00.RAM[124][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4307_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0178_),
    .Q(\tms1x00.RAM[124][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4308_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0179_),
    .Q(\tms1x00.RAM[123][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4309_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0180_),
    .Q(\tms1x00.RAM[123][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4310_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0181_),
    .Q(\tms1x00.RAM[123][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4311_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0182_),
    .Q(\tms1x00.RAM[123][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4312_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0183_),
    .Q(\tms1x00.RAM[122][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4313_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0184_),
    .Q(\tms1x00.RAM[122][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4314_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0185_),
    .Q(\tms1x00.RAM[122][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4315_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0186_),
    .Q(\tms1x00.RAM[122][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4316_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0187_),
    .Q(\tms1x00.RAM[121][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4317_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0188_),
    .Q(\tms1x00.RAM[121][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4318_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0189_),
    .Q(\tms1x00.RAM[121][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4319_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0190_),
    .Q(\tms1x00.RAM[121][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4320_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0191_),
    .Q(\tms1x00.RAM[120][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4321_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0192_),
    .Q(\tms1x00.RAM[120][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4322_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0193_),
    .Q(\tms1x00.RAM[120][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4323_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0194_),
    .Q(\tms1x00.RAM[120][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4324_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0195_),
    .Q(\tms1x00.RAM[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4325_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0196_),
    .Q(\tms1x00.RAM[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4326_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0197_),
    .Q(\tms1x00.RAM[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4327_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0198_),
    .Q(\tms1x00.RAM[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4328_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0199_),
    .Q(\tms1x00.RAM[118][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4329_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0200_),
    .Q(\tms1x00.RAM[118][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4330_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0201_),
    .Q(\tms1x00.RAM[118][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4331_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0202_),
    .Q(\tms1x00.RAM[118][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4332_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0203_),
    .Q(\tms1x00.RAM[117][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4333_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0204_),
    .Q(\tms1x00.RAM[117][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4334_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0205_),
    .Q(\tms1x00.RAM[117][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4335_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0206_),
    .Q(\tms1x00.RAM[117][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4336_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0207_),
    .Q(\tms1x00.RAM[116][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4337_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0208_),
    .Q(\tms1x00.RAM[116][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4338_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0209_),
    .Q(\tms1x00.RAM[116][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4339_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0210_),
    .Q(\tms1x00.RAM[116][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4340_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0211_),
    .Q(\tms1x00.RAM[126][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4341_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0212_),
    .Q(\tms1x00.RAM[126][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4342_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0213_),
    .Q(\tms1x00.RAM[126][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4343_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0214_),
    .Q(\tms1x00.RAM[126][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4344_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0215_),
    .Q(\tms1x00.RAM[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4345_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0216_),
    .Q(\tms1x00.RAM[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4346_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0217_),
    .Q(\tms1x00.RAM[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4347_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0218_),
    .Q(\tms1x00.RAM[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4348_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0219_),
    .Q(\tms1x00.RAM[23][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4349_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0220_),
    .Q(\tms1x00.RAM[23][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4350_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0221_),
    .Q(\tms1x00.RAM[23][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4351_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0222_),
    .Q(\tms1x00.RAM[23][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4352_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0223_),
    .Q(\tms1x00.RAM[22][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4353_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0224_),
    .Q(\tms1x00.RAM[22][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4354_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0225_),
    .Q(\tms1x00.RAM[22][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4355_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0226_),
    .Q(\tms1x00.RAM[22][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4356_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0227_),
    .Q(\tms1x00.RAM[21][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4357_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0228_),
    .Q(\tms1x00.RAM[21][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4358_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0229_),
    .Q(\tms1x00.RAM[21][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4359_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0230_),
    .Q(\tms1x00.RAM[21][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4360_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0231_),
    .Q(\tms1x00.RAM[20][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4361_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0232_),
    .Q(\tms1x00.RAM[20][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4362_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0233_),
    .Q(\tms1x00.RAM[20][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4363_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0234_),
    .Q(\tms1x00.RAM[20][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4364_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0235_),
    .Q(\tms1x00.RAM[28][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4365_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0236_),
    .Q(\tms1x00.RAM[28][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4366_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0237_),
    .Q(\tms1x00.RAM[28][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4367_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0238_),
    .Q(\tms1x00.RAM[28][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4368_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0239_),
    .Q(\tms1x00.RAM[27][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4369_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0240_),
    .Q(\tms1x00.RAM[27][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4370_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0241_),
    .Q(\tms1x00.RAM[27][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4371_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0242_),
    .Q(\tms1x00.RAM[27][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4372_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0243_),
    .Q(\tms1x00.RAM[26][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4373_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0244_),
    .Q(\tms1x00.RAM[26][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4374_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0245_),
    .Q(\tms1x00.RAM[26][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4375_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0246_),
    .Q(\tms1x00.RAM[26][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4376_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0247_),
    .Q(\tms1x00.RAM[25][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4377_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0248_),
    .Q(\tms1x00.RAM[25][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4378_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0249_),
    .Q(\tms1x00.RAM[25][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4379_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0250_),
    .Q(\tms1x00.RAM[25][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4380_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0251_),
    .Q(\tms1x00.RAM[24][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4381_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0252_),
    .Q(\tms1x00.RAM[24][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4382_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0253_),
    .Q(\tms1x00.RAM[24][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4383_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0254_),
    .Q(\tms1x00.RAM[24][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4384_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0255_),
    .Q(\tms1x00.RAM[32][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4385_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0256_),
    .Q(\tms1x00.RAM[32][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4386_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0257_),
    .Q(\tms1x00.RAM[32][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4387_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0258_),
    .Q(\tms1x00.RAM[32][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4388_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0259_),
    .Q(\tms1x00.RAM[31][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4389_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0260_),
    .Q(\tms1x00.RAM[31][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4390_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0261_),
    .Q(\tms1x00.RAM[31][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4391_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0262_),
    .Q(\tms1x00.RAM[31][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4392_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0263_),
    .Q(\tms1x00.RAM[30][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4393_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0264_),
    .Q(\tms1x00.RAM[30][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4394_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0265_),
    .Q(\tms1x00.RAM[30][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4395_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0266_),
    .Q(\tms1x00.RAM[30][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4396_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0267_),
    .Q(\tms1x00.RAM[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4397_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0268_),
    .Q(\tms1x00.RAM[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4398_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0269_),
    .Q(\tms1x00.RAM[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4399_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0270_),
    .Q(\tms1x00.RAM[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4400_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0271_),
    .Q(\tms1x00.RAM[36][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4401_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0272_),
    .Q(\tms1x00.RAM[36][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4402_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0273_),
    .Q(\tms1x00.RAM[36][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4403_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0274_),
    .Q(\tms1x00.RAM[36][3] ));
 sky130_fd_sc_hd__dfxtp_2 _4404_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0007_),
    .Q(_0000_));
 sky130_fd_sc_hd__dfxtp_2 _4405_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0008_),
    .Q(_0001_));
 sky130_fd_sc_hd__dfxtp_1 _4406_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0009_),
    .Q(_0002_));
 sky130_fd_sc_hd__dfxtp_2 _4407_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0010_),
    .Q(_0003_));
 sky130_fd_sc_hd__dfxtp_4 _4408_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0011_),
    .Q(_0004_));
 sky130_fd_sc_hd__dfxtp_1 _4409_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0012_),
    .Q(_0005_));
 sky130_fd_sc_hd__dfxtp_2 _4410_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0013_),
    .Q(_0006_));
 sky130_fd_sc_hd__dfxtp_1 _4411_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0275_),
    .Q(\tms1x00.RAM[35][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4412_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0276_),
    .Q(\tms1x00.RAM[35][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4413_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0277_),
    .Q(\tms1x00.RAM[35][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4414_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0278_),
    .Q(\tms1x00.RAM[35][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4415_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0279_),
    .Q(\tms1x00.RAM[34][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4416_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0280_),
    .Q(\tms1x00.RAM[34][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4417_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0281_),
    .Q(\tms1x00.RAM[34][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4418_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0282_),
    .Q(\tms1x00.RAM[34][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4419_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0283_),
    .Q(\tms1x00.RAM[33][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4420_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0284_),
    .Q(\tms1x00.RAM[33][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4421_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0285_),
    .Q(\tms1x00.RAM[33][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4422_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0286_),
    .Q(\tms1x00.RAM[33][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4423_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0287_),
    .Q(\tms1x00.RAM[41][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4424_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0288_),
    .Q(\tms1x00.RAM[41][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4425_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0289_),
    .Q(\tms1x00.RAM[41][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4426_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0290_),
    .Q(\tms1x00.RAM[41][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4427_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0291_),
    .Q(\tms1x00.RAM[40][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4428_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0292_),
    .Q(\tms1x00.RAM[40][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4429_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0293_),
    .Q(\tms1x00.RAM[40][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4430_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0294_),
    .Q(\tms1x00.RAM[40][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4431_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0295_),
    .Q(\tms1x00.RAM[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4432_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0296_),
    .Q(\tms1x00.RAM[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4433_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0297_),
    .Q(\tms1x00.RAM[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4434_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0298_),
    .Q(\tms1x00.RAM[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4435_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0299_),
    .Q(\tms1x00.RAM[38][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4436_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0300_),
    .Q(\tms1x00.RAM[38][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4437_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0301_),
    .Q(\tms1x00.RAM[38][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4438_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0302_),
    .Q(\tms1x00.RAM[38][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4439_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0303_),
    .Q(\tms1x00.RAM[37][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4440_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0304_),
    .Q(\tms1x00.RAM[37][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4441_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0305_),
    .Q(\tms1x00.RAM[37][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4442_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0306_),
    .Q(\tms1x00.RAM[37][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4443_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0307_),
    .Q(\tms1x00.RAM[45][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4444_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0308_),
    .Q(\tms1x00.RAM[45][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4445_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0309_),
    .Q(\tms1x00.RAM[45][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4446_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0310_),
    .Q(\tms1x00.RAM[45][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4447_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0311_),
    .Q(\tms1x00.RAM[44][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4448_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0312_),
    .Q(\tms1x00.RAM[44][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4449_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0313_),
    .Q(\tms1x00.RAM[44][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4450_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0314_),
    .Q(\tms1x00.RAM[44][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4451_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0315_),
    .Q(\tms1x00.RAM[43][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4452_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0316_),
    .Q(\tms1x00.RAM[43][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4453_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0317_),
    .Q(\tms1x00.RAM[43][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4454_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0318_),
    .Q(\tms1x00.RAM[43][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4455_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0319_),
    .Q(\tms1x00.RAM[42][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4456_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0320_),
    .Q(\tms1x00.RAM[42][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4457_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0321_),
    .Q(\tms1x00.RAM[42][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4458_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0322_),
    .Q(\tms1x00.RAM[42][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4459_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0323_),
    .Q(\tms1x00.RAM[50][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4460_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0324_),
    .Q(\tms1x00.RAM[50][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4461_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0325_),
    .Q(\tms1x00.RAM[50][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4462_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0326_),
    .Q(\tms1x00.RAM[50][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4463_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0327_),
    .Q(\tms1x00.RAM[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4464_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0328_),
    .Q(\tms1x00.RAM[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4465_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0329_),
    .Q(\tms1x00.RAM[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4466_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0330_),
    .Q(\tms1x00.RAM[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4467_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0331_),
    .Q(\tms1x00.RAM[48][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4468_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0332_),
    .Q(\tms1x00.RAM[48][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4469_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0333_),
    .Q(\tms1x00.RAM[48][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4470_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0334_),
    .Q(\tms1x00.RAM[48][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4471_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0335_),
    .Q(\tms1x00.RAM[47][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4472_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0336_),
    .Q(\tms1x00.RAM[47][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4473_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0337_),
    .Q(\tms1x00.RAM[47][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4474_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0338_),
    .Q(\tms1x00.RAM[47][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4475_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0339_),
    .Q(\tms1x00.RAM[46][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4476_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0340_),
    .Q(\tms1x00.RAM[46][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4477_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0341_),
    .Q(\tms1x00.RAM[46][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4478_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0342_),
    .Q(\tms1x00.RAM[46][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4479_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0343_),
    .Q(\tms1x00.RAM[54][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4480_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0344_),
    .Q(\tms1x00.RAM[54][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4481_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0345_),
    .Q(\tms1x00.RAM[54][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4482_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0346_),
    .Q(\tms1x00.RAM[54][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4483_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0347_),
    .Q(\tms1x00.RAM[53][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4484_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0348_),
    .Q(\tms1x00.RAM[53][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4485_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0349_),
    .Q(\tms1x00.RAM[53][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4486_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0350_),
    .Q(\tms1x00.RAM[53][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4487_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0351_),
    .Q(\tms1x00.RAM[52][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4488_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0352_),
    .Q(\tms1x00.RAM[52][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4489_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0353_),
    .Q(\tms1x00.RAM[52][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4490_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0354_),
    .Q(\tms1x00.RAM[52][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4491_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0355_),
    .Q(\tms1x00.RAM[51][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4492_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0356_),
    .Q(\tms1x00.RAM[51][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4493_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0357_),
    .Q(\tms1x00.RAM[51][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4494_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0358_),
    .Q(\tms1x00.RAM[51][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4495_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0359_),
    .Q(\tms1x00.RAM[58][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4496_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0360_),
    .Q(\tms1x00.RAM[58][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4497_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0361_),
    .Q(\tms1x00.RAM[58][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4498_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0362_),
    .Q(\tms1x00.RAM[58][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4499_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0363_),
    .Q(\tms1x00.RAM[57][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4500_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0364_),
    .Q(\tms1x00.RAM[57][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4501_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0365_),
    .Q(\tms1x00.RAM[57][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4502_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0366_),
    .Q(\tms1x00.RAM[57][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4503_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0367_),
    .Q(\tms1x00.RAM[56][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4504_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0368_),
    .Q(\tms1x00.RAM[56][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4505_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0369_),
    .Q(\tms1x00.RAM[56][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4506_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0370_),
    .Q(\tms1x00.RAM[56][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4507_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0371_),
    .Q(\tms1x00.RAM[55][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4508_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0372_),
    .Q(\tms1x00.RAM[55][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4509_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0373_),
    .Q(\tms1x00.RAM[55][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4510_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0374_),
    .Q(\tms1x00.RAM[55][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4511_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0375_),
    .Q(\tms1x00.RAM[63][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4512_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0376_),
    .Q(\tms1x00.RAM[63][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4513_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0377_),
    .Q(\tms1x00.RAM[63][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4514_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0378_),
    .Q(\tms1x00.RAM[63][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4515_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0379_),
    .Q(\tms1x00.RAM[62][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4516_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0380_),
    .Q(\tms1x00.RAM[62][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4517_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0381_),
    .Q(\tms1x00.RAM[62][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4518_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0382_),
    .Q(\tms1x00.RAM[62][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4519_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0383_),
    .Q(\tms1x00.RAM[61][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4520_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0384_),
    .Q(\tms1x00.RAM[61][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4521_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0385_),
    .Q(\tms1x00.RAM[61][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4522_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0386_),
    .Q(\tms1x00.RAM[61][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4523_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0387_),
    .Q(\tms1x00.RAM[60][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4524_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0388_),
    .Q(\tms1x00.RAM[60][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4525_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0389_),
    .Q(\tms1x00.RAM[60][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4526_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0390_),
    .Q(\tms1x00.RAM[60][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4527_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0391_),
    .Q(\tms1x00.RAM[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4528_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0392_),
    .Q(\tms1x00.RAM[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4529_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0393_),
    .Q(\tms1x00.RAM[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4530_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0394_),
    .Q(\tms1x00.RAM[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4531_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0395_),
    .Q(\tms1x00.RAM[67][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4532_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0396_),
    .Q(\tms1x00.RAM[67][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4533_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0397_),
    .Q(\tms1x00.RAM[67][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4534_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0398_),
    .Q(\tms1x00.RAM[67][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4535_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0399_),
    .Q(\tms1x00.RAM[66][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4536_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0400_),
    .Q(\tms1x00.RAM[66][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4537_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0401_),
    .Q(\tms1x00.RAM[66][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4538_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0402_),
    .Q(\tms1x00.RAM[66][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4539_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0403_),
    .Q(\tms1x00.RAM[65][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4540_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0404_),
    .Q(\tms1x00.RAM[65][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4541_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0405_),
    .Q(\tms1x00.RAM[65][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4542_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0406_),
    .Q(\tms1x00.RAM[65][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4543_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0407_),
    .Q(\tms1x00.RAM[64][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4544_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0408_),
    .Q(\tms1x00.RAM[64][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4545_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0409_),
    .Q(\tms1x00.RAM[64][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4546_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0410_),
    .Q(\tms1x00.RAM[64][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4547_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0411_),
    .Q(\tms1x00.RAM[71][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4548_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0412_),
    .Q(\tms1x00.RAM[71][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4549_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0413_),
    .Q(\tms1x00.RAM[71][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4550_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0414_),
    .Q(\tms1x00.RAM[71][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4551_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0415_),
    .Q(\tms1x00.RAM[70][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4552_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0416_),
    .Q(\tms1x00.RAM[70][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4553_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0417_),
    .Q(\tms1x00.RAM[70][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4554_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0418_),
    .Q(\tms1x00.RAM[70][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4555_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0419_),
    .Q(\tms1x00.RAM[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4556_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0420_),
    .Q(\tms1x00.RAM[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4557_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0421_),
    .Q(\tms1x00.RAM[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4558_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0422_),
    .Q(\tms1x00.RAM[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4559_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0423_),
    .Q(\tms1x00.RAM[68][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4560_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0424_),
    .Q(\tms1x00.RAM[68][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4561_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0425_),
    .Q(\tms1x00.RAM[68][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4562_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0426_),
    .Q(\tms1x00.RAM[68][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4563_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0427_),
    .Q(\tms1x00.RAM[76][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4564_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0428_),
    .Q(\tms1x00.RAM[76][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4565_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0429_),
    .Q(\tms1x00.RAM[76][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4566_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0430_),
    .Q(\tms1x00.RAM[76][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4567_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0431_),
    .Q(\tms1x00.RAM[75][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4568_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0432_),
    .Q(\tms1x00.RAM[75][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4569_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0433_),
    .Q(\tms1x00.RAM[75][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4570_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0434_),
    .Q(\tms1x00.RAM[75][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4571_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0435_),
    .Q(\tms1x00.RAM[74][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4572_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0436_),
    .Q(\tms1x00.RAM[74][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4573_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0437_),
    .Q(\tms1x00.RAM[74][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4574_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0438_),
    .Q(\tms1x00.RAM[74][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4575_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0439_),
    .Q(\tms1x00.RAM[73][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4576_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0440_),
    .Q(\tms1x00.RAM[73][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4577_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0441_),
    .Q(\tms1x00.RAM[73][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4578_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0442_),
    .Q(\tms1x00.RAM[73][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4579_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0443_),
    .Q(\tms1x00.RAM[72][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4580_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0444_),
    .Q(\tms1x00.RAM[72][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4581_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0445_),
    .Q(\tms1x00.RAM[72][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4582_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0446_),
    .Q(\tms1x00.RAM[72][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4583_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0447_),
    .Q(\tms1x00.RAM[77][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4584_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0448_),
    .Q(\tms1x00.RAM[77][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4585_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0449_),
    .Q(\tms1x00.RAM[77][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4586_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0450_),
    .Q(\tms1x00.RAM[77][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4587_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0451_),
    .Q(\tms1x00.RAM[80][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4588_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0452_),
    .Q(\tms1x00.RAM[80][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4589_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0453_),
    .Q(\tms1x00.RAM[80][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4590_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0454_),
    .Q(\tms1x00.RAM[80][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4591_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0455_),
    .Q(\tms1x00.RAM[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4592_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0456_),
    .Q(\tms1x00.RAM[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4593_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0457_),
    .Q(\tms1x00.RAM[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4594_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0458_),
    .Q(\tms1x00.RAM[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4595_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0459_),
    .Q(\tms1x00.RAM[78][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4596_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0460_),
    .Q(\tms1x00.RAM[78][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4597_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0461_),
    .Q(\tms1x00.RAM[78][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4598_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0462_),
    .Q(\tms1x00.RAM[78][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4599_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0463_),
    .Q(\tms1x00.RAM[85][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4600_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0464_),
    .Q(\tms1x00.RAM[85][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4601_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0465_),
    .Q(\tms1x00.RAM[85][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4602_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0466_),
    .Q(\tms1x00.RAM[85][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4603_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0467_),
    .Q(\tms1x00.RAM[84][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4604_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0468_),
    .Q(\tms1x00.RAM[84][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4605_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0469_),
    .Q(\tms1x00.RAM[84][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4606_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0470_),
    .Q(\tms1x00.RAM[84][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4607_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0471_),
    .Q(\tms1x00.RAM[83][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4608_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0472_),
    .Q(\tms1x00.RAM[83][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4609_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0473_),
    .Q(\tms1x00.RAM[83][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4610_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0474_),
    .Q(\tms1x00.RAM[83][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4611_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0475_),
    .Q(\tms1x00.RAM[82][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4612_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0476_),
    .Q(\tms1x00.RAM[82][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4613_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0477_),
    .Q(\tms1x00.RAM[82][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4614_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0478_),
    .Q(\tms1x00.RAM[82][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4615_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0479_),
    .Q(\tms1x00.RAM[81][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4616_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0480_),
    .Q(\tms1x00.RAM[81][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4617_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0481_),
    .Q(\tms1x00.RAM[81][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4618_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0482_),
    .Q(\tms1x00.RAM[81][3] ));
 sky130_fd_sc_hd__dfxtp_2 _4619_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0483_),
    .Q(\tms1x00.ram_addr_buff[0] ));
 sky130_fd_sc_hd__dfxtp_2 _4620_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0484_),
    .Q(\tms1x00.ram_addr_buff[1] ));
 sky130_fd_sc_hd__dfxtp_2 _4621_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0485_),
    .Q(\tms1x00.ram_addr_buff[2] ));
 sky130_fd_sc_hd__dfxtp_2 _4622_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0486_),
    .Q(\tms1x00.ram_addr_buff[3] ));
 sky130_fd_sc_hd__dfxtp_4 _4623_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0487_),
    .Q(\tms1x00.ram_addr_buff[4] ));
 sky130_fd_sc_hd__dfxtp_4 _4624_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0488_),
    .Q(\tms1x00.ram_addr_buff[5] ));
 sky130_fd_sc_hd__dfxtp_4 _4625_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0489_),
    .Q(\tms1x00.ram_addr_buff[6] ));
 sky130_fd_sc_hd__dfxtp_4 _4626_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0490_),
    .Q(net33));
 sky130_fd_sc_hd__dfxtp_4 _4627_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0491_),
    .Q(net34));
 sky130_fd_sc_hd__dfxtp_2 _4628_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0492_),
    .Q(net35));
 sky130_fd_sc_hd__dfxtp_2 _4629_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0493_),
    .Q(\tms1x00.ins_in[0] ));
 sky130_fd_sc_hd__dfxtp_2 _4630_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0494_),
    .Q(\tms1x00.ins_in[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4631_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0495_),
    .Q(\tms1x00.ins_in[2] ));
 sky130_fd_sc_hd__dfxtp_2 _4632_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0496_),
    .Q(\tms1x00.ins_in[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4633_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0497_),
    .Q(\tms1x00.ins_in[4] ));
 sky130_fd_sc_hd__dfxtp_1 _4634_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0498_),
    .Q(\tms1x00.ins_in[5] ));
 sky130_fd_sc_hd__dfxtp_1 _4635_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0499_),
    .Q(\tms1x00.ins_in[6] ));
 sky130_fd_sc_hd__dfxtp_2 _4636_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0500_),
    .Q(\tms1x00.ins_in[7] ));
 sky130_fd_sc_hd__dfxtp_1 _4637_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net1),
    .Q(\tms1x00.K_latch[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4638_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net2),
    .Q(\tms1x00.K_latch[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4639_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net3),
    .Q(\tms1x00.K_latch[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4640_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net4),
    .Q(\tms1x00.K_latch[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4641_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0501_),
    .Q(net37));
 sky130_fd_sc_hd__dfxtp_1 _4642_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0502_),
    .Q(net38));
 sky130_fd_sc_hd__dfxtp_1 _4643_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0503_),
    .Q(net39));
 sky130_fd_sc_hd__dfxtp_1 _4644_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0504_),
    .Q(net40));
 sky130_fd_sc_hd__dfxtp_1 _4645_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0505_),
    .Q(net41));
 sky130_fd_sc_hd__dfxtp_1 _4646_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0506_),
    .Q(net42));
 sky130_fd_sc_hd__dfxtp_1 _4647_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0507_),
    .Q(net43));
 sky130_fd_sc_hd__dfxtp_1 _4648_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0508_),
    .Q(net44));
 sky130_fd_sc_hd__dfxtp_1 _4649_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0509_),
    .Q(net45));
 sky130_fd_sc_hd__dfxtp_1 _4650_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0510_),
    .Q(net46));
 sky130_fd_sc_hd__dfxtp_1 _4651_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0511_),
    .Q(net47));
 sky130_fd_sc_hd__dfxtp_1 _4652_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0512_),
    .Q(net48));
 sky130_fd_sc_hd__dfxtp_1 _4653_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0513_),
    .Q(net49));
 sky130_fd_sc_hd__dfxtp_1 _4654_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0514_),
    .Q(net50));
 sky130_fd_sc_hd__dfxtp_1 _4655_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0515_),
    .Q(net51));
 sky130_fd_sc_hd__dfxtp_1 _4656_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0516_),
    .Q(net28));
 sky130_fd_sc_hd__dfxtp_1 _4657_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0517_),
    .Q(net29));
 sky130_fd_sc_hd__dfxtp_1 _4658_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0518_),
    .Q(net30));
 sky130_fd_sc_hd__dfxtp_1 _4659_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0519_),
    .Q(net31));
 sky130_fd_sc_hd__dfxtp_1 _4660_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0520_),
    .Q(net32));
 sky130_fd_sc_hd__dfxtp_1 _4661_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0521_),
    .Q(\tms1x00.CL ));
 sky130_fd_sc_hd__dfxtp_1 _4662_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0522_),
    .Q(\tms1x00.status ));
 sky130_fd_sc_hd__dfxtp_1 _4663_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0523_),
    .Q(\tms1x00.PB[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4664_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0524_),
    .Q(\tms1x00.PB[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4665_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0525_),
    .Q(\tms1x00.PB[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4666_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0526_),
    .Q(\tms1x00.PB[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4667_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0527_),
    .Q(\tms1x00.SR[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4668_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0528_),
    .Q(\tms1x00.SR[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4669_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0529_),
    .Q(\tms1x00.SR[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4670_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0530_),
    .Q(\tms1x00.SR[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4671_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0531_),
    .Q(\tms1x00.SR[4] ));
 sky130_fd_sc_hd__dfxtp_1 _4672_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0532_),
    .Q(\tms1x00.SR[5] ));
 sky130_fd_sc_hd__dfxtp_1 _4673_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0533_),
    .Q(\tms1x00.PA[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4674_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0534_),
    .Q(\tms1x00.PA[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4675_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0535_),
    .Q(\tms1x00.PA[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4676_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0536_),
    .Q(\tms1x00.PA[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4677_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0537_),
    .Q(\tms1x00.PC[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4678_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0538_),
    .Q(\tms1x00.PC[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4679_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0539_),
    .Q(\tms1x00.PC[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4680_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0540_),
    .Q(\tms1x00.PC[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4681_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0541_),
    .Q(\tms1x00.PC[4] ));
 sky130_fd_sc_hd__dfxtp_1 _4682_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0542_),
    .Q(\tms1x00.PC[5] ));
 sky130_fd_sc_hd__dfxtp_1 _4683_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0543_),
    .Q(\tms1x00.P[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4684_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0544_),
    .Q(\tms1x00.P[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4685_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0545_),
    .Q(\tms1x00.P[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4686_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0546_),
    .Q(\tms1x00.P[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4687_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0547_),
    .Q(\tms1x00.Y[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4688_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0548_),
    .Q(\tms1x00.Y[1] ));
 sky130_fd_sc_hd__dfxtp_2 _4689_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0549_),
    .Q(\tms1x00.Y[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4690_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0550_),
    .Q(\tms1x00.Y[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4691_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0551_),
    .Q(\tms1x00.X[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4692_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0552_),
    .Q(\tms1x00.X[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4693_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0553_),
    .Q(\tms1x00.X[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4694_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0554_),
    .Q(\tms1x00.N[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4695_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0555_),
    .Q(\tms1x00.N[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4696_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0556_),
    .Q(\tms1x00.N[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4697_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0557_),
    .Q(\tms1x00.N[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4698_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0558_),
    .Q(\tms1x00.A[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4699_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0559_),
    .Q(\tms1x00.A[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4700_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0560_),
    .Q(\tms1x00.A[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4701_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0561_),
    .Q(\tms1x00.A[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4702_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0562_),
    .Q(\tms1x00.RAM[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4703_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0563_),
    .Q(\tms1x00.RAM[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4704_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_0564_),
    .Q(\tms1x00.RAM[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4705_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0565_),
    .Q(\tms1x00.RAM[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4706_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0566_),
    .Q(\tms1x00.RAM[18][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4707_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0567_),
    .Q(\tms1x00.RAM[18][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4708_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0568_),
    .Q(\tms1x00.RAM[18][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4709_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0569_),
    .Q(\tms1x00.RAM[18][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4710_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0570_),
    .Q(\tms1x00.RAM[39][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4711_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0571_),
    .Q(\tms1x00.RAM[39][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4712_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0572_),
    .Q(\tms1x00.RAM[39][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4713_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0573_),
    .Q(\tms1x00.RAM[39][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4714_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0574_),
    .Q(\tms1x00.RAM[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4715_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0575_),
    .Q(\tms1x00.RAM[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4716_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0576_),
    .Q(\tms1x00.RAM[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4717_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0577_),
    .Q(\tms1x00.RAM[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4718_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0578_),
    .Q(\tms1x00.RAM[17][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4719_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0579_),
    .Q(\tms1x00.RAM[17][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4720_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0580_),
    .Q(\tms1x00.RAM[17][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4721_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0581_),
    .Q(\tms1x00.RAM[17][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4722_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0582_),
    .Q(\tms1x00.RAM[29][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4723_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0583_),
    .Q(\tms1x00.RAM[29][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4724_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0584_),
    .Q(\tms1x00.RAM[29][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4725_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0585_),
    .Q(\tms1x00.RAM[29][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4726_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0586_),
    .Q(\tms1x00.RAM[16][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4727_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0587_),
    .Q(\tms1x00.RAM[16][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4728_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0588_),
    .Q(\tms1x00.RAM[16][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4729_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0589_),
    .Q(\tms1x00.RAM[16][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4730_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0590_),
    .Q(\tms1x00.RAM[119][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4731_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0591_),
    .Q(\tms1x00.RAM[119][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4732_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0592_),
    .Q(\tms1x00.RAM[119][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4733_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0593_),
    .Q(\tms1x00.RAM[119][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4734_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0594_),
    .Q(\tms1x00.RAM[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4735_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0595_),
    .Q(\tms1x00.RAM[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4736_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0596_),
    .Q(\tms1x00.RAM[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4737_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0597_),
    .Q(\tms1x00.RAM[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4738_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0598_),
    .Q(\tms1x00.RAM[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4739_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0599_),
    .Q(\tms1x00.RAM[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4740_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0600_),
    .Q(\tms1x00.RAM[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4741_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0601_),
    .Q(\tms1x00.RAM[15][3] ));
 sky130_fd_sc_hd__dfxtp_4 _4742_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0602_),
    .Q(\tms1x00.rom_addr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4743_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0603_),
    .Q(\tms1x00.rom_addr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4744_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_0604_),
    .Q(net52));
 sky130_fd_sc_hd__dfxtp_1 _4745_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_0605_),
    .Q(net53));
 sky130_fd_sc_hd__dfxtp_1 _4746_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_0606_),
    .Q(net54));
 sky130_fd_sc_hd__dfxtp_1 _4747_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0607_),
    .Q(net55));
 sky130_fd_sc_hd__dfxtp_1 _4748_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_0608_),
    .Q(net56));
 sky130_fd_sc_hd__dfxtp_1 _4749_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0609_),
    .Q(net57));
 sky130_fd_sc_hd__dfxtp_1 _4750_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0610_),
    .Q(net58));
 sky130_fd_sc_hd__dfxtp_1 _4751_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0611_),
    .Q(net59));
 sky130_fd_sc_hd__dfxtp_1 _4752_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0612_),
    .Q(\tms1x00.RAM[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4753_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0613_),
    .Q(\tms1x00.RAM[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4754_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0614_),
    .Q(\tms1x00.RAM[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4755_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0615_),
    .Q(\tms1x00.RAM[9][3] ));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_120 (.HI(net120));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_121 (.HI(net121));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_122 (.HI(net122));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_123 (.HI(net123));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_124 (.HI(net124));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_125 (.HI(net125));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_126 (.HI(net126));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_127 (.HI(net127));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_128 (.HI(net128));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_73 (.LO(net73));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_74 (.LO(net74));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_75 (.LO(net75));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_76 (.LO(net76));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_77 (.LO(net77));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_78 (.LO(net78));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_79 (.LO(net79));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_80 (.LO(net80));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_81 (.LO(net81));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_82 (.LO(net82));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_83 (.LO(net83));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_84 (.LO(net84));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_85 (.LO(net85));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_86 (.LO(net86));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_87 (.LO(net87));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_88 (.LO(net88));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_89 (.LO(net89));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_90 (.LO(net90));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_91 (.LO(net91));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_92 (.LO(net92));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_93 (.LO(net93));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_94 (.LO(net94));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_95 (.LO(net95));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_96 (.LO(net96));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_97 (.LO(net97));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_98 (.LO(net98));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_99 (.LO(net99));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_100 (.LO(net100));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_101 (.LO(net101));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_102 (.LO(net102));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_103 (.LO(net103));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_104 (.LO(net104));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_105 (.LO(net105));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_106 (.LO(net106));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_107 (.LO(net107));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_108 (.LO(net108));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_109 (.LO(net109));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_110 (.LO(net110));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_111 (.LO(net111));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_112 (.LO(net112));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_113 (.LO(net113));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_114 (.LO(net114));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_115 (.LO(net115));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_116 (.LO(net116));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_117 (.LO(net117));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_118 (.LO(net118));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_119 (.HI(net119));
 sky130_fd_sc_hd__clkbuf_1 _4813_ (.A(net16),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_2 _4814_ (.A(net17),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_2 _4815_ (.A(net19),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_2 _4816_ (.A(net20),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_2 _4817_ (.A(net21),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_2 _4818_ (.A(net22),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_2 _4819_ (.A(net23),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_2 _4820_ (.A(net24),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_2 _4821_ (.A(net25),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_2 _4822_ (.A(net26),
    .X(net69));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(io_in[6]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(io_in[7]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(io_in[8]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(io_in[9]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(oram_value[0]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(oram_value[10]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(oram_value[1]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(oram_value[2]),
    .X(net8));
 sky130_fd_sc_hd__dlymetal6s2s_1 input9 (.A(oram_value[3]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(oram_value[4]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(oram_value[5]),
    .X(net11));
 sky130_fd_sc_hd__dlymetal6s2s_1 input12 (.A(oram_value[6]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(oram_value[7]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(oram_value[8]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(oram_value[9]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_4 input16 (.A(wb_rst_i),
    .X(net16));
 sky130_fd_sc_hd__dlymetal6s2s_1 input17 (.A(wbs_adr_i[0]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(wbs_adr_i[16]),
    .X(net18));
 sky130_fd_sc_hd__dlymetal6s2s_1 input19 (.A(wbs_adr_i[1]),
    .X(net19));
 sky130_fd_sc_hd__dlymetal6s2s_1 input20 (.A(wbs_adr_i[2]),
    .X(net20));
 sky130_fd_sc_hd__dlymetal6s2s_1 input21 (.A(wbs_adr_i[3]),
    .X(net21));
 sky130_fd_sc_hd__dlymetal6s2s_1 input22 (.A(wbs_adr_i[4]),
    .X(net22));
 sky130_fd_sc_hd__dlymetal6s2s_1 input23 (.A(wbs_adr_i[5]),
    .X(net23));
 sky130_fd_sc_hd__dlymetal6s2s_1 input24 (.A(wbs_adr_i[6]),
    .X(net24));
 sky130_fd_sc_hd__dlymetal6s2s_1 input25 (.A(wbs_adr_i[7]),
    .X(net25));
 sky130_fd_sc_hd__dlymetal6s2s_1 input26 (.A(wbs_adr_i[8]),
    .X(net26));
 sky130_fd_sc_hd__dlymetal6s2s_1 input27 (.A(wbs_we_i),
    .X(net27));
 sky130_fd_sc_hd__buf_2 output28 (.A(net28),
    .X(io_out[10]));
 sky130_fd_sc_hd__buf_2 output29 (.A(net29),
    .X(io_out[11]));
 sky130_fd_sc_hd__buf_2 output30 (.A(net30),
    .X(io_out[12]));
 sky130_fd_sc_hd__buf_2 output31 (.A(net31),
    .X(io_out[13]));
 sky130_fd_sc_hd__buf_2 output32 (.A(net32),
    .X(io_out[14]));
 sky130_fd_sc_hd__buf_2 output33 (.A(net33),
    .X(io_out[15]));
 sky130_fd_sc_hd__buf_2 output34 (.A(net34),
    .X(io_out[16]));
 sky130_fd_sc_hd__buf_2 output35 (.A(net35),
    .X(io_out[17]));
 sky130_fd_sc_hd__buf_2 output36 (.A(net36),
    .X(io_out[18]));
 sky130_fd_sc_hd__buf_2 output37 (.A(net37),
    .X(io_out[19]));
 sky130_fd_sc_hd__buf_2 output38 (.A(net38),
    .X(io_out[20]));
 sky130_fd_sc_hd__buf_2 output39 (.A(net39),
    .X(io_out[21]));
 sky130_fd_sc_hd__buf_2 output40 (.A(net40),
    .X(io_out[22]));
 sky130_fd_sc_hd__buf_2 output41 (.A(net41),
    .X(io_out[23]));
 sky130_fd_sc_hd__buf_2 output42 (.A(net42),
    .X(io_out[24]));
 sky130_fd_sc_hd__buf_2 output43 (.A(net43),
    .X(io_out[25]));
 sky130_fd_sc_hd__buf_2 output44 (.A(net44),
    .X(io_out[26]));
 sky130_fd_sc_hd__buf_2 output45 (.A(net45),
    .X(io_out[27]));
 sky130_fd_sc_hd__buf_2 output46 (.A(net46),
    .X(io_out[28]));
 sky130_fd_sc_hd__buf_2 output47 (.A(net47),
    .X(io_out[29]));
 sky130_fd_sc_hd__buf_2 output48 (.A(net48),
    .X(io_out[30]));
 sky130_fd_sc_hd__buf_2 output49 (.A(net49),
    .X(io_out[31]));
 sky130_fd_sc_hd__buf_2 output50 (.A(net50),
    .X(io_out[32]));
 sky130_fd_sc_hd__buf_2 output51 (.A(net51),
    .X(io_out[33]));
 sky130_fd_sc_hd__buf_2 output52 (.A(net52),
    .X(oram_addr[0]));
 sky130_fd_sc_hd__buf_2 output53 (.A(net53),
    .X(oram_addr[1]));
 sky130_fd_sc_hd__buf_2 output54 (.A(net54),
    .X(oram_addr[2]));
 sky130_fd_sc_hd__buf_2 output55 (.A(net55),
    .X(oram_addr[3]));
 sky130_fd_sc_hd__buf_2 output56 (.A(net56),
    .X(oram_addr[4]));
 sky130_fd_sc_hd__buf_2 output57 (.A(net57),
    .X(oram_addr[5]));
 sky130_fd_sc_hd__buf_2 output58 (.A(net58),
    .X(oram_addr[6]));
 sky130_fd_sc_hd__buf_2 output59 (.A(net59),
    .X(oram_addr[7]));
 sky130_fd_sc_hd__buf_2 output60 (.A(net60),
    .X(oram_csb));
 sky130_fd_sc_hd__buf_2 output61 (.A(net61),
    .X(ram_adrb[0]));
 sky130_fd_sc_hd__buf_2 output62 (.A(net62),
    .X(ram_adrb[1]));
 sky130_fd_sc_hd__buf_2 output63 (.A(net63),
    .X(ram_adrb[2]));
 sky130_fd_sc_hd__buf_2 output64 (.A(net64),
    .X(ram_adrb[3]));
 sky130_fd_sc_hd__buf_2 output65 (.A(net65),
    .X(ram_adrb[4]));
 sky130_fd_sc_hd__buf_2 output66 (.A(net66),
    .X(ram_adrb[5]));
 sky130_fd_sc_hd__buf_2 output67 (.A(net67),
    .X(ram_adrb[6]));
 sky130_fd_sc_hd__buf_2 output68 (.A(net68),
    .X(ram_adrb[7]));
 sky130_fd_sc_hd__buf_2 output69 (.A(net69),
    .X(ram_adrb[8]));
 sky130_fd_sc_hd__buf_2 output70 (.A(net70),
    .X(ram_csb));
 sky130_fd_sc_hd__buf_2 output71 (.A(net71),
    .X(ram_web));
 sky130_fd_sc_hd__conb_1 wrapped_tms1x00_72 (.LO(net72));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_21_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_23_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_25_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_26_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_28_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_29_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_32_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_33_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_34_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_37_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__2510__S1 (.DIODE(_0001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2206__A (.DIODE(_0001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2198__A (.DIODE(_0001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2169__A (.DIODE(_0001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2164__A (.DIODE(_0001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2149__A (.DIODE(_0001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2126__A (.DIODE(_0001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2528__B1 (.DIODE(_0003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2385__B1 (.DIODE(_0003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2208__A (.DIODE(_0003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2177__A (.DIODE(_0003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2158__A (.DIODE(_0003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2144__A (.DIODE(_0003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2591__C1 (.DIODE(_0004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2534__A1 (.DIODE(_0004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2522__B1 (.DIODE(_0004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2310__C1 (.DIODE(_0004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2222__A (.DIODE(_0004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2163__A (.DIODE(_0004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2161__A (.DIODE(_0004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2211__A (.DIODE(_0005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2125__A (.DIODE(_0005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2594__A1 (.DIODE(_0006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2593__A (.DIODE(_0006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2448__B1 (.DIODE(_0006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2345__C1 (.DIODE(_0006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2256__A (.DIODE(_0006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2225__C1 (.DIODE(_0006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3974__A1 (.DIODE(_0616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3953__A1 (.DIODE(_0616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3806__B (.DIODE(_0616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3797__B (.DIODE(_0616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3796__B (.DIODE(_0616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3792__C_N (.DIODE(_0616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3735__A0 (.DIODE(_0616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2113__C (.DIODE(_0616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2102__C (.DIODE(_0616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2081__A0 (.DIODE(_0616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3893__C (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3833__A (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3799__A (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3775__A (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2119__A (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2079__A (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3739__S (.DIODE(_0622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3737__S (.DIODE(_0622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3735__S (.DIODE(_0622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2098__S (.DIODE(_0622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2096__S (.DIODE(_0622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2094__S (.DIODE(_0622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2092__S (.DIODE(_0622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2088__S (.DIODE(_0622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2085__S (.DIODE(_0622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2081__S (.DIODE(_0622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3981__A1 (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3958__A1 (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3806__A (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3796__C_N (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3793__B (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3792__B (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3737__A0 (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2113__B (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2102__B (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2085__A0 (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3988__A1 (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3806__C_N (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3797__A (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3796__A (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3793__A (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3792__A (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3739__A0 (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2113__A (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2102__A (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2088__A0 (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3966__A1 (.DIODE(_0629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3844__A1 (.DIODE(_0629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3841__A1 (.DIODE(_0629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3838__A1 (.DIODE(_0629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3835__A1 (.DIODE(_0629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3831__A1 (.DIODE(_0629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3829__A1 (.DIODE(_0629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3827__A1 (.DIODE(_0629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3825__A1 (.DIODE(_0629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2091__A (.DIODE(_0629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3993__A1 (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3843__A (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3840__A (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3837__A (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3809__A1 (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3800__A1 (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3795__A1 (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3741__A0 (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2120__A1 (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2092__A0 (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4000__A (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3941__A1 (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3890__A0 (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3862__A2 (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3859__A1 (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3856__A1 (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3853__A1 (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3850__A1 (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3791__A1 (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2109__A (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3997__A (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3949__B (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3938__A1 (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3886__A0 (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3847__D (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3788__A1 (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2596__B (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2497__A (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2280__A2 (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2109__B (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3836__A2 (.DIODE(_0642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3832__B (.DIODE(_0642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3822__B (.DIODE(_0642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3817__B (.DIODE(_0642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3812__B (.DIODE(_0642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3803__B (.DIODE(_0642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2110__A (.DIODE(_0642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3831__A2 (.DIODE(_0649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3825__A3 (.DIODE(_0649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3821__A2 (.DIODE(_0649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3816__A2 (.DIODE(_0649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3811__A2 (.DIODE(_0649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3802__A2 (.DIODE(_0649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2117__A (.DIODE(_0649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4004__C1 (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4002__C1 (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3999__C1 (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3993__C1 (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3988__C1 (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3981__C1 (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3974__C1 (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3863__C1 (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3795__C1 (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2120__C1 (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2592__C1 (.DIODE(_0657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2572__C1 (.DIODE(_0657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2534__B1 (.DIODE(_0657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2513__B1 (.DIODE(_0657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2473__B1 (.DIODE(_0657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2448__A1 (.DIODE(_0657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2370__B1 (.DIODE(_0657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2345__A1 (.DIODE(_0657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2255__B1 (.DIODE(_0657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2225__A1 (.DIODE(_0657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2527__S1 (.DIODE(_0658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2519__S1 (.DIODE(_0658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2440__S1 (.DIODE(_0658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2384__S1 (.DIODE(_0658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2337__S1 (.DIODE(_0658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2235__A (.DIODE(_0658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2215__S1 (.DIODE(_0658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2156__A (.DIODE(_0658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2142__A (.DIODE(_0658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2127__A (.DIODE(_0658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2524__A (.DIODE(_0659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2518__S1 (.DIODE(_0659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2509__S1 (.DIODE(_0659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2506__A1 (.DIODE(_0659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2504__A_N (.DIODE(_0659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2327__A (.DIODE(_0659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2252__S1 (.DIODE(_0659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2226__A (.DIODE(_0659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2132__A (.DIODE(_0659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2128__A (.DIODE(_0659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2568__A1 (.DIODE(_0660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2526__A (.DIODE(_0660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2475__A (.DIODE(_0660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2428__A (.DIODE(_0660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2406__A1 (.DIODE(_0660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2372__A (.DIODE(_0660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2325__A (.DIODE(_0660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2303__A1 (.DIODE(_0660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2195__A (.DIODE(_0660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2138__A1 (.DIODE(_0660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2527__S0 (.DIODE(_0661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2523__S (.DIODE(_0661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2505__S (.DIODE(_0661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2440__S0 (.DIODE(_0661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2402__S (.DIODE(_0661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2384__S0 (.DIODE(_0661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2337__S0 (.DIODE(_0661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2215__S0 (.DIODE(_0661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2155__A (.DIODE(_0661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2130__S (.DIODE(_0661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2562__A1 (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2458__A1 (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2423__A1 (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2405__A (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2355__A1 (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2320__A1 (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2302__A (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2239__A1 (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2184__A1 (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2136__A (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2519__S0 (.DIODE(_0665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2510__S0 (.DIODE(_0665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2503__S (.DIODE(_0665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2299__S (.DIODE(_0665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2265__A (.DIODE(_0665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2181__A (.DIODE(_0665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2171__A (.DIODE(_0665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2166__A (.DIODE(_0665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2141__A (.DIODE(_0665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2134__A (.DIODE(_0665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2575__S (.DIODE(_0666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2565__S (.DIODE(_0666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2561__S (.DIODE(_0666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2543__S (.DIODE(_0666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2518__S0 (.DIODE(_0666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2457__S (.DIODE(_0666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2420__S (.DIODE(_0666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2404__S (.DIODE(_0666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2179__S (.DIODE(_0666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2135__S (.DIODE(_0666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2512__A1 (.DIODE(_0669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2508__B2 (.DIODE(_0669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2490__A (.DIODE(_0669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2483__A1 (.DIODE(_0669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2436__A1 (.DIODE(_0669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2406__C1 (.DIODE(_0669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2303__C1 (.DIODE(_0669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2274__A (.DIODE(_0669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2267__A1 (.DIODE(_0669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2138__C1 (.DIODE(_0669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2162__A1 (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2528__A1 (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2441__A1 (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2385__A1 (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2338__A1 (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2329__A1 (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2216__A1 (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2200__A1 (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2176__A (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2146__A (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2140__A (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2529__A1 (.DIODE(_0672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2480__A1 (.DIODE(_0672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2468__A1 (.DIODE(_0672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2433__A1 (.DIODE(_0672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2408__A1 (.DIODE(_0672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2377__A1 (.DIODE(_0672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2330__A1 (.DIODE(_0672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2305__A1 (.DIODE(_0672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2201__A1 (.DIODE(_0672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2145__A1 (.DIODE(_0672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2539__S0 (.DIODE(_0673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2474__S (.DIODE(_0673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2464__S (.DIODE(_0673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2427__S (.DIODE(_0673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2407__S0 (.DIODE(_0673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2361__S (.DIODE(_0673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2304__S0 (.DIODE(_0673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2257__S (.DIODE(_0673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2246__S (.DIODE(_0673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2143__S0 (.DIODE(_0673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2539__S1 (.DIODE(_0674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2453__S1 (.DIODE(_0674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2411__S1 (.DIODE(_0674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2407__S1 (.DIODE(_0674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2374__A (.DIODE(_0674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2350__S1 (.DIODE(_0674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2308__S1 (.DIODE(_0674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2304__S1 (.DIODE(_0674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2197__A (.DIODE(_0674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2143__S1 (.DIODE(_0674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2521__C1 (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2512__C1 (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2483__B1 (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2467__B1 (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2408__B1 (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2364__B1 (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2305__B1 (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2267__B1 (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2249__B1 (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2145__B1 (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2578__B2 (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2564__B2 (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2546__B2 (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2533__A1 (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2460__B2 (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2410__A (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2357__B2 (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2322__B2 (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2307__A (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2152__A (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2580__S0 (.DIODE(_0679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2444__S0 (.DIODE(_0679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2388__S0 (.DIODE(_0679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2341__S0 (.DIODE(_0679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2328__S0 (.DIODE(_0679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2326__S (.DIODE(_0679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2220__S0 (.DIODE(_0679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2199__S0 (.DIODE(_0679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2196__S (.DIODE(_0679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2148__A (.DIODE(_0679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2563__S0 (.DIODE(_0680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2545__S0 (.DIODE(_0680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2530__S0 (.DIODE(_0680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2459__S0 (.DIODE(_0680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2409__S0 (.DIODE(_0680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2356__S0 (.DIODE(_0680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2321__S0 (.DIODE(_0680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2306__S0 (.DIODE(_0680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2240__S0 (.DIODE(_0680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2151__S0 (.DIODE(_0680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2587__S1 (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2531__S1 (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2438__S1 (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2431__S1 (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2382__S1 (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2375__S1 (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2335__S1 (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2271__S1 (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2213__S1 (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2150__A (.DIODE(_0681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2579__S1 (.DIODE(_0682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2569__S1 (.DIODE(_0682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2536__A_N (.DIODE(_0682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2451__A_N (.DIODE(_0682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2424__S1 (.DIODE(_0682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2331__S1 (.DIODE(_0682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2240__S1 (.DIODE(_0682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2203__S1 (.DIODE(_0682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2187__S1 (.DIODE(_0682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2151__S1 (.DIODE(_0682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2152__B (.DIODE(_0683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2521__A1 (.DIODE(_0686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2515__A (.DIODE(_0686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2471__A1 (.DIODE(_0686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2452__C1 (.DIODE(_0686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2412__A1 (.DIODE(_0686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2368__A1 (.DIODE(_0686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2309__A1 (.DIODE(_0686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2270__A (.DIODE(_0686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2253__A1 (.DIODE(_0686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2160__A1 (.DIODE(_0686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2577__S0 (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2453__S0 (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2418__S0 (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2411__S0 (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2350__S0 (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2315__S0 (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2308__S0 (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2233__S0 (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2175__S0 (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2157__S0 (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2577__S1 (.DIODE(_0688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2545__S1 (.DIODE(_0688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2530__S1 (.DIODE(_0688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2477__A (.DIODE(_0688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2430__A (.DIODE(_0688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2418__S1 (.DIODE(_0688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2315__S1 (.DIODE(_0688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2233__S1 (.DIODE(_0688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2175__S1 (.DIODE(_0688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2157__S1 (.DIODE(_0688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2578__C1 (.DIODE(_0691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2508__C1 (.DIODE(_0691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2471__B1 (.DIODE(_0691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2412__B1 (.DIODE(_0691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2368__B1 (.DIODE(_0691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2309__B1 (.DIODE(_0691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2276__B1 (.DIODE(_0691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2262__B1 (.DIODE(_0691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2253__B1 (.DIODE(_0691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2160__B1 (.DIODE(_0691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2494__A1 (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2473__A1 (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2447__A1 (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2413__C1 (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2391__A1 (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2370__A1 (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2344__A1 (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2278__A1 (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2224__A1 (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2162__C1 (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2589__S1 (.DIODE(_0696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2585__S1 (.DIODE(_0696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2491__S1 (.DIODE(_0696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2478__S1 (.DIODE(_0696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2442__S1 (.DIODE(_0696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2386__S1 (.DIODE(_0696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2339__S1 (.DIODE(_0696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2275__S1 (.DIODE(_0696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2217__S1 (.DIODE(_0696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2165__A (.DIODE(_0696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2574__A_N (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2542__A_N (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2538__A1 (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2434__S1 (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2415__A_N (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2378__S1 (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2348__A_N (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2312__A_N (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2231__A_N (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2168__A_N (.DIODE(_0697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2537__S (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2514__S0 (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2450__S (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2435__S0 (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2414__S (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2347__S (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2311__S (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2269__S0 (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2230__S (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2167__S (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2514__S1 (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2489__S1 (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2482__S1 (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2470__S1 (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2435__S1 (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2367__S1 (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2273__S1 (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2269__S1 (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2266__S1 (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2170__A (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2576__A1 (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2566__A_N (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2556__S1 (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2544__A1 (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2421__A_N (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2417__A1 (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2314__A1 (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2251__S1 (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2180__A_N (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2174__A1 (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2551__S (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2509__S0 (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2416__S (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2367__S0 (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2317__S (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2313__S (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2301__S (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2252__S0 (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2236__S (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2172__S (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2576__B1 (.DIODE(_0705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2544__B1 (.DIODE(_0705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2538__B1 (.DIODE(_0705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2445__A1 (.DIODE(_0705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2417__B1 (.DIODE(_0705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2389__A1 (.DIODE(_0705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2342__A1 (.DIODE(_0705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2314__B1 (.DIODE(_0705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2202__A (.DIODE(_0705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2174__B1 (.DIODE(_0705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2540__B2 (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2454__A (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2419__B2 (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2365__A1 (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2351__A (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2316__B2 (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2263__A1 (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2250__A1 (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2234__A (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2178__B2 (.DIODE(_0708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2567__S (.DIODE(_0713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2525__S (.DIODE(_0713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2422__S (.DIODE(_0713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2371__S (.DIODE(_0713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2354__S (.DIODE(_0713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2324__S (.DIODE(_0713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2319__S (.DIODE(_0713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2238__S (.DIODE(_0713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2194__S (.DIODE(_0713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2182__S (.DIODE(_0713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2590__A1 (.DIODE(_0715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2568__B1 (.DIODE(_0715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2532__A1 (.DIODE(_0715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2492__A1 (.DIODE(_0715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2486__A (.DIODE(_0715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2439__A (.DIODE(_0715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2336__A (.DIODE(_0715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2276__A1 (.DIODE(_0715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2214__A (.DIODE(_0715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2184__B1 (.DIODE(_0715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2587__S0 (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2583__S0 (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2531__S0 (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2487__S0 (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2438__S0 (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2431__S0 (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2382__S0 (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2375__S0 (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2271__S0 (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2186__A (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2579__S0 (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2569__S0 (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2481__S0 (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2469__S0 (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2434__S0 (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2424__S0 (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2378__S0 (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2331__S0 (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2203__S0 (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2187__S0 (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2192__B1 (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2588__A (.DIODE(_0720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2586__A1 (.DIODE(_0720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2488__A1 (.DIODE(_0720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2443__A (.DIODE(_0720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2432__A1 (.DIODE(_0720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2387__A (.DIODE(_0720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2376__A1 (.DIODE(_0720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2340__A (.DIODE(_0720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2272__A1 (.DIODE(_0720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2189__A (.DIODE(_0720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2582__A1 (.DIODE(_0721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2570__B2 (.DIODE(_0721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2558__A1 (.DIODE(_0721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2554__A1 (.DIODE(_0721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2472__A1 (.DIODE(_0721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2425__B2 (.DIODE(_0721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2369__A1 (.DIODE(_0721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2254__A1 (.DIODE(_0721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2241__B2 (.DIODE(_0721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2192__B2 (.DIODE(_0721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2590__B1 (.DIODE(_0722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2492__B1 (.DIODE(_0722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2479__B1 (.DIODE(_0722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2432__B1 (.DIODE(_0722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2376__B1 (.DIODE(_0722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2342__B1 (.DIODE(_0722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2329__B1 (.DIODE(_0722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2221__B1 (.DIODE(_0722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2200__B1 (.DIODE(_0722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2191__A (.DIODE(_0722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2570__C1 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2557__B1 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2546__C1 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2522__A1 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2461__A1 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2425__C1 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2358__A1 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2322__C1 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2242__A1 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2192__C1 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2583__S1 (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2580__S1 (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2487__S1 (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2444__S1 (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2388__S1 (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2341__S1 (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2328__S1 (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2243__A (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2220__S1 (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2199__S1 (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2557__A1 (.DIODE(_0734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2553__C1 (.DIODE(_0734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2484__A1 (.DIODE(_0734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2437__A1 (.DIODE(_0734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2381__A1 (.DIODE(_0734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2349__C1 (.DIODE(_0734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2334__A1 (.DIODE(_0734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2268__A1 (.DIODE(_0734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2232__C1 (.DIODE(_0734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2210__A1 (.DIODE(_0734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2517__A (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2479__A1 (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2467__A1 (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2380__A1 (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2364__A1 (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2333__A1 (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2262__A1 (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2249__A1 (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2218__A (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2209__A1 (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2589__S0 (.DIODE(_0737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2535__S (.DIODE(_0737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2476__S (.DIODE(_0737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2466__S0 (.DIODE(_0737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2363__S0 (.DIODE(_0737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2332__S0 (.DIODE(_0737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2275__S0 (.DIODE(_0737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2261__S0 (.DIODE(_0737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2217__S0 (.DIODE(_0737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2207__S0 (.DIODE(_0737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2516__S1 (.DIODE(_0738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2507__S1 (.DIODE(_0738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2485__S1 (.DIODE(_0738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2466__S1 (.DIODE(_0738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2379__S1 (.DIODE(_0738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2363__S1 (.DIODE(_0738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2332__S1 (.DIODE(_0738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2261__S1 (.DIODE(_0738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2248__S1 (.DIODE(_0738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2207__S1 (.DIODE(_0738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2494__B1 (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2447__C1 (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2391__C1 (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2344__B1 (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2278__B1 (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2224__B1 (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2585__S0 (.DIODE(_0744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2491__S0 (.DIODE(_0744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2478__S0 (.DIODE(_0744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2442__S0 (.DIODE(_0744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2429__S (.DIODE(_0744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2386__S0 (.DIODE(_0744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2373__S (.DIODE(_0744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2339__S0 (.DIODE(_0744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2335__S0 (.DIODE(_0744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2213__S0 (.DIODE(_0744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2216__A2 (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2584__A (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2581__A (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2562__B1 (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2458__B1 (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2423__B1 (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2383__A (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2355__B1 (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2320__B1 (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2239__B1 (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2221__A1 (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2592__A1 (.DIODE(_0754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2513__A1 (.DIODE(_0754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2493__C1 (.DIODE(_0754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2446__C1 (.DIODE(_0754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2390__C1 (.DIODE(_0754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2343__C1 (.DIODE(_0754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2277__C1 (.DIODE(_0754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2223__C1 (.DIODE(_0754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3945__A (.DIODE(_0757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2280__B1 (.DIODE(_0757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2555__S1 (.DIODE(_0758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2553__A1 (.DIODE(_0758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2549__S1 (.DIODE(_0758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2465__A (.DIODE(_0758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2452__A1 (.DIODE(_0758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2362__A (.DIODE(_0758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2349__A1 (.DIODE(_0758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2258__A (.DIODE(_0758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2247__A (.DIODE(_0758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2232__A1 (.DIODE(_0758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2516__S0 (.DIODE(_0759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2507__S0 (.DIODE(_0759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2485__S0 (.DIODE(_0759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2462__S (.DIODE(_0759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2379__S0 (.DIODE(_0759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2359__S (.DIODE(_0759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2259__S (.DIODE(_0759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2248__S0 (.DIODE(_0759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2244__S (.DIODE(_0759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2228__A (.DIODE(_0759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2556__S0 (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2555__S0 (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2550__S (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2549__S0 (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2449__S (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2366__S0 (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2346__S (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2264__S0 (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2251__S0 (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2229__S (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2560__A_N (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2552__A_N (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2481__S1 (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2469__S1 (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2456__A_N (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2366__S1 (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2353__A_N (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2318__A_N (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2264__S1 (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2237__A_N (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2563__S1 (.DIODE(_0775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2463__A (.DIODE(_0775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2459__S1 (.DIODE(_0775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2409__S1 (.DIODE(_0775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2360__A (.DIODE(_0775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2356__S1 (.DIODE(_0775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2321__S1 (.DIODE(_0775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2306__S1 (.DIODE(_0775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2260__A (.DIODE(_0775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2245__A (.DIODE(_0775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2245__B_N (.DIODE(_0776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2250__A3 (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2250__B1 (.DIODE(_0781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2254__A2 (.DIODE(_0783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2268__A2 (.DIODE(_0796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2573__S (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2559__S (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2541__S (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2489__S0 (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2482__S0 (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2470__S0 (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2455__S (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2352__S (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2273__S0 (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2266__S0 (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2277__A2 (.DIODE(_0804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2274__B (.DIODE(_0805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3945__B (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2280__B2 (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3695__A (.DIODE(_0820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3547__A (.DIODE(_0820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3417__A (.DIODE(_0820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3305__A (.DIODE(_0820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3151__A (.DIODE(_0820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3036__A (.DIODE(_0820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2914__A (.DIODE(_0820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2726__A (.DIODE(_0820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2602__A (.DIODE(_0820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2289__A (.DIODE(_0820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2718__A0 (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2709__A0 (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2699__A0 (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2690__A0 (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2680__A0 (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2670__A0 (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2659__A0 (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2649__A0 (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2636__A0 (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2297__A0 (.DIODE(_0821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2972__A (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2954__A (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2945__A (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2896__A (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2887__A (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2878__A (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2291__A (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2990__A (.DIODE(_0823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2981__A (.DIODE(_0823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2858__A (.DIODE(_0823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2848__A (.DIODE(_0823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2839__A (.DIODE(_0823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2830__A (.DIODE(_0823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2815__A (.DIODE(_0823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2804__A (.DIODE(_0823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2635__A (.DIODE(_0823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2296__A (.DIODE(_0823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3051__A (.DIODE(_0825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3038__A (.DIODE(_0825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3027__A (.DIODE(_0825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2793__A (.DIODE(_0825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2782__B (.DIODE(_0825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2647__B (.DIODE(_0825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2633__A_N (.DIODE(_0825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2605__B (.DIODE(_0825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2294__C (.DIODE(_0825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3708__A (.DIODE(_0827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3529__A (.DIODE(_0827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3439__A (.DIODE(_0827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3296__A (.DIODE(_0827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3251__A (.DIODE(_0827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2905__A (.DIODE(_0827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2689__A (.DIODE(_0827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2296__B (.DIODE(_0827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2307__B (.DIODE(_0837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2316__B1 (.DIODE(_0846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2322__B1 (.DIODE(_0852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2338__A2 (.DIODE(_0868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3956__A (.DIODE(_0876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2394__A1 (.DIODE(_0876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2360__B_N (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2365__A3 (.DIODE(_0893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2365__B1 (.DIODE(_0895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2369__A2 (.DIODE(_0897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2381__A2 (.DIODE(_0909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2381__B1 (.DIODE(_0911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2385__A2 (.DIODE(_0915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2387__B (.DIODE(_0917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2389__A2 (.DIODE(_0919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3956__B (.DIODE(_0923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2394__A2 (.DIODE(_0923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4013__A (.DIODE(_0926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4003__A2 (.DIODE(_0926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3994__A (.DIODE(_0926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3968__C_N (.DIODE(_0926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3957__A1 (.DIODE(_0926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3935__A1 (.DIODE(_0926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3882__A0 (.DIODE(_0926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3847__A_N (.DIODE(_0926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3783__A0 (.DIODE(_0926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2396__A1 (.DIODE(_0926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3699__A (.DIODE(_0929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3551__A (.DIODE(_0929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3421__A (.DIODE(_0929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3309__A (.DIODE(_0929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3155__A (.DIODE(_0929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3041__A (.DIODE(_0929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2918__A (.DIODE(_0929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2731__A (.DIODE(_0929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2611__A (.DIODE(_0929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2399__A (.DIODE(_0929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2720__A0 (.DIODE(_0930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2711__A0 (.DIODE(_0930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2701__A0 (.DIODE(_0930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2692__A0 (.DIODE(_0930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2682__A0 (.DIODE(_0930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2672__A0 (.DIODE(_0930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2661__A0 (.DIODE(_0930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2651__A0 (.DIODE(_0930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2638__A0 (.DIODE(_0930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2400__A0 (.DIODE(_0930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2413__A1 (.DIODE(_0936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2410__B (.DIODE(_0939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2419__B1 (.DIODE(_0948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2425__B1 (.DIODE(_0954_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2441__A2 (.DIODE(_0970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3960__A (.DIODE(_0978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2496__A1 (.DIODE(_0978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2463__B_N (.DIODE(_0992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2465__B (.DIODE(_0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2468__B1 (.DIODE(_0997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2472__A2 (.DIODE(_0999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2484__A2 (.DIODE(_1011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2488__A2 (.DIODE(_1017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2490__B (.DIODE(_1019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2492__A2 (.DIODE(_1021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3960__B (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2496__A2 (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3702__A (.DIODE(_1029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3554__A (.DIODE(_1029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3424__A (.DIODE(_1029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3312__A (.DIODE(_1029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3158__A (.DIODE(_1029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3044__A (.DIODE(_1029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2921__A (.DIODE(_1029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2734__A (.DIODE(_1029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2614__A (.DIODE(_1029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2500__A (.DIODE(_1029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2722__A0 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2713__A0 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2703__A0 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2694__A0 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2684__A0 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2674__A0 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2663__A0 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2653__A0 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2640__A0 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2501__A0 (.DIODE(_1030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2521__A2 (.DIODE(_1047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2520__B (.DIODE(_1048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2533__A2 (.DIODE(_1059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2554__A2 (.DIODE(_1078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2554__B1 (.DIODE(_1082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2558__A2 (.DIODE(_1084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2578__A1 (.DIODE(_1103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2582__A2 (.DIODE(_1108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2588__B (.DIODE(_1116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3965__A (.DIODE(_1123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2597__B1 (.DIODE(_1123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3705__A (.DIODE(_1127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3557__A (.DIODE(_1127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3427__A (.DIODE(_1127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3315__A (.DIODE(_1127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3161__A (.DIODE(_1127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3047__A (.DIODE(_1127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2924__A (.DIODE(_1127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2737__A (.DIODE(_1127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2617__A (.DIODE(_1127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2599__A (.DIODE(_1127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2724__A0 (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2715__A0 (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2705__A0 (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2696__A0 (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2686__A0 (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2676__A0 (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2665__A0 (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2655__A0 (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2642__A0 (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2600__A0 (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4105__A0 (.DIODE(_1130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4096__A0 (.DIODE(_1130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2805__A1 (.DIODE(_1130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2785__A1 (.DIODE(_1130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2774__A1 (.DIODE(_1130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2765__A1 (.DIODE(_1130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2752__A1 (.DIODE(_1130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2741__A1 (.DIODE(_1130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2625__A1 (.DIODE(_1130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2609__A1 (.DIODE(_1130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3726__A (.DIODE(_1131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3717__A (.DIODE(_1131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3708__B (.DIODE(_1131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3696__A (.DIODE(_1131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3686__A (.DIODE(_1131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3659__A (.DIODE(_1131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2604__A (.DIODE(_1131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2795__A (.DIODE(_1132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2784__A (.DIODE(_1132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2773__A (.DIODE(_1132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2751__A (.DIODE(_1132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2740__A (.DIODE(_1132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2728__A (.DIODE(_1132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2717__A (.DIODE(_1132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2708__A (.DIODE(_1132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2698__A (.DIODE(_1132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2608__A (.DIODE(_1132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4134__A (.DIODE(_1135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3632__A (.DIODE(_1135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3457__A (.DIODE(_1135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3278__A (.DIODE(_1135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3182__A (.DIODE(_1135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2804__B (.DIODE(_1135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2608__B (.DIODE(_1135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4107__A0 (.DIODE(_1138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4098__A0 (.DIODE(_1138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2807__A1 (.DIODE(_1138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2787__A1 (.DIODE(_1138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2776__A1 (.DIODE(_1138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2767__A1 (.DIODE(_1138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2754__A1 (.DIODE(_1138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2743__A1 (.DIODE(_1138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2627__A1 (.DIODE(_1138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2612__A1 (.DIODE(_1138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4109__A0 (.DIODE(_1140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4100__A0 (.DIODE(_1140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2809__A1 (.DIODE(_1140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2789__A1 (.DIODE(_1140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2778__A1 (.DIODE(_1140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2769__A1 (.DIODE(_1140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2756__A1 (.DIODE(_1140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2745__A1 (.DIODE(_1140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2629__A1 (.DIODE(_1140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2615__A1 (.DIODE(_1140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4111__A0 (.DIODE(_1142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4102__A0 (.DIODE(_1142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2811__A1 (.DIODE(_1142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2791__A1 (.DIODE(_1142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2780__A1 (.DIODE(_1142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2771__A1 (.DIODE(_1142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2758__A1 (.DIODE(_1142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2747__A1 (.DIODE(_1142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2631__A1 (.DIODE(_1142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2618__A1 (.DIODE(_1142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3475__A (.DIODE(_1145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3466__A (.DIODE(_1145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3457__B (.DIODE(_1145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3448__A (.DIODE(_1145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3418__A (.DIODE(_1145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3408__A (.DIODE(_1145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3381__A (.DIODE(_1145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3363__A (.DIODE(_1145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2679__A (.DIODE(_1145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2624__A (.DIODE(_1145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3614__A (.DIODE(_1147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3345__A (.DIODE(_1147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3164__A (.DIODE(_1147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3060__A (.DIODE(_1147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3017__A (.DIODE(_1147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2981__B (.DIODE(_1147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2740__B (.DIODE(_1147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2624__B (.DIODE(_1147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4068__A (.DIODE(_1154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4023__A (.DIODE(_1154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3650__A (.DIODE(_1154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3502__B (.DIODE(_1154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3327__A (.DIODE(_1154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2999__A (.DIODE(_1154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2717__B (.DIODE(_1154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2635__B (.DIODE(_1154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3677__A (.DIODE(_1160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3650__B (.DIODE(_1160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3605__A (.DIODE(_1160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3596__A (.DIODE(_1160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3578__A (.DIODE(_1160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3529__B (.DIODE(_1160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2645__A (.DIODE(_1160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3641__A (.DIODE(_1161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3632__B (.DIODE(_1161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3623__A (.DIODE(_1161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3614__B (.DIODE(_1161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3569__A (.DIODE(_1161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3560__A (.DIODE(_1161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3548__A (.DIODE(_1161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3538__A (.DIODE(_1161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2658__A (.DIODE(_1161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2648__A (.DIODE(_1161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3686__B (.DIODE(_1163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3520__A (.DIODE(_1163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3418__B (.DIODE(_1163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3318__A (.DIODE(_1163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3133__A (.DIODE(_1163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3078__A (.DIODE(_1163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2848__B (.DIODE(_1163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2648__B (.DIODE(_1163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4104__A (.DIODE(_1169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3484__B (.DIODE(_1169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3390__A (.DIODE(_1169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3215__A (.DIODE(_1169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2945__B (.DIODE(_1169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2698__B (.DIODE(_1169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2669__A (.DIODE(_1169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2658__B (.DIODE(_1169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3078__B (.DIODE(_1175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3051__B (.DIODE(_1175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3038__C (.DIODE(_1175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3027__B (.DIODE(_1175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3017__B (.DIODE(_1175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2999__B (.DIODE(_1175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2668__A (.DIODE(_1175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4086__A (.DIODE(_1176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3096__A (.DIODE(_1176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3087__A (.DIODE(_1176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3069__A (.DIODE(_1176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3008__A (.DIODE(_1176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2936__A (.DIODE(_1176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2927__A (.DIODE(_1176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2915__A (.DIODE(_1176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2905__B (.DIODE(_1176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2669__B (.DIODE(_1176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4059__A (.DIODE(_1182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3726__B (.DIODE(_1182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3548__B (.DIODE(_1182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3269__A (.DIODE(_1182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3105__A (.DIODE(_1182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2927__B (.DIODE(_1182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2887__B (.DIODE(_1182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2679__B (.DIODE(_1182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4077__A (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4068__B (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4059__B (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3215__B (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3133__B (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3114__A (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2689__B (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4050__A (.DIODE(_1199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3677__B (.DIODE(_1199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3493__B (.DIODE(_1199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3399__A (.DIODE(_1199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3224__B (.DIODE(_1199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3096__B (.DIODE(_1199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2954__B (.DIODE(_1199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2708__B (.DIODE(_1199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2906__A0 (.DIODE(_1210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2897__A0 (.DIODE(_1210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2888__A0 (.DIODE(_1210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2879__A0 (.DIODE(_1210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2869__A0 (.DIODE(_1210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2859__A0 (.DIODE(_1210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2849__A0 (.DIODE(_1210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2840__A0 (.DIODE(_1210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2796__A0 (.DIODE(_1210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2729__A0 (.DIODE(_1210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4095__A (.DIODE(_1211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3605__B (.DIODE(_1211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3511__B (.DIODE(_1211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3336__A (.DIODE(_1211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3152__B (.DIODE(_1211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3008__B (.DIODE(_1211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2972__B (.DIODE(_1211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2728__B (.DIODE(_1211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2908__A0 (.DIODE(_1214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2899__A0 (.DIODE(_1214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2890__A0 (.DIODE(_1214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2881__A0 (.DIODE(_1214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2871__A0 (.DIODE(_1214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2861__A0 (.DIODE(_1214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2851__A0 (.DIODE(_1214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2842__A0 (.DIODE(_1214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2798__A0 (.DIODE(_1214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2732__A0 (.DIODE(_1214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2910__A0 (.DIODE(_1216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2901__A0 (.DIODE(_1216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2892__A0 (.DIODE(_1216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2883__A0 (.DIODE(_1216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2873__A0 (.DIODE(_1216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2863__A0 (.DIODE(_1216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2853__A0 (.DIODE(_1216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2844__A0 (.DIODE(_1216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2800__A0 (.DIODE(_1216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2735__A0 (.DIODE(_1216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2912__A0 (.DIODE(_1218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2903__A0 (.DIODE(_1218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2894__A0 (.DIODE(_1218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2885__A0 (.DIODE(_1218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2875__A0 (.DIODE(_1218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2865__A0 (.DIODE(_1218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2855__A0 (.DIODE(_1218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2846__A0 (.DIODE(_1218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2802__A0 (.DIODE(_1218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2738__A0 (.DIODE(_1218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3623__B (.DIODE(_1226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3448__B (.DIODE(_1226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3354__A (.DIODE(_1226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3173__B (.DIODE(_1226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2990__B (.DIODE(_1226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2963__A (.DIODE(_1226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2751__B (.DIODE(_1226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4104__B (.DIODE(_1232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4095__B (.DIODE(_1232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4050__B (.DIODE(_1232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4023__B (.DIODE(_1232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3520__B (.DIODE(_1232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3296__B (.DIODE(_1232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2761__A (.DIODE(_1232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4134__B (.DIODE(_1233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3668__A (.DIODE(_1233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3587__A (.DIODE(_1233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3372__A (.DIODE(_1233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3233__A (.DIODE(_1233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3105__B (.DIODE(_1233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3060__B (.DIODE(_1233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2963__B (.DIODE(_1233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2868__A (.DIODE(_1233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2764__A (.DIODE(_1233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3641__B (.DIODE(_1235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3466__B (.DIODE(_1235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3287__A (.DIODE(_1235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3192__B (.DIODE(_1235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2815__B (.DIODE(_1235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2773__B (.DIODE(_1235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2764__B (.DIODE(_1235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4086__B (.DIODE(_1247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4041__A (.DIODE(_1247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3668__B (.DIODE(_1247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3569__B (.DIODE(_1247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3475__B (.DIODE(_1247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3115__B (.DIODE(_1247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2830__B (.DIODE(_1247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2784__B (.DIODE(_1247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3587__B (.DIODE(_1254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3578__B (.DIODE(_1254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3408__B (.DIODE(_1254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3306__A (.DIODE(_1254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3124__B (.DIODE(_1254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3069__B (.DIODE(_1254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2839__B (.DIODE(_1254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2795__B (.DIODE(_1254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4135__A1 (.DIODE(_1265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4087__A1 (.DIODE(_1265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4042__A1 (.DIODE(_1265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3669__A1 (.DIODE(_1265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3642__A1 (.DIODE(_1265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3633__A1 (.DIODE(_1265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3624__A1 (.DIODE(_1265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3615__A1 (.DIODE(_1265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3191__A (.DIODE(_1265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2814__A (.DIODE(_1265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3183__A1 (.DIODE(_1266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3174__A1 (.DIODE(_1266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3165__A1 (.DIODE(_1266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3116__A1 (.DIODE(_1266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3061__A1 (.DIODE(_1266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2991__A1 (.DIODE(_1266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2982__A1 (.DIODE(_1266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2964__A1 (.DIODE(_1266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2831__A1 (.DIODE(_1266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2816__A1 (.DIODE(_1266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4137__A1 (.DIODE(_1269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4089__A1 (.DIODE(_1269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4044__A1 (.DIODE(_1269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3671__A1 (.DIODE(_1269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3644__A1 (.DIODE(_1269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3635__A1 (.DIODE(_1269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3626__A1 (.DIODE(_1269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3617__A1 (.DIODE(_1269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3195__A (.DIODE(_1269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2819__A (.DIODE(_1269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3185__A1 (.DIODE(_1270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3176__A1 (.DIODE(_1270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3167__A1 (.DIODE(_1270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3118__A1 (.DIODE(_1270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3063__A1 (.DIODE(_1270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2993__A1 (.DIODE(_1270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2984__A1 (.DIODE(_1270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2966__A1 (.DIODE(_1270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2833__A1 (.DIODE(_1270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2820__A1 (.DIODE(_1270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4139__A1 (.DIODE(_1272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4091__A1 (.DIODE(_1272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4046__A1 (.DIODE(_1272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3673__A1 (.DIODE(_1272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3646__A1 (.DIODE(_1272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3637__A1 (.DIODE(_1272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3628__A1 (.DIODE(_1272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3619__A1 (.DIODE(_1272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3198__A (.DIODE(_1272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2823__A (.DIODE(_1272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3187__A1 (.DIODE(_1273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3178__A1 (.DIODE(_1273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3169__A1 (.DIODE(_1273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3120__A1 (.DIODE(_1273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3065__A1 (.DIODE(_1273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2995__A1 (.DIODE(_1273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2986__A1 (.DIODE(_1273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2968__A1 (.DIODE(_1273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2835__A1 (.DIODE(_1273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2824__A1 (.DIODE(_1273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4141__A1 (.DIODE(_1275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4093__A1 (.DIODE(_1275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4048__A1 (.DIODE(_1275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3675__A1 (.DIODE(_1275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3648__A1 (.DIODE(_1275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3639__A1 (.DIODE(_1275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3630__A1 (.DIODE(_1275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3621__A1 (.DIODE(_1275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3201__A (.DIODE(_1275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2827__A (.DIODE(_1275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3189__A1 (.DIODE(_1276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3180__A1 (.DIODE(_1276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3171__A1 (.DIODE(_1276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3122__A1 (.DIODE(_1276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3067__A1 (.DIODE(_1276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2997__A1 (.DIODE(_1276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2988__A1 (.DIODE(_1276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2970__A1 (.DIODE(_1276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2837__A1 (.DIODE(_1276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2828__A1 (.DIODE(_1276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3696__B (.DIODE(_1293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3596__B (.DIODE(_1293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3430__B (.DIODE(_1293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3372__B (.DIODE(_1293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3242__A (.DIODE(_1293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3142__B (.DIODE(_1293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3087__B (.DIODE(_1293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2858__B (.DIODE(_1293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4077__B (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3659__B (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3560__B (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3381__B (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3206__A (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2936__B (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2896__B (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2868__B (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4032__B (.DIODE(_1305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3717__B (.DIODE(_1305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3538__B (.DIODE(_1305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3363__B (.DIODE(_1305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3260__A (.DIODE(_1305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3233__B (.DIODE(_1305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2915__B (.DIODE(_1305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2878__B (.DIODE(_1305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3028__A0 (.DIODE(_1326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3018__A0 (.DIODE(_1326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3009__A0 (.DIODE(_1326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3000__A0 (.DIODE(_1326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2973__A0 (.DIODE(_1326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2955__A0 (.DIODE(_1326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2946__A0 (.DIODE(_1326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2937__A0 (.DIODE(_1326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2928__A0 (.DIODE(_1326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2916__A0 (.DIODE(_1326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3030__A0 (.DIODE(_1329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3020__A0 (.DIODE(_1329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3011__A0 (.DIODE(_1329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3002__A0 (.DIODE(_1329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2975__A0 (.DIODE(_1329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2957__A0 (.DIODE(_1329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2948__A0 (.DIODE(_1329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2939__A0 (.DIODE(_1329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2930__A0 (.DIODE(_1329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2919__A0 (.DIODE(_1329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3032__A0 (.DIODE(_1331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3022__A0 (.DIODE(_1331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3013__A0 (.DIODE(_1331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3004__A0 (.DIODE(_1331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2977__A0 (.DIODE(_1331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2959__A0 (.DIODE(_1331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2950__A0 (.DIODE(_1331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2941__A0 (.DIODE(_1331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2932__A0 (.DIODE(_1331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2922__A0 (.DIODE(_1331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3034__A0 (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3024__A0 (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3015__A0 (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3006__A0 (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2979__A0 (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2961__A0 (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2952__A0 (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2943__A0 (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2934__A0 (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2925__A0 (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3006__S (.DIODE(_1375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3004__S (.DIODE(_1375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3002__S (.DIODE(_1375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3000__S (.DIODE(_1375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3034__S (.DIODE(_1391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3032__S (.DIODE(_1391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3030__S (.DIODE(_1391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3028__S (.DIODE(_1391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3143__A0 (.DIODE(_1396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3134__A0 (.DIODE(_1396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3125__A0 (.DIODE(_1396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3106__A0 (.DIODE(_1396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3097__A0 (.DIODE(_1396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3088__A0 (.DIODE(_1396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3079__A0 (.DIODE(_1396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3070__A0 (.DIODE(_1396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3052__A0 (.DIODE(_1396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3039__A0 (.DIODE(_1396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3048__S (.DIODE(_1398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3045__S (.DIODE(_1398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3042__S (.DIODE(_1398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3039__S (.DIODE(_1398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3145__A0 (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3136__A0 (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3127__A0 (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3108__A0 (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3099__A0 (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3090__A0 (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3081__A0 (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3072__A0 (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3054__A0 (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3042__A0 (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3147__A0 (.DIODE(_1402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3138__A0 (.DIODE(_1402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3129__A0 (.DIODE(_1402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3110__A0 (.DIODE(_1402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3101__A0 (.DIODE(_1402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3092__A0 (.DIODE(_1402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3083__A0 (.DIODE(_1402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3074__A0 (.DIODE(_1402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3056__A0 (.DIODE(_1402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3045__A0 (.DIODE(_1402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3149__A0 (.DIODE(_1404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3140__A0 (.DIODE(_1404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3131__A0 (.DIODE(_1404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3112__A0 (.DIODE(_1404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3103__A0 (.DIODE(_1404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3094__A0 (.DIODE(_1404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3085__A0 (.DIODE(_1404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3076__A0 (.DIODE(_1404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3058__A0 (.DIODE(_1404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3048__A0 (.DIODE(_1404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3058__S (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3056__S (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3054__S (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3052__S (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4032__A (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3224__A (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3192__A (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3182__B (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3173__A (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3164__B (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3152__A (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3142__A (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3124__A (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3115__A (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3140__S (.DIODE(_1453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3138__S (.DIODE(_1453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3136__S (.DIODE(_1453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3134__S (.DIODE(_1453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3297__A0 (.DIODE(_1463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3270__A0 (.DIODE(_1463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3261__A0 (.DIODE(_1463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3252__A0 (.DIODE(_1463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3243__A0 (.DIODE(_1463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3234__A0 (.DIODE(_1463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3225__A0 (.DIODE(_1463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3216__A0 (.DIODE(_1463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3207__A0 (.DIODE(_1463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3153__A0 (.DIODE(_1463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3299__A0 (.DIODE(_1466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3272__A0 (.DIODE(_1466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3263__A0 (.DIODE(_1466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3254__A0 (.DIODE(_1466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3245__A0 (.DIODE(_1466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3236__A0 (.DIODE(_1466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3227__A0 (.DIODE(_1466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3218__A0 (.DIODE(_1466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3209__A0 (.DIODE(_1466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3156__A0 (.DIODE(_1466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3301__A0 (.DIODE(_1468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3274__A0 (.DIODE(_1468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3265__A0 (.DIODE(_1468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3256__A0 (.DIODE(_1468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3247__A0 (.DIODE(_1468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3238__A0 (.DIODE(_1468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3229__A0 (.DIODE(_1468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3220__A0 (.DIODE(_1468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3211__A0 (.DIODE(_1468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3159__A0 (.DIODE(_1468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3303__A0 (.DIODE(_1470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3276__A0 (.DIODE(_1470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3267__A0 (.DIODE(_1470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3258__A0 (.DIODE(_1470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3249__A0 (.DIODE(_1470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3240__A0 (.DIODE(_1470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3231__A0 (.DIODE(_1470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3222__A0 (.DIODE(_1470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3213__A0 (.DIODE(_1470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3162__A0 (.DIODE(_1470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3570__A1 (.DIODE(_1487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3476__A1 (.DIODE(_1487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3467__A1 (.DIODE(_1487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3458__A1 (.DIODE(_1487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3449__A1 (.DIODE(_1487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3355__A1 (.DIODE(_1487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3346__A1 (.DIODE(_1487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3288__A1 (.DIODE(_1487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3279__A1 (.DIODE(_1487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3193__A1 (.DIODE(_1487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3572__A1 (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3478__A1 (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3469__A1 (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3460__A1 (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3451__A1 (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3357__A1 (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3348__A1 (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3290__A1 (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3281__A1 (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3196__A1 (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3574__A1 (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3480__A1 (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3471__A1 (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3462__A1 (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3453__A1 (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3359__A1 (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3350__A1 (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3292__A1 (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3283__A1 (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3199__A1 (.DIODE(_1492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3576__A1 (.DIODE(_1494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3482__A1 (.DIODE(_1494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3473__A1 (.DIODE(_1494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3464__A1 (.DIODE(_1494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3455__A1 (.DIODE(_1494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3361__A1 (.DIODE(_1494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3352__A1 (.DIODE(_1494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3294__A1 (.DIODE(_1494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3285__A1 (.DIODE(_1494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3202__A1 (.DIODE(_1494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3399__B (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3390__B (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3336__B (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3327__B (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3318__B (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3306__B (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3205__A (.DIODE(_1496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4041__B (.DIODE(_1497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3354__B (.DIODE(_1497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3345__B (.DIODE(_1497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3287__B (.DIODE(_1497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3278__B (.DIODE(_1497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3269__B (.DIODE(_1497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3260__B (.DIODE(_1497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3251__B (.DIODE(_1497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3242__B (.DIODE(_1497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3206__B (.DIODE(_1497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3240__S (.DIODE(_1513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3238__S (.DIODE(_1513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3236__S (.DIODE(_1513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3234__S (.DIODE(_1513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3409__A0 (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3400__A0 (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3391__A0 (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3382__A0 (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3373__A0 (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3364__A0 (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3337__A0 (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3328__A0 (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3319__A0 (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3307__A0 (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3411__A0 (.DIODE(_1556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3402__A0 (.DIODE(_1556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3393__A0 (.DIODE(_1556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3384__A0 (.DIODE(_1556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3375__A0 (.DIODE(_1556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3366__A0 (.DIODE(_1556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3339__A0 (.DIODE(_1556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3330__A0 (.DIODE(_1556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3321__A0 (.DIODE(_1556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3310__A0 (.DIODE(_1556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3413__A0 (.DIODE(_1558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3404__A0 (.DIODE(_1558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3395__A0 (.DIODE(_1558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3386__A0 (.DIODE(_1558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3377__A0 (.DIODE(_1558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3368__A0 (.DIODE(_1558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3341__A0 (.DIODE(_1558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3332__A0 (.DIODE(_1558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3323__A0 (.DIODE(_1558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3313__A0 (.DIODE(_1558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3415__A0 (.DIODE(_1560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3406__A0 (.DIODE(_1560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3397__A0 (.DIODE(_1560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3388__A0 (.DIODE(_1560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3379__A0 (.DIODE(_1560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3370__A0 (.DIODE(_1560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3343__A0 (.DIODE(_1560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3334__A0 (.DIODE(_1560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3325__A0 (.DIODE(_1560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3316__A0 (.DIODE(_1560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3539__A0 (.DIODE(_1617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3530__A0 (.DIODE(_1617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3521__A0 (.DIODE(_1617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3512__A0 (.DIODE(_1617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3503__A0 (.DIODE(_1617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3494__A0 (.DIODE(_1617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3485__A0 (.DIODE(_1617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3440__A0 (.DIODE(_1617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3431__A0 (.DIODE(_1617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3419__A0 (.DIODE(_1617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3541__A0 (.DIODE(_1620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3532__A0 (.DIODE(_1620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3523__A0 (.DIODE(_1620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3514__A0 (.DIODE(_1620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3505__A0 (.DIODE(_1620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3496__A0 (.DIODE(_1620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3487__A0 (.DIODE(_1620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3442__A0 (.DIODE(_1620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3433__A0 (.DIODE(_1620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3422__A0 (.DIODE(_1620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3543__A0 (.DIODE(_1622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3534__A0 (.DIODE(_1622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3525__A0 (.DIODE(_1622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3516__A0 (.DIODE(_1622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3507__A0 (.DIODE(_1622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3498__A0 (.DIODE(_1622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3489__A0 (.DIODE(_1622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3444__A0 (.DIODE(_1622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3435__A0 (.DIODE(_1622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3425__A0 (.DIODE(_1622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3545__A0 (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3536__A0 (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3527__A0 (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3518__A0 (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3509__A0 (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3500__A0 (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3491__A0 (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3446__A0 (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3437__A0 (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3428__A0 (.DIODE(_1624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3687__A0 (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3678__A0 (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3660__A0 (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3651__A0 (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3606__A0 (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3597__A0 (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3588__A0 (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3579__A0 (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3561__A0 (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3549__A0 (.DIODE(_1691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3689__A0 (.DIODE(_1694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3680__A0 (.DIODE(_1694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3662__A0 (.DIODE(_1694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3653__A0 (.DIODE(_1694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3608__A0 (.DIODE(_1694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3599__A0 (.DIODE(_1694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3590__A0 (.DIODE(_1694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3581__A0 (.DIODE(_1694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3563__A0 (.DIODE(_1694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3552__A0 (.DIODE(_1694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3691__A0 (.DIODE(_1696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3682__A0 (.DIODE(_1696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3664__A0 (.DIODE(_1696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3655__A0 (.DIODE(_1696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3610__A0 (.DIODE(_1696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3601__A0 (.DIODE(_1696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3592__A0 (.DIODE(_1696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3583__A0 (.DIODE(_1696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3565__A0 (.DIODE(_1696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3555__A0 (.DIODE(_1696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3693__A0 (.DIODE(_1698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3684__A0 (.DIODE(_1698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3666__A0 (.DIODE(_1698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3657__A0 (.DIODE(_1698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3612__A0 (.DIODE(_1698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3603__A0 (.DIODE(_1698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3594__A0 (.DIODE(_1698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3585__A0 (.DIODE(_1698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3567__A0 (.DIODE(_1698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3558__A0 (.DIODE(_1698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4078__A0 (.DIODE(_1775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4069__A0 (.DIODE(_1775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4060__A0 (.DIODE(_1775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4051__A0 (.DIODE(_1775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4033__A0 (.DIODE(_1775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4024__A0 (.DIODE(_1775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3727__A0 (.DIODE(_1775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3718__A0 (.DIODE(_1775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3709__A0 (.DIODE(_1775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3697__A0 (.DIODE(_1775_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4080__A0 (.DIODE(_1778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4071__A0 (.DIODE(_1778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4062__A0 (.DIODE(_1778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4053__A0 (.DIODE(_1778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4035__A0 (.DIODE(_1778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4026__A0 (.DIODE(_1778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3729__A0 (.DIODE(_1778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3720__A0 (.DIODE(_1778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3711__A0 (.DIODE(_1778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3700__A0 (.DIODE(_1778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4082__A0 (.DIODE(_1780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4073__A0 (.DIODE(_1780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4064__A0 (.DIODE(_1780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4055__A0 (.DIODE(_1780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4037__A0 (.DIODE(_1780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4028__A0 (.DIODE(_1780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3731__A0 (.DIODE(_1780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3722__A0 (.DIODE(_1780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3713__A0 (.DIODE(_1780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3703__A0 (.DIODE(_1780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4084__A0 (.DIODE(_1782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4075__A0 (.DIODE(_1782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4066__A0 (.DIODE(_1782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4057__A0 (.DIODE(_1782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4039__A0 (.DIODE(_1782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4030__A0 (.DIODE(_1782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3733__A0 (.DIODE(_1782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3724__A0 (.DIODE(_1782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3715__A0 (.DIODE(_1782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3706__A0 (.DIODE(_1782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3924__B1 (.DIODE(_1807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3883__A (.DIODE(_1807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3879__A (.DIODE(_1807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3871__C1 (.DIODE(_1807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3784__A (.DIODE(_1807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3763__A (.DIODE(_1807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3759__A (.DIODE(_1807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3755__B1 (.DIODE(_1807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3754__A (.DIODE(_1807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3751__B (.DIODE(_1807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3860__C1 (.DIODE(_1826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3857__C1 (.DIODE(_1826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3854__C1 (.DIODE(_1826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3851__C1 (.DIODE(_1826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3845__C1 (.DIODE(_1826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3842__C1 (.DIODE(_1826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3839__C1 (.DIODE(_1826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3791__C1 (.DIODE(_1826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3788__C1 (.DIODE(_1826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3776__C1 (.DIODE(_1826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4013__D_N (.DIODE(_1830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3994__B (.DIODE(_1830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3969__A2 (.DIODE(_1830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3968__A (.DIODE(_1830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3952__A1 (.DIODE(_1830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3949__D (.DIODE(_1830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3930__A1 (.DIODE(_1830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3878__A0 (.DIODE(_1830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3847__B (.DIODE(_1830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3781__B2 (.DIODE(_1830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3836__C1 (.DIODE(_1844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3830__C1 (.DIODE(_1844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3828__C1 (.DIODE(_1844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3826__C1 (.DIODE(_1844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3823__A (.DIODE(_1844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3818__A (.DIODE(_1844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3813__A (.DIODE(_1844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3809__C1 (.DIODE(_1844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3804__A (.DIODE(_1844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3800__C1 (.DIODE(_1844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3904__S (.DIODE(_1913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3902__S (.DIODE(_1913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3900__S (.DIODE(_1913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3898__S (.DIODE(_1913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3896__S (.DIODE(_1913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3894__S (.DIODE(_1913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3993__A2 (.DIODE(_1968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3992__A (.DIODE(_1968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3988__A2 (.DIODE(_1968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3987__A (.DIODE(_1968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3981__A2 (.DIODE(_1968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3980__A (.DIODE(_1968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3974__A2 (.DIODE(_1968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3973__A (.DIODE(_1968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4132__S (.DIODE(_2058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4130__S (.DIODE(_2058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4128__S (.DIODE(_2058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4126__S (.DIODE(_2058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4124__S (.DIODE(_2058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4122__S (.DIODE(_2058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4120__S (.DIODE(_2058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4118__S (.DIODE(_2058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4116__S (.DIODE(_2058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4114__S (.DIODE(_2058_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(io_in[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(io_in[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(io_in[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(io_in[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(oram_value[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(oram_value[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(oram_value[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(oram_value[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(oram_value[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(oram_value[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(oram_value[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(oram_value[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(oram_value[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(oram_value[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(oram_value[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA__4747__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4750__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4681__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4671__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4707__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4719__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4706__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4613__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4670__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4669__CLK (.DIODE(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__3234__A1 (.DIODE(\tms1x00.RAM[2][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2233__A2 (.DIODE(\tms1x00.RAM[2][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3236__A1 (.DIODE(\tms1x00.RAM[2][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2350__A2 (.DIODE(\tms1x00.RAM[2][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3238__A1 (.DIODE(\tms1x00.RAM[2][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2453__A2 (.DIODE(\tms1x00.RAM[2][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3297__A1 (.DIODE(\tms1x00.RAM[3][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2233__A3 (.DIODE(\tms1x00.RAM[3][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3299__A1 (.DIODE(\tms1x00.RAM[3][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2350__A3 (.DIODE(\tms1x00.RAM[3][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3301__A1 (.DIODE(\tms1x00.RAM[3][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2453__A3 (.DIODE(\tms1x00.RAM[3][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3820__C (.DIODE(\tms1x00.Y[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3815__A_N (.DIODE(\tms1x00.Y[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3810__B (.DIODE(\tms1x00.Y[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3807__B (.DIODE(\tms1x00.Y[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3801__C (.DIODE(\tms1x00.Y[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3793__C_N (.DIODE(\tms1x00.Y[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2074__A (.DIODE(\tms1x00.Y[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3962__B2 (.DIODE(\tms1x00.Y[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3820__A (.DIODE(\tms1x00.Y[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3815__C (.DIODE(\tms1x00.Y[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3810__C (.DIODE(\tms1x00.Y[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3807__C_N (.DIODE(\tms1x00.Y[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3801__A_N (.DIODE(\tms1x00.Y[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2087__A (.DIODE(\tms1x00.Y[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3961__A1 (.DIODE(\tms1x00.ins_in[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3950__A (.DIODE(\tms1x00.ins_in[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3928__A1 (.DIODE(\tms1x00.ins_in[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3876__C (.DIODE(\tms1x00.ins_in[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3776__A1 (.DIODE(\tms1x00.ins_in[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2282__A (.DIODE(\tms1x00.ins_in[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2122__A_N (.DIODE(\tms1x00.ins_in[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2105__A (.DIODE(\tms1x00.ins_in[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3050__B (.DIODE(\tms1x00.ram_addr_buff[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3037__A (.DIODE(\tms1x00.ram_addr_buff[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3026__D_N (.DIODE(\tms1x00.ram_addr_buff[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2762__B (.DIODE(\tms1x00.ram_addr_buff[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2749__C_N (.DIODE(\tms1x00.ram_addr_buff[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2647__A (.DIODE(\tms1x00.ram_addr_buff[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2606__A (.DIODE(\tms1x00.ram_addr_buff[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2292__B (.DIODE(\tms1x00.ram_addr_buff[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2084__A (.DIODE(\tms1x00.ram_addr_buff[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3741__A1 (.DIODE(\tms1x00.ram_addr_buff[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3050__D_N (.DIODE(\tms1x00.ram_addr_buff[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3037__C_N (.DIODE(\tms1x00.ram_addr_buff[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3026__C_N (.DIODE(\tms1x00.ram_addr_buff[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2646__A (.DIODE(\tms1x00.ram_addr_buff[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2633__B (.DIODE(\tms1x00.ram_addr_buff[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2605__C_N (.DIODE(\tms1x00.ram_addr_buff[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2294__B (.DIODE(\tms1x00.ram_addr_buff[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2092__A1 (.DIODE(\tms1x00.ram_addr_buff[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3743__A1 (.DIODE(\tms1x00.ram_addr_buff[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3204__A (.DIODE(\tms1x00.ram_addr_buff[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2760__A (.DIODE(\tms1x00.ram_addr_buff[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2688__C_N (.DIODE(\tms1x00.ram_addr_buff[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2667__A (.DIODE(\tms1x00.ram_addr_buff[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2644__A (.DIODE(\tms1x00.ram_addr_buff[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2620__C (.DIODE(\tms1x00.ram_addr_buff[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2603__C (.DIODE(\tms1x00.ram_addr_buff[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2290__A_N (.DIODE(\tms1x00.ram_addr_buff[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2094__A1 (.DIODE(\tms1x00.ram_addr_buff[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3745__A1 (.DIODE(\tms1x00.ram_addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3204__C_N (.DIODE(\tms1x00.ram_addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2760__B (.DIODE(\tms1x00.ram_addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2688__A (.DIODE(\tms1x00.ram_addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2667__B (.DIODE(\tms1x00.ram_addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2644__B (.DIODE(\tms1x00.ram_addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2620__B (.DIODE(\tms1x00.ram_addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2603__A_N (.DIODE(\tms1x00.ram_addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2290__B (.DIODE(\tms1x00.ram_addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2096__A1 (.DIODE(\tms1x00.ram_addr_buff[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3747__A1 (.DIODE(\tms1x00.ram_addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3204__B (.DIODE(\tms1x00.ram_addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2760__C (.DIODE(\tms1x00.ram_addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2688__B (.DIODE(\tms1x00.ram_addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2667__C (.DIODE(\tms1x00.ram_addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2644__C_N (.DIODE(\tms1x00.ram_addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2620__A_N (.DIODE(\tms1x00.ram_addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2603__B (.DIODE(\tms1x00.ram_addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2290__C (.DIODE(\tms1x00.ram_addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2098__A1 (.DIODE(\tms1x00.ram_addr_buff[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_wb_clk_i_A (.DIODE(wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(wb_rst_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(wbs_adr_i[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(wbs_adr_i[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(wbs_adr_i[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(wbs_adr_i[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(wbs_adr_i[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(wbs_adr_i[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(wbs_adr_i[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(wbs_adr_i[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(wbs_adr_i[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(wbs_adr_i[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(wbs_we_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__3757__A0 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__4813__A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__4013__B (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__3943__C (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__3749__A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__2283__B (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__2124__B (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__2076__A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__4814__A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__4815__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__4816__A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__4817__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__4818__A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__4819__A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__4820__A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__4821__A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__4822__A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__2101__A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_output33_A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__3951__A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__3944__A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__3753__B (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__3752__A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__3751__A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__2123__B (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__2108__B (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__2077__A_N (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_output34_A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__3943__B (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__3765__A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__3753__A_N (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__3752__B (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__2123__C_N (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__2108__C (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__2078__A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_output35_A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__3943__A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__3753__C (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__2124__A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__2108__A_N (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__2077__B (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_output36_A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__2118__B1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_output37_A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__3794__B1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_output40_A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__3808__B1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_output44_A (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__3825__B1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_output45_A (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__3827__B1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_output46_A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__3829__B1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_output47_A (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__3831__B1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_output48_A (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__3835__B1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_output49_A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__3838__B1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_output50_A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__3841__B1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_output51_A (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__3844__B1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_output61_A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_output62_A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_output63_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_output64_A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_output65_A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_output66_A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_output67_A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_output68_A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_output69_A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_output71_A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__4545__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4539__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4541__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4536__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4718__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4532__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4540__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4726__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4177__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4610__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4587__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4589__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4614__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4615__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4609__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4611__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4607__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4727__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4709__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4729__CLK (.DIODE(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4531__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4533__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4538__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4534__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4592__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4399__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4527__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4591__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4555__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4593__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4557__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4216__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4558__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4606__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4556__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4594__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4179__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4176__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4590__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4546__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4544__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4542__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4543__CLK (.DIODE(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4521__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4522__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4520__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4513__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4396__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4516__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4524__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4488__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4490__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4411__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4419__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4485__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4489__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4514__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4483__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4487__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4486__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4464__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4463__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4528__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4518__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4525__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4434__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4526__CLK (.DIODE(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4666__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4661__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4678__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4393__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4398__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4431__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4517__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4515__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4667__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4433__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4662__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4511__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4365__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4519__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4523__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4395__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4535__CLK (.DIODE(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4633__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4636__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4635__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4692__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4683__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4691__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4418__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4693__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4415__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4417__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4421__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4413__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4409__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4410__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4408__CLK (.DIODE(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4690__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4659__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4688__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4660__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4143__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4420__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4401__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4621__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4711__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4438__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4441__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4402__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4437__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4385__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4387__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4414__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4623__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4422__CLK (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4459__CLK (.DIODE(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4470__CLK (.DIODE(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4345__CLK (.DIODE(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4479__CLK (.DIODE(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4482__CLK (.DIODE(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4344__CLK (.DIODE(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4347__CLK (.DIODE(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4247__CLK (.DIODE(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4246__CLK (.DIODE(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4245__CLK (.DIODE(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4244__CLK (.DIODE(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4530__CLK (.DIODE(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4491__CLK (.DIODE(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4466__CLK (.DIODE(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4468__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4175__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4469__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4172__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4330__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4467__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4404__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4407__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4405__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4447__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4302__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4259__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4341__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4331__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4342__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4733__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4730__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4508__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4481__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4732__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4480__CLK (.DIODE(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4269__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4258__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4261__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4263__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4271__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4257__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4275__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4280__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4283__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4314__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4256__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4304__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4168__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4170__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4301__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4300__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4305__CLK (.DIODE(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4333__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4332__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4323__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4336__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4337__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4339__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4239__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4243__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4338__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4334__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4306__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4169__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4171__CLK (.DIODE(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4359__CLK (.DIODE(clknet_leaf_25_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4346__CLK (.DIODE(clknet_leaf_25_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4507__CLK (.DIODE(clknet_leaf_25_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4355__CLK (.DIODE(clknet_leaf_25_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4510__CLK (.DIODE(clknet_leaf_25_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4350__CLK (.DIODE(clknet_leaf_25_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4167__CLK (.DIODE(clknet_leaf_25_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4164__CLK (.DIODE(clknet_leaf_25_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4351__CLK (.DIODE(clknet_leaf_25_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4595__CLK (.DIODE(clknet_leaf_25_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4349__CLK (.DIODE(clknet_leaf_25_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4363__CLK (.DIODE(clknet_leaf_25_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4353__CLK (.DIODE(clknet_leaf_25_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4352__CLK (.DIODE(clknet_leaf_25_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4362__CLK (.DIODE(clknet_leaf_25_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4354__CLK (.DIODE(clknet_leaf_25_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4509__CLK (.DIODE(clknet_leaf_25_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4358__CLK (.DIODE(clknet_leaf_25_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4329__CLK (.DIODE(clknet_leaf_25_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4731__CLK (.DIODE(clknet_leaf_25_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4328__CLK (.DIODE(clknet_leaf_25_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4562__CLK (.DIODE(clknet_leaf_26_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4596__CLK (.DIODE(clknet_leaf_26_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4597__CLK (.DIODE(clknet_leaf_26_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4166__CLK (.DIODE(clknet_leaf_26_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4165__CLK (.DIODE(clknet_leaf_26_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4566__CLK (.DIODE(clknet_leaf_26_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4598__CLK (.DIODE(clknet_leaf_26_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4219__CLK (.DIODE(clknet_leaf_26_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4217__CLK (.DIODE(clknet_leaf_26_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4218__CLK (.DIODE(clknet_leaf_26_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4163__CLK (.DIODE(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4559__CLK (.DIODE(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4161__CLK (.DIODE(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4375__CLK (.DIODE(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4162__CLK (.DIODE(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4383__CLK (.DIODE(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4374__CLK (.DIODE(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4506__CLK (.DIODE(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4502__CLK (.DIODE(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4500__CLK (.DIODE(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4501__CLK (.DIODE(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4499__CLK (.DIODE(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4324__CLK (.DIODE(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4495__CLK (.DIODE(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4553__CLK (.DIODE(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4498__CLK (.DIODE(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4496__CLK (.DIODE(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4549__CLK (.DIODE(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4554__CLK (.DIODE(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4560__CLK (.DIODE(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4561__CLK (.DIODE(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4550__CLK (.DIODE(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4547__CLK (.DIODE(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4551__CLK (.DIODE(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4208__CLK (.DIODE(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4210__CLK (.DIODE(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4226__CLK (.DIODE(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4293__CLK (.DIODE(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4224__CLK (.DIODE(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4297__CLK (.DIODE(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4292__CLK (.DIODE(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4294__CLK (.DIODE(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4298__CLK (.DIODE(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4296__CLK (.DIODE(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4209__CLK (.DIODE(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4222__CLK (.DIODE(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4220__CLK (.DIODE(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4151__CLK (.DIODE(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4154__CLK (.DIODE(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4153__CLK (.DIODE(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4223__CLK (.DIODE(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4221__CLK (.DIODE(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4737__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4738__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4206__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4198__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4205__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4202__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4201__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4200__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4196__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4197__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4287__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4203__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4199__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4211__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4149__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4150__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4148__CLK (.DIODE(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4741__CLK (.DIODE(clknet_leaf_33_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4582__CLK (.DIODE(clknet_leaf_33_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4754__CLK (.DIODE(clknet_leaf_33_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4753__CLK (.DIODE(clknet_leaf_33_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4752__CLK (.DIODE(clknet_leaf_33_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4213__CLK (.DIODE(clknet_leaf_33_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4214__CLK (.DIODE(clknet_leaf_33_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4552__CLK (.DIODE(clknet_leaf_33_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4548__CLK (.DIODE(clknet_leaf_33_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4755__CLK (.DIODE(clknet_leaf_33_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4284__CLK (.DIODE(clknet_leaf_33_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4497__CLK (.DIODE(clknet_leaf_33_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4155__CLK (.DIODE(clknet_leaf_33_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4285__CLK (.DIODE(clknet_leaf_33_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4152__CLK (.DIODE(clknet_leaf_33_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4574__CLK (.DIODE(clknet_leaf_34_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4570__CLK (.DIODE(clknet_leaf_34_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4577__CLK (.DIODE(clknet_leaf_34_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4581__CLK (.DIODE(clknet_leaf_34_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4579__CLK (.DIODE(clknet_leaf_34_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4600__CLK (.DIODE(clknet_leaf_34_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4575__CLK (.DIODE(clknet_leaf_34_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4605__CLK (.DIODE(clknet_leaf_34_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4604__CLK (.DIODE(clknet_leaf_34_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4567__CLK (.DIODE(clknet_leaf_34_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4178__CLK (.DIODE(clknet_leaf_34_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4599__CLK (.DIODE(clknet_leaf_34_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4212__CLK (.DIODE(clknet_leaf_34_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4603__CLK (.DIODE(clknet_leaf_34_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4565__CLK (.DIODE(clknet_leaf_34_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4602__CLK (.DIODE(clknet_leaf_34_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4563__CLK (.DIODE(clknet_leaf_34_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4583__CLK (.DIODE(clknet_leaf_34_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4564__CLK (.DIODE(clknet_leaf_34_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4584__CLK (.DIODE(clknet_leaf_34_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4585__CLK (.DIODE(clknet_leaf_34_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4586__CLK (.DIODE(clknet_leaf_34_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4601__CLK (.DIODE(clknet_leaf_34_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4578__CLK (.DIODE(clknet_leaf_34_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4215__CLK (.DIODE(clknet_leaf_34_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4734__CLK (.DIODE(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4716__CLK (.DIODE(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4714__CLK (.DIODE(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4703__CLK (.DIODE(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4702__CLK (.DIODE(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4715__CLK (.DIODE(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4705__CLK (.DIODE(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4616__CLK (.DIODE(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4612__CLK (.DIODE(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4608__CLK (.DIODE(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4617__CLK (.DIODE(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4568__CLK (.DIODE(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4569__CLK (.DIODE(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4588__CLK (.DIODE(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4618__CLK (.DIODE(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4571__CLK (.DIODE(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4573__CLK (.DIODE(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4572__CLK (.DIODE(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4580__CLK (.DIODE(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4576__CLK (.DIODE(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_37_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__4704__CLK (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_639 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_534 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_690 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_826 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_639 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_760 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_796 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_796 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_534 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_814 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_774 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_450 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_618 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_667 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_663 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_676 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_796 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_693 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_663 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_695 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_704 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_676 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_555 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_690 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_807 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_826 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_555 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_560 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_841 ();
 assign io_oeb[0] = net119;
 assign io_oeb[10] = net77;
 assign io_oeb[11] = net78;
 assign io_oeb[12] = net79;
 assign io_oeb[13] = net80;
 assign io_oeb[14] = net81;
 assign io_oeb[15] = net82;
 assign io_oeb[16] = net83;
 assign io_oeb[17] = net84;
 assign io_oeb[18] = net85;
 assign io_oeb[19] = net86;
 assign io_oeb[1] = net120;
 assign io_oeb[20] = net87;
 assign io_oeb[21] = net88;
 assign io_oeb[22] = net89;
 assign io_oeb[23] = net90;
 assign io_oeb[24] = net91;
 assign io_oeb[25] = net92;
 assign io_oeb[26] = net93;
 assign io_oeb[27] = net94;
 assign io_oeb[28] = net95;
 assign io_oeb[29] = net96;
 assign io_oeb[2] = net121;
 assign io_oeb[30] = net97;
 assign io_oeb[31] = net98;
 assign io_oeb[32] = net99;
 assign io_oeb[33] = net100;
 assign io_oeb[34] = net101;
 assign io_oeb[35] = net102;
 assign io_oeb[36] = net103;
 assign io_oeb[37] = net124;
 assign io_oeb[3] = net122;
 assign io_oeb[4] = net123;
 assign io_oeb[5] = net72;
 assign io_oeb[6] = net73;
 assign io_oeb[7] = net74;
 assign io_oeb[8] = net75;
 assign io_oeb[9] = net76;
 assign io_out[0] = net104;
 assign io_out[1] = net105;
 assign io_out[2] = net106;
 assign io_out[34] = net114;
 assign io_out[35] = net115;
 assign io_out[36] = net116;
 assign io_out[37] = net117;
 assign io_out[3] = net107;
 assign io_out[4] = net108;
 assign io_out[5] = net109;
 assign io_out[6] = net110;
 assign io_out[7] = net111;
 assign io_out[8] = net112;
 assign io_out[9] = net113;
 assign oram_addr[8] = net118;
 assign ram_wmask[0] = net125;
 assign ram_wmask[1] = net126;
 assign ram_wmask[2] = net127;
 assign ram_wmask[3] = net128;
endmodule

