magic
tech sky130B
magscale 1 2
timestamp 1672430794
<< obsli1 >>
rect 1104 2159 198812 197489
<< obsm1 >>
rect 1104 212 199074 197520
<< metal2 >>
rect 1214 199200 1270 200000
rect 2962 199200 3018 200000
rect 4710 199200 4766 200000
rect 6458 199200 6514 200000
rect 8206 199200 8262 200000
rect 9954 199200 10010 200000
rect 11702 199200 11758 200000
rect 13450 199200 13506 200000
rect 15198 199200 15254 200000
rect 16946 199200 17002 200000
rect 18694 199200 18750 200000
rect 20442 199200 20498 200000
rect 22190 199200 22246 200000
rect 23938 199200 23994 200000
rect 25686 199200 25742 200000
rect 27434 199200 27490 200000
rect 29182 199200 29238 200000
rect 30930 199200 30986 200000
rect 32678 199200 32734 200000
rect 34426 199200 34482 200000
rect 36174 199200 36230 200000
rect 37922 199200 37978 200000
rect 39670 199200 39726 200000
rect 41418 199200 41474 200000
rect 43166 199200 43222 200000
rect 44914 199200 44970 200000
rect 46662 199200 46718 200000
rect 48410 199200 48466 200000
rect 50158 199200 50214 200000
rect 51906 199200 51962 200000
rect 53654 199200 53710 200000
rect 55402 199200 55458 200000
rect 57150 199200 57206 200000
rect 58898 199200 58954 200000
rect 60646 199200 60702 200000
rect 62394 199200 62450 200000
rect 64142 199200 64198 200000
rect 65890 199200 65946 200000
rect 67638 199200 67694 200000
rect 69386 199200 69442 200000
rect 71134 199200 71190 200000
rect 72882 199200 72938 200000
rect 74630 199200 74686 200000
rect 76378 199200 76434 200000
rect 78126 199200 78182 200000
rect 79874 199200 79930 200000
rect 81622 199200 81678 200000
rect 83370 199200 83426 200000
rect 85118 199200 85174 200000
rect 86866 199200 86922 200000
rect 88614 199200 88670 200000
rect 90362 199200 90418 200000
rect 92110 199200 92166 200000
rect 93858 199200 93914 200000
rect 95606 199200 95662 200000
rect 97354 199200 97410 200000
rect 99102 199200 99158 200000
rect 100850 199200 100906 200000
rect 102598 199200 102654 200000
rect 104346 199200 104402 200000
rect 106094 199200 106150 200000
rect 107842 199200 107898 200000
rect 109590 199200 109646 200000
rect 111338 199200 111394 200000
rect 113086 199200 113142 200000
rect 114834 199200 114890 200000
rect 116582 199200 116638 200000
rect 118330 199200 118386 200000
rect 120078 199200 120134 200000
rect 121826 199200 121882 200000
rect 123574 199200 123630 200000
rect 125322 199200 125378 200000
rect 127070 199200 127126 200000
rect 128818 199200 128874 200000
rect 130566 199200 130622 200000
rect 132314 199200 132370 200000
rect 134062 199200 134118 200000
rect 135810 199200 135866 200000
rect 137558 199200 137614 200000
rect 139306 199200 139362 200000
rect 141054 199200 141110 200000
rect 142802 199200 142858 200000
rect 144550 199200 144606 200000
rect 146298 199200 146354 200000
rect 148046 199200 148102 200000
rect 149794 199200 149850 200000
rect 151542 199200 151598 200000
rect 153290 199200 153346 200000
rect 155038 199200 155094 200000
rect 156786 199200 156842 200000
rect 158534 199200 158590 200000
rect 160282 199200 160338 200000
rect 162030 199200 162086 200000
rect 163778 199200 163834 200000
rect 165526 199200 165582 200000
rect 167274 199200 167330 200000
rect 169022 199200 169078 200000
rect 170770 199200 170826 200000
rect 172518 199200 172574 200000
rect 174266 199200 174322 200000
rect 176014 199200 176070 200000
rect 177762 199200 177818 200000
rect 179510 199200 179566 200000
rect 181258 199200 181314 200000
rect 183006 199200 183062 200000
rect 184754 199200 184810 200000
rect 186502 199200 186558 200000
rect 188250 199200 188306 200000
rect 189998 199200 190054 200000
rect 191746 199200 191802 200000
rect 193494 199200 193550 200000
rect 195242 199200 195298 200000
rect 196990 199200 197046 200000
rect 198738 199200 198794 200000
rect 2410 0 2466 800
rect 4342 0 4398 800
rect 6274 0 6330 800
rect 8206 0 8262 800
rect 10138 0 10194 800
rect 12070 0 12126 800
rect 14002 0 14058 800
rect 15934 0 15990 800
rect 17866 0 17922 800
rect 19798 0 19854 800
rect 21730 0 21786 800
rect 23662 0 23718 800
rect 25594 0 25650 800
rect 27526 0 27582 800
rect 29458 0 29514 800
rect 31390 0 31446 800
rect 33322 0 33378 800
rect 35254 0 35310 800
rect 37186 0 37242 800
rect 39118 0 39174 800
rect 41050 0 41106 800
rect 42982 0 43038 800
rect 44914 0 44970 800
rect 46846 0 46902 800
rect 48778 0 48834 800
rect 50710 0 50766 800
rect 52642 0 52698 800
rect 54574 0 54630 800
rect 56506 0 56562 800
rect 58438 0 58494 800
rect 60370 0 60426 800
rect 62302 0 62358 800
rect 64234 0 64290 800
rect 66166 0 66222 800
rect 68098 0 68154 800
rect 70030 0 70086 800
rect 71962 0 72018 800
rect 73894 0 73950 800
rect 75826 0 75882 800
rect 77758 0 77814 800
rect 79690 0 79746 800
rect 81622 0 81678 800
rect 83554 0 83610 800
rect 85486 0 85542 800
rect 87418 0 87474 800
rect 89350 0 89406 800
rect 91282 0 91338 800
rect 93214 0 93270 800
rect 95146 0 95202 800
rect 97078 0 97134 800
rect 99010 0 99066 800
rect 100942 0 100998 800
rect 102874 0 102930 800
rect 104806 0 104862 800
rect 106738 0 106794 800
rect 108670 0 108726 800
rect 110602 0 110658 800
rect 112534 0 112590 800
rect 114466 0 114522 800
rect 116398 0 116454 800
rect 118330 0 118386 800
rect 120262 0 120318 800
rect 122194 0 122250 800
rect 124126 0 124182 800
rect 126058 0 126114 800
rect 127990 0 128046 800
rect 129922 0 129978 800
rect 131854 0 131910 800
rect 133786 0 133842 800
rect 135718 0 135774 800
rect 137650 0 137706 800
rect 139582 0 139638 800
rect 141514 0 141570 800
rect 143446 0 143502 800
rect 145378 0 145434 800
rect 147310 0 147366 800
rect 149242 0 149298 800
rect 151174 0 151230 800
rect 153106 0 153162 800
rect 155038 0 155094 800
rect 156970 0 157026 800
rect 158902 0 158958 800
rect 160834 0 160890 800
rect 162766 0 162822 800
rect 164698 0 164754 800
rect 166630 0 166686 800
rect 168562 0 168618 800
rect 170494 0 170550 800
rect 172426 0 172482 800
rect 174358 0 174414 800
rect 176290 0 176346 800
rect 178222 0 178278 800
rect 180154 0 180210 800
rect 182086 0 182142 800
rect 184018 0 184074 800
rect 185950 0 186006 800
rect 187882 0 187938 800
rect 189814 0 189870 800
rect 191746 0 191802 800
rect 193678 0 193734 800
rect 195610 0 195666 800
rect 197542 0 197598 800
<< obsm2 >>
rect 1398 199144 2906 199322
rect 3074 199144 4654 199322
rect 4822 199144 6402 199322
rect 6570 199144 8150 199322
rect 8318 199144 9898 199322
rect 10066 199144 11646 199322
rect 11814 199144 13394 199322
rect 13562 199144 15142 199322
rect 15310 199144 16890 199322
rect 17058 199144 18638 199322
rect 18806 199144 20386 199322
rect 20554 199144 22134 199322
rect 22302 199144 23882 199322
rect 24050 199144 25630 199322
rect 25798 199144 27378 199322
rect 27546 199144 29126 199322
rect 29294 199144 30874 199322
rect 31042 199144 32622 199322
rect 32790 199144 34370 199322
rect 34538 199144 36118 199322
rect 36286 199144 37866 199322
rect 38034 199144 39614 199322
rect 39782 199144 41362 199322
rect 41530 199144 43110 199322
rect 43278 199144 44858 199322
rect 45026 199144 46606 199322
rect 46774 199144 48354 199322
rect 48522 199144 50102 199322
rect 50270 199144 51850 199322
rect 52018 199144 53598 199322
rect 53766 199144 55346 199322
rect 55514 199144 57094 199322
rect 57262 199144 58842 199322
rect 59010 199144 60590 199322
rect 60758 199144 62338 199322
rect 62506 199144 64086 199322
rect 64254 199144 65834 199322
rect 66002 199144 67582 199322
rect 67750 199144 69330 199322
rect 69498 199144 71078 199322
rect 71246 199144 72826 199322
rect 72994 199144 74574 199322
rect 74742 199144 76322 199322
rect 76490 199144 78070 199322
rect 78238 199144 79818 199322
rect 79986 199144 81566 199322
rect 81734 199144 83314 199322
rect 83482 199144 85062 199322
rect 85230 199144 86810 199322
rect 86978 199144 88558 199322
rect 88726 199144 90306 199322
rect 90474 199144 92054 199322
rect 92222 199144 93802 199322
rect 93970 199144 95550 199322
rect 95718 199144 97298 199322
rect 97466 199144 99046 199322
rect 99214 199144 100794 199322
rect 100962 199144 102542 199322
rect 102710 199144 104290 199322
rect 104458 199144 106038 199322
rect 106206 199144 107786 199322
rect 107954 199144 109534 199322
rect 109702 199144 111282 199322
rect 111450 199144 113030 199322
rect 113198 199144 114778 199322
rect 114946 199144 116526 199322
rect 116694 199144 118274 199322
rect 118442 199144 120022 199322
rect 120190 199144 121770 199322
rect 121938 199144 123518 199322
rect 123686 199144 125266 199322
rect 125434 199144 127014 199322
rect 127182 199144 128762 199322
rect 128930 199144 130510 199322
rect 130678 199144 132258 199322
rect 132426 199144 134006 199322
rect 134174 199144 135754 199322
rect 135922 199144 137502 199322
rect 137670 199144 139250 199322
rect 139418 199144 140998 199322
rect 141166 199144 142746 199322
rect 142914 199144 144494 199322
rect 144662 199144 146242 199322
rect 146410 199144 147990 199322
rect 148158 199144 149738 199322
rect 149906 199144 151486 199322
rect 151654 199144 153234 199322
rect 153402 199144 154982 199322
rect 155150 199144 156730 199322
rect 156898 199144 158478 199322
rect 158646 199144 160226 199322
rect 160394 199144 161974 199322
rect 162142 199144 163722 199322
rect 163890 199144 165470 199322
rect 165638 199144 167218 199322
rect 167386 199144 168966 199322
rect 169134 199144 170714 199322
rect 170882 199144 172462 199322
rect 172630 199144 174210 199322
rect 174378 199144 175958 199322
rect 176126 199144 177706 199322
rect 177874 199144 179454 199322
rect 179622 199144 181202 199322
rect 181370 199144 182950 199322
rect 183118 199144 184698 199322
rect 184866 199144 186446 199322
rect 186614 199144 188194 199322
rect 188362 199144 189942 199322
rect 190110 199144 191690 199322
rect 191858 199144 193438 199322
rect 193606 199144 195186 199322
rect 195354 199144 196934 199322
rect 197102 199144 198682 199322
rect 198850 199144 199068 199322
rect 1398 856 199068 199144
rect 1398 31 2354 856
rect 2522 31 4286 856
rect 4454 31 6218 856
rect 6386 31 8150 856
rect 8318 31 10082 856
rect 10250 31 12014 856
rect 12182 31 13946 856
rect 14114 31 15878 856
rect 16046 31 17810 856
rect 17978 31 19742 856
rect 19910 31 21674 856
rect 21842 31 23606 856
rect 23774 31 25538 856
rect 25706 31 27470 856
rect 27638 31 29402 856
rect 29570 31 31334 856
rect 31502 31 33266 856
rect 33434 31 35198 856
rect 35366 31 37130 856
rect 37298 31 39062 856
rect 39230 31 40994 856
rect 41162 31 42926 856
rect 43094 31 44858 856
rect 45026 31 46790 856
rect 46958 31 48722 856
rect 48890 31 50654 856
rect 50822 31 52586 856
rect 52754 31 54518 856
rect 54686 31 56450 856
rect 56618 31 58382 856
rect 58550 31 60314 856
rect 60482 31 62246 856
rect 62414 31 64178 856
rect 64346 31 66110 856
rect 66278 31 68042 856
rect 68210 31 69974 856
rect 70142 31 71906 856
rect 72074 31 73838 856
rect 74006 31 75770 856
rect 75938 31 77702 856
rect 77870 31 79634 856
rect 79802 31 81566 856
rect 81734 31 83498 856
rect 83666 31 85430 856
rect 85598 31 87362 856
rect 87530 31 89294 856
rect 89462 31 91226 856
rect 91394 31 93158 856
rect 93326 31 95090 856
rect 95258 31 97022 856
rect 97190 31 98954 856
rect 99122 31 100886 856
rect 101054 31 102818 856
rect 102986 31 104750 856
rect 104918 31 106682 856
rect 106850 31 108614 856
rect 108782 31 110546 856
rect 110714 31 112478 856
rect 112646 31 114410 856
rect 114578 31 116342 856
rect 116510 31 118274 856
rect 118442 31 120206 856
rect 120374 31 122138 856
rect 122306 31 124070 856
rect 124238 31 126002 856
rect 126170 31 127934 856
rect 128102 31 129866 856
rect 130034 31 131798 856
rect 131966 31 133730 856
rect 133898 31 135662 856
rect 135830 31 137594 856
rect 137762 31 139526 856
rect 139694 31 141458 856
rect 141626 31 143390 856
rect 143558 31 145322 856
rect 145490 31 147254 856
rect 147422 31 149186 856
rect 149354 31 151118 856
rect 151286 31 153050 856
rect 153218 31 154982 856
rect 155150 31 156914 856
rect 157082 31 158846 856
rect 159014 31 160778 856
rect 160946 31 162710 856
rect 162878 31 164642 856
rect 164810 31 166574 856
rect 166742 31 168506 856
rect 168674 31 170438 856
rect 170606 31 172370 856
rect 172538 31 174302 856
rect 174470 31 176234 856
rect 176402 31 178166 856
rect 178334 31 180098 856
rect 180266 31 182030 856
rect 182198 31 183962 856
rect 184130 31 185894 856
rect 186062 31 187826 856
rect 187994 31 189758 856
rect 189926 31 191690 856
rect 191858 31 193622 856
rect 193790 31 195554 856
rect 195722 31 197486 856
rect 197654 31 199068 856
<< metal3 >>
rect 0 197480 800 197600
rect 199200 196936 200000 197056
rect 0 192720 800 192840
rect 199200 192312 200000 192432
rect 0 187960 800 188080
rect 199200 187688 200000 187808
rect 0 183200 800 183320
rect 199200 183064 200000 183184
rect 0 178440 800 178560
rect 199200 178440 200000 178560
rect 0 173680 800 173800
rect 199200 173816 200000 173936
rect 199200 169192 200000 169312
rect 0 168920 800 169040
rect 199200 164568 200000 164688
rect 0 164160 800 164280
rect 199200 159944 200000 160064
rect 0 159400 800 159520
rect 199200 155320 200000 155440
rect 0 154640 800 154760
rect 199200 150696 200000 150816
rect 0 149880 800 150000
rect 199200 146072 200000 146192
rect 0 145120 800 145240
rect 199200 141448 200000 141568
rect 0 140360 800 140480
rect 199200 136824 200000 136944
rect 0 135600 800 135720
rect 199200 132200 200000 132320
rect 0 130840 800 130960
rect 199200 127576 200000 127696
rect 0 126080 800 126200
rect 199200 122952 200000 123072
rect 0 121320 800 121440
rect 199200 118328 200000 118448
rect 0 116560 800 116680
rect 199200 113704 200000 113824
rect 0 111800 800 111920
rect 199200 109080 200000 109200
rect 0 107040 800 107160
rect 199200 104456 200000 104576
rect 0 102280 800 102400
rect 199200 99832 200000 99952
rect 0 97520 800 97640
rect 199200 95208 200000 95328
rect 0 92760 800 92880
rect 199200 90584 200000 90704
rect 0 88000 800 88120
rect 199200 85960 200000 86080
rect 0 83240 800 83360
rect 199200 81336 200000 81456
rect 0 78480 800 78600
rect 199200 76712 200000 76832
rect 0 73720 800 73840
rect 199200 72088 200000 72208
rect 0 68960 800 69080
rect 199200 67464 200000 67584
rect 0 64200 800 64320
rect 199200 62840 200000 62960
rect 0 59440 800 59560
rect 199200 58216 200000 58336
rect 0 54680 800 54800
rect 199200 53592 200000 53712
rect 0 49920 800 50040
rect 199200 48968 200000 49088
rect 0 45160 800 45280
rect 199200 44344 200000 44464
rect 0 40400 800 40520
rect 199200 39720 200000 39840
rect 0 35640 800 35760
rect 199200 35096 200000 35216
rect 0 30880 800 31000
rect 199200 30472 200000 30592
rect 0 26120 800 26240
rect 199200 25848 200000 25968
rect 0 21360 800 21480
rect 199200 21224 200000 21344
rect 0 16600 800 16720
rect 199200 16600 200000 16720
rect 0 11840 800 11960
rect 199200 11976 200000 12096
rect 199200 7352 200000 7472
rect 0 7080 800 7200
rect 199200 2728 200000 2848
rect 0 2320 800 2440
<< obsm3 >>
rect 880 197400 199200 197573
rect 800 197136 199200 197400
rect 800 196856 199120 197136
rect 800 192920 199200 196856
rect 880 192640 199200 192920
rect 800 192512 199200 192640
rect 800 192232 199120 192512
rect 800 188160 199200 192232
rect 880 187888 199200 188160
rect 880 187880 199120 187888
rect 800 187608 199120 187880
rect 800 183400 199200 187608
rect 880 183264 199200 183400
rect 880 183120 199120 183264
rect 800 182984 199120 183120
rect 800 178640 199200 182984
rect 880 178360 199120 178640
rect 800 174016 199200 178360
rect 800 173880 199120 174016
rect 880 173736 199120 173880
rect 880 173600 199200 173736
rect 800 169392 199200 173600
rect 800 169120 199120 169392
rect 880 169112 199120 169120
rect 880 168840 199200 169112
rect 800 164768 199200 168840
rect 800 164488 199120 164768
rect 800 164360 199200 164488
rect 880 164080 199200 164360
rect 800 160144 199200 164080
rect 800 159864 199120 160144
rect 800 159600 199200 159864
rect 880 159320 199200 159600
rect 800 155520 199200 159320
rect 800 155240 199120 155520
rect 800 154840 199200 155240
rect 880 154560 199200 154840
rect 800 150896 199200 154560
rect 800 150616 199120 150896
rect 800 150080 199200 150616
rect 880 149800 199200 150080
rect 800 146272 199200 149800
rect 800 145992 199120 146272
rect 800 145320 199200 145992
rect 880 145040 199200 145320
rect 800 141648 199200 145040
rect 800 141368 199120 141648
rect 800 140560 199200 141368
rect 880 140280 199200 140560
rect 800 137024 199200 140280
rect 800 136744 199120 137024
rect 800 135800 199200 136744
rect 880 135520 199200 135800
rect 800 132400 199200 135520
rect 800 132120 199120 132400
rect 800 131040 199200 132120
rect 880 130760 199200 131040
rect 800 127776 199200 130760
rect 800 127496 199120 127776
rect 800 126280 199200 127496
rect 880 126000 199200 126280
rect 800 123152 199200 126000
rect 800 122872 199120 123152
rect 800 121520 199200 122872
rect 880 121240 199200 121520
rect 800 118528 199200 121240
rect 800 118248 199120 118528
rect 800 116760 199200 118248
rect 880 116480 199200 116760
rect 800 113904 199200 116480
rect 800 113624 199120 113904
rect 800 112000 199200 113624
rect 880 111720 199200 112000
rect 800 109280 199200 111720
rect 800 109000 199120 109280
rect 800 107240 199200 109000
rect 880 106960 199200 107240
rect 800 104656 199200 106960
rect 800 104376 199120 104656
rect 800 102480 199200 104376
rect 880 102200 199200 102480
rect 800 100032 199200 102200
rect 800 99752 199120 100032
rect 800 97720 199200 99752
rect 880 97440 199200 97720
rect 800 95408 199200 97440
rect 800 95128 199120 95408
rect 800 92960 199200 95128
rect 880 92680 199200 92960
rect 800 90784 199200 92680
rect 800 90504 199120 90784
rect 800 88200 199200 90504
rect 880 87920 199200 88200
rect 800 86160 199200 87920
rect 800 85880 199120 86160
rect 800 83440 199200 85880
rect 880 83160 199200 83440
rect 800 81536 199200 83160
rect 800 81256 199120 81536
rect 800 78680 199200 81256
rect 880 78400 199200 78680
rect 800 76912 199200 78400
rect 800 76632 199120 76912
rect 800 73920 199200 76632
rect 880 73640 199200 73920
rect 800 72288 199200 73640
rect 800 72008 199120 72288
rect 800 69160 199200 72008
rect 880 68880 199200 69160
rect 800 67664 199200 68880
rect 800 67384 199120 67664
rect 800 64400 199200 67384
rect 880 64120 199200 64400
rect 800 63040 199200 64120
rect 800 62760 199120 63040
rect 800 59640 199200 62760
rect 880 59360 199200 59640
rect 800 58416 199200 59360
rect 800 58136 199120 58416
rect 800 54880 199200 58136
rect 880 54600 199200 54880
rect 800 53792 199200 54600
rect 800 53512 199120 53792
rect 800 50120 199200 53512
rect 880 49840 199200 50120
rect 800 49168 199200 49840
rect 800 48888 199120 49168
rect 800 45360 199200 48888
rect 880 45080 199200 45360
rect 800 44544 199200 45080
rect 800 44264 199120 44544
rect 800 40600 199200 44264
rect 880 40320 199200 40600
rect 800 39920 199200 40320
rect 800 39640 199120 39920
rect 800 35840 199200 39640
rect 880 35560 199200 35840
rect 800 35296 199200 35560
rect 800 35016 199120 35296
rect 800 31080 199200 35016
rect 880 30800 199200 31080
rect 800 30672 199200 30800
rect 800 30392 199120 30672
rect 800 26320 199200 30392
rect 880 26048 199200 26320
rect 880 26040 199120 26048
rect 800 25768 199120 26040
rect 800 21560 199200 25768
rect 880 21424 199200 21560
rect 880 21280 199120 21424
rect 800 21144 199120 21280
rect 800 16800 199200 21144
rect 880 16520 199120 16800
rect 800 12176 199200 16520
rect 800 12040 199120 12176
rect 880 11896 199120 12040
rect 880 11760 199200 11896
rect 800 7552 199200 11760
rect 800 7280 199120 7552
rect 880 7272 199120 7280
rect 880 7000 199200 7272
rect 800 2928 199200 7000
rect 800 2648 199120 2928
rect 800 2520 199200 2648
rect 880 2240 199200 2520
rect 800 35 199200 2240
<< metal4 >>
rect 4208 2128 4528 197520
rect 19568 2128 19888 197520
rect 34928 2128 35248 197520
rect 50288 2128 50608 197520
rect 65648 2128 65968 197520
rect 81008 2128 81328 197520
rect 96368 2128 96688 197520
rect 111728 2128 112048 197520
rect 127088 2128 127408 197520
rect 142448 2128 142768 197520
rect 157808 2128 158128 197520
rect 173168 2128 173488 197520
rect 188528 2128 188848 197520
<< obsm4 >>
rect 1715 2048 4128 197301
rect 4608 2048 19488 197301
rect 19968 2048 34848 197301
rect 35328 2048 50208 197301
rect 50688 2048 65568 197301
rect 66048 2048 80928 197301
rect 81408 2048 96288 197301
rect 96768 2048 111648 197301
rect 112128 2048 127008 197301
rect 127488 2048 142368 197301
rect 142848 2048 157728 197301
rect 158208 2048 161493 197301
rect 1715 35 161493 2048
<< labels >>
rlabel metal2 s 1214 199200 1270 200000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 53654 199200 53710 200000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 58898 199200 58954 200000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 64142 199200 64198 200000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 69386 199200 69442 200000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 74630 199200 74686 200000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 79874 199200 79930 200000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 85118 199200 85174 200000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 90362 199200 90418 200000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 95606 199200 95662 200000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 100850 199200 100906 200000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 6458 199200 6514 200000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 106094 199200 106150 200000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 111338 199200 111394 200000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 116582 199200 116638 200000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 121826 199200 121882 200000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 127070 199200 127126 200000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 132314 199200 132370 200000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 137558 199200 137614 200000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 142802 199200 142858 200000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 148046 199200 148102 200000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 153290 199200 153346 200000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 11702 199200 11758 200000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 158534 199200 158590 200000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 163778 199200 163834 200000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 169022 199200 169078 200000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 174266 199200 174322 200000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 179510 199200 179566 200000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 184754 199200 184810 200000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 189998 199200 190054 200000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 195242 199200 195298 200000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 16946 199200 17002 200000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 22190 199200 22246 200000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 27434 199200 27490 200000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 32678 199200 32734 200000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 37922 199200 37978 200000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 43166 199200 43222 200000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 48410 199200 48466 200000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 2962 199200 3018 200000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 55402 199200 55458 200000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 60646 199200 60702 200000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 65890 199200 65946 200000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 71134 199200 71190 200000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 76378 199200 76434 200000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 81622 199200 81678 200000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 86866 199200 86922 200000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 92110 199200 92166 200000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 97354 199200 97410 200000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 102598 199200 102654 200000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 8206 199200 8262 200000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 107842 199200 107898 200000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 113086 199200 113142 200000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 118330 199200 118386 200000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 123574 199200 123630 200000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 128818 199200 128874 200000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 134062 199200 134118 200000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 139306 199200 139362 200000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 144550 199200 144606 200000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 149794 199200 149850 200000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 155038 199200 155094 200000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 13450 199200 13506 200000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 160282 199200 160338 200000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 165526 199200 165582 200000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 170770 199200 170826 200000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 176014 199200 176070 200000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 181258 199200 181314 200000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 186502 199200 186558 200000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 191746 199200 191802 200000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 196990 199200 197046 200000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 18694 199200 18750 200000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 23938 199200 23994 200000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 29182 199200 29238 200000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 34426 199200 34482 200000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 39670 199200 39726 200000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 44914 199200 44970 200000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 50158 199200 50214 200000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 4710 199200 4766 200000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 57150 199200 57206 200000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 62394 199200 62450 200000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 67638 199200 67694 200000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 72882 199200 72938 200000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 78126 199200 78182 200000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 83370 199200 83426 200000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 88614 199200 88670 200000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 93858 199200 93914 200000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 99102 199200 99158 200000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 104346 199200 104402 200000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 9954 199200 10010 200000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 109590 199200 109646 200000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 114834 199200 114890 200000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 120078 199200 120134 200000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 125322 199200 125378 200000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 130566 199200 130622 200000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 135810 199200 135866 200000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 141054 199200 141110 200000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 146298 199200 146354 200000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 151542 199200 151598 200000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 156786 199200 156842 200000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 15198 199200 15254 200000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 162030 199200 162086 200000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 167274 199200 167330 200000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 172518 199200 172574 200000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 177762 199200 177818 200000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 183006 199200 183062 200000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 188250 199200 188306 200000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 193494 199200 193550 200000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 198738 199200 198794 200000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 20442 199200 20498 200000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 25686 199200 25742 200000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 30930 199200 30986 200000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 36174 199200 36230 200000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 41418 199200 41474 200000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 46662 199200 46718 200000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 51906 199200 51962 200000 6 io_out[9]
port 114 nsew signal output
rlabel metal3 s 0 7080 800 7200 6 oram_addr[0]
port 115 nsew signal output
rlabel metal3 s 0 16600 800 16720 6 oram_addr[1]
port 116 nsew signal output
rlabel metal3 s 0 26120 800 26240 6 oram_addr[2]
port 117 nsew signal output
rlabel metal3 s 0 35640 800 35760 6 oram_addr[3]
port 118 nsew signal output
rlabel metal3 s 0 45160 800 45280 6 oram_addr[4]
port 119 nsew signal output
rlabel metal3 s 0 54680 800 54800 6 oram_addr[5]
port 120 nsew signal output
rlabel metal3 s 0 64200 800 64320 6 oram_addr[6]
port 121 nsew signal output
rlabel metal3 s 0 73720 800 73840 6 oram_addr[7]
port 122 nsew signal output
rlabel metal3 s 0 83240 800 83360 6 oram_addr[8]
port 123 nsew signal output
rlabel metal3 s 0 2320 800 2440 6 oram_csb
port 124 nsew signal output
rlabel metal3 s 0 11840 800 11960 6 oram_value[0]
port 125 nsew signal input
rlabel metal3 s 0 97520 800 97640 6 oram_value[10]
port 126 nsew signal input
rlabel metal3 s 0 102280 800 102400 6 oram_value[11]
port 127 nsew signal input
rlabel metal3 s 0 107040 800 107160 6 oram_value[12]
port 128 nsew signal input
rlabel metal3 s 0 111800 800 111920 6 oram_value[13]
port 129 nsew signal input
rlabel metal3 s 0 116560 800 116680 6 oram_value[14]
port 130 nsew signal input
rlabel metal3 s 0 121320 800 121440 6 oram_value[15]
port 131 nsew signal input
rlabel metal3 s 0 126080 800 126200 6 oram_value[16]
port 132 nsew signal input
rlabel metal3 s 0 130840 800 130960 6 oram_value[17]
port 133 nsew signal input
rlabel metal3 s 0 135600 800 135720 6 oram_value[18]
port 134 nsew signal input
rlabel metal3 s 0 140360 800 140480 6 oram_value[19]
port 135 nsew signal input
rlabel metal3 s 0 21360 800 21480 6 oram_value[1]
port 136 nsew signal input
rlabel metal3 s 0 145120 800 145240 6 oram_value[20]
port 137 nsew signal input
rlabel metal3 s 0 149880 800 150000 6 oram_value[21]
port 138 nsew signal input
rlabel metal3 s 0 154640 800 154760 6 oram_value[22]
port 139 nsew signal input
rlabel metal3 s 0 159400 800 159520 6 oram_value[23]
port 140 nsew signal input
rlabel metal3 s 0 164160 800 164280 6 oram_value[24]
port 141 nsew signal input
rlabel metal3 s 0 168920 800 169040 6 oram_value[25]
port 142 nsew signal input
rlabel metal3 s 0 173680 800 173800 6 oram_value[26]
port 143 nsew signal input
rlabel metal3 s 0 178440 800 178560 6 oram_value[27]
port 144 nsew signal input
rlabel metal3 s 0 183200 800 183320 6 oram_value[28]
port 145 nsew signal input
rlabel metal3 s 0 187960 800 188080 6 oram_value[29]
port 146 nsew signal input
rlabel metal3 s 0 30880 800 31000 6 oram_value[2]
port 147 nsew signal input
rlabel metal3 s 0 192720 800 192840 6 oram_value[30]
port 148 nsew signal input
rlabel metal3 s 0 197480 800 197600 6 oram_value[31]
port 149 nsew signal input
rlabel metal3 s 0 40400 800 40520 6 oram_value[3]
port 150 nsew signal input
rlabel metal3 s 0 49920 800 50040 6 oram_value[4]
port 151 nsew signal input
rlabel metal3 s 0 59440 800 59560 6 oram_value[5]
port 152 nsew signal input
rlabel metal3 s 0 68960 800 69080 6 oram_value[6]
port 153 nsew signal input
rlabel metal3 s 0 78480 800 78600 6 oram_value[7]
port 154 nsew signal input
rlabel metal3 s 0 88000 800 88120 6 oram_value[8]
port 155 nsew signal input
rlabel metal3 s 0 92760 800 92880 6 oram_value[9]
port 156 nsew signal input
rlabel metal3 s 199200 11976 200000 12096 6 ram_adrb[0]
port 157 nsew signal output
rlabel metal3 s 199200 21224 200000 21344 6 ram_adrb[1]
port 158 nsew signal output
rlabel metal3 s 199200 30472 200000 30592 6 ram_adrb[2]
port 159 nsew signal output
rlabel metal3 s 199200 39720 200000 39840 6 ram_adrb[3]
port 160 nsew signal output
rlabel metal3 s 199200 48968 200000 49088 6 ram_adrb[4]
port 161 nsew signal output
rlabel metal3 s 199200 58216 200000 58336 6 ram_adrb[5]
port 162 nsew signal output
rlabel metal3 s 199200 67464 200000 67584 6 ram_adrb[6]
port 163 nsew signal output
rlabel metal3 s 199200 76712 200000 76832 6 ram_adrb[7]
port 164 nsew signal output
rlabel metal3 s 199200 85960 200000 86080 6 ram_adrb[8]
port 165 nsew signal output
rlabel metal3 s 199200 2728 200000 2848 6 ram_csb
port 166 nsew signal output
rlabel metal3 s 199200 16600 200000 16720 6 ram_val[0]
port 167 nsew signal input
rlabel metal3 s 199200 99832 200000 99952 6 ram_val[10]
port 168 nsew signal input
rlabel metal3 s 199200 104456 200000 104576 6 ram_val[11]
port 169 nsew signal input
rlabel metal3 s 199200 109080 200000 109200 6 ram_val[12]
port 170 nsew signal input
rlabel metal3 s 199200 113704 200000 113824 6 ram_val[13]
port 171 nsew signal input
rlabel metal3 s 199200 118328 200000 118448 6 ram_val[14]
port 172 nsew signal input
rlabel metal3 s 199200 122952 200000 123072 6 ram_val[15]
port 173 nsew signal input
rlabel metal3 s 199200 127576 200000 127696 6 ram_val[16]
port 174 nsew signal input
rlabel metal3 s 199200 132200 200000 132320 6 ram_val[17]
port 175 nsew signal input
rlabel metal3 s 199200 136824 200000 136944 6 ram_val[18]
port 176 nsew signal input
rlabel metal3 s 199200 141448 200000 141568 6 ram_val[19]
port 177 nsew signal input
rlabel metal3 s 199200 25848 200000 25968 6 ram_val[1]
port 178 nsew signal input
rlabel metal3 s 199200 146072 200000 146192 6 ram_val[20]
port 179 nsew signal input
rlabel metal3 s 199200 150696 200000 150816 6 ram_val[21]
port 180 nsew signal input
rlabel metal3 s 199200 155320 200000 155440 6 ram_val[22]
port 181 nsew signal input
rlabel metal3 s 199200 159944 200000 160064 6 ram_val[23]
port 182 nsew signal input
rlabel metal3 s 199200 164568 200000 164688 6 ram_val[24]
port 183 nsew signal input
rlabel metal3 s 199200 169192 200000 169312 6 ram_val[25]
port 184 nsew signal input
rlabel metal3 s 199200 173816 200000 173936 6 ram_val[26]
port 185 nsew signal input
rlabel metal3 s 199200 178440 200000 178560 6 ram_val[27]
port 186 nsew signal input
rlabel metal3 s 199200 183064 200000 183184 6 ram_val[28]
port 187 nsew signal input
rlabel metal3 s 199200 187688 200000 187808 6 ram_val[29]
port 188 nsew signal input
rlabel metal3 s 199200 35096 200000 35216 6 ram_val[2]
port 189 nsew signal input
rlabel metal3 s 199200 192312 200000 192432 6 ram_val[30]
port 190 nsew signal input
rlabel metal3 s 199200 196936 200000 197056 6 ram_val[31]
port 191 nsew signal input
rlabel metal3 s 199200 44344 200000 44464 6 ram_val[3]
port 192 nsew signal input
rlabel metal3 s 199200 53592 200000 53712 6 ram_val[4]
port 193 nsew signal input
rlabel metal3 s 199200 62840 200000 62960 6 ram_val[5]
port 194 nsew signal input
rlabel metal3 s 199200 72088 200000 72208 6 ram_val[6]
port 195 nsew signal input
rlabel metal3 s 199200 81336 200000 81456 6 ram_val[7]
port 196 nsew signal input
rlabel metal3 s 199200 90584 200000 90704 6 ram_val[8]
port 197 nsew signal input
rlabel metal3 s 199200 95208 200000 95328 6 ram_val[9]
port 198 nsew signal input
rlabel metal3 s 199200 7352 200000 7472 6 ram_web
port 199 nsew signal output
rlabel metal4 s 4208 2128 4528 197520 6 vccd1
port 200 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 197520 6 vccd1
port 200 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 197520 6 vccd1
port 200 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 197520 6 vccd1
port 200 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 197520 6 vccd1
port 200 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 197520 6 vccd1
port 200 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 197520 6 vccd1
port 200 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 197520 6 vssd1
port 201 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 197520 6 vssd1
port 201 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 197520 6 vssd1
port 201 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 197520 6 vssd1
port 201 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 197520 6 vssd1
port 201 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 197520 6 vssd1
port 201 nsew ground bidirectional
rlabel metal2 s 2410 0 2466 800 6 wb_clk_i
port 202 nsew signal input
rlabel metal2 s 4342 0 4398 800 6 wb_rst_i
port 203 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 wbs_ack_o
port 204 nsew signal output
rlabel metal2 s 14002 0 14058 800 6 wbs_adr_i[0]
port 205 nsew signal input
rlabel metal2 s 71962 0 72018 800 6 wbs_adr_i[10]
port 206 nsew signal input
rlabel metal2 s 77758 0 77814 800 6 wbs_adr_i[11]
port 207 nsew signal input
rlabel metal2 s 83554 0 83610 800 6 wbs_adr_i[12]
port 208 nsew signal input
rlabel metal2 s 89350 0 89406 800 6 wbs_adr_i[13]
port 209 nsew signal input
rlabel metal2 s 95146 0 95202 800 6 wbs_adr_i[14]
port 210 nsew signal input
rlabel metal2 s 100942 0 100998 800 6 wbs_adr_i[15]
port 211 nsew signal input
rlabel metal2 s 106738 0 106794 800 6 wbs_adr_i[16]
port 212 nsew signal input
rlabel metal2 s 112534 0 112590 800 6 wbs_adr_i[17]
port 213 nsew signal input
rlabel metal2 s 118330 0 118386 800 6 wbs_adr_i[18]
port 214 nsew signal input
rlabel metal2 s 124126 0 124182 800 6 wbs_adr_i[19]
port 215 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 wbs_adr_i[1]
port 216 nsew signal input
rlabel metal2 s 129922 0 129978 800 6 wbs_adr_i[20]
port 217 nsew signal input
rlabel metal2 s 135718 0 135774 800 6 wbs_adr_i[21]
port 218 nsew signal input
rlabel metal2 s 141514 0 141570 800 6 wbs_adr_i[22]
port 219 nsew signal input
rlabel metal2 s 147310 0 147366 800 6 wbs_adr_i[23]
port 220 nsew signal input
rlabel metal2 s 153106 0 153162 800 6 wbs_adr_i[24]
port 221 nsew signal input
rlabel metal2 s 158902 0 158958 800 6 wbs_adr_i[25]
port 222 nsew signal input
rlabel metal2 s 164698 0 164754 800 6 wbs_adr_i[26]
port 223 nsew signal input
rlabel metal2 s 170494 0 170550 800 6 wbs_adr_i[27]
port 224 nsew signal input
rlabel metal2 s 176290 0 176346 800 6 wbs_adr_i[28]
port 225 nsew signal input
rlabel metal2 s 182086 0 182142 800 6 wbs_adr_i[29]
port 226 nsew signal input
rlabel metal2 s 25594 0 25650 800 6 wbs_adr_i[2]
port 227 nsew signal input
rlabel metal2 s 187882 0 187938 800 6 wbs_adr_i[30]
port 228 nsew signal input
rlabel metal2 s 193678 0 193734 800 6 wbs_adr_i[31]
port 229 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 wbs_adr_i[3]
port 230 nsew signal input
rlabel metal2 s 37186 0 37242 800 6 wbs_adr_i[4]
port 231 nsew signal input
rlabel metal2 s 42982 0 43038 800 6 wbs_adr_i[5]
port 232 nsew signal input
rlabel metal2 s 48778 0 48834 800 6 wbs_adr_i[6]
port 233 nsew signal input
rlabel metal2 s 54574 0 54630 800 6 wbs_adr_i[7]
port 234 nsew signal input
rlabel metal2 s 60370 0 60426 800 6 wbs_adr_i[8]
port 235 nsew signal input
rlabel metal2 s 66166 0 66222 800 6 wbs_adr_i[9]
port 236 nsew signal input
rlabel metal2 s 8206 0 8262 800 6 wbs_cyc_i
port 237 nsew signal input
rlabel metal2 s 15934 0 15990 800 6 wbs_dat_i[0]
port 238 nsew signal input
rlabel metal2 s 73894 0 73950 800 6 wbs_dat_i[10]
port 239 nsew signal input
rlabel metal2 s 79690 0 79746 800 6 wbs_dat_i[11]
port 240 nsew signal input
rlabel metal2 s 85486 0 85542 800 6 wbs_dat_i[12]
port 241 nsew signal input
rlabel metal2 s 91282 0 91338 800 6 wbs_dat_i[13]
port 242 nsew signal input
rlabel metal2 s 97078 0 97134 800 6 wbs_dat_i[14]
port 243 nsew signal input
rlabel metal2 s 102874 0 102930 800 6 wbs_dat_i[15]
port 244 nsew signal input
rlabel metal2 s 108670 0 108726 800 6 wbs_dat_i[16]
port 245 nsew signal input
rlabel metal2 s 114466 0 114522 800 6 wbs_dat_i[17]
port 246 nsew signal input
rlabel metal2 s 120262 0 120318 800 6 wbs_dat_i[18]
port 247 nsew signal input
rlabel metal2 s 126058 0 126114 800 6 wbs_dat_i[19]
port 248 nsew signal input
rlabel metal2 s 21730 0 21786 800 6 wbs_dat_i[1]
port 249 nsew signal input
rlabel metal2 s 131854 0 131910 800 6 wbs_dat_i[20]
port 250 nsew signal input
rlabel metal2 s 137650 0 137706 800 6 wbs_dat_i[21]
port 251 nsew signal input
rlabel metal2 s 143446 0 143502 800 6 wbs_dat_i[22]
port 252 nsew signal input
rlabel metal2 s 149242 0 149298 800 6 wbs_dat_i[23]
port 253 nsew signal input
rlabel metal2 s 155038 0 155094 800 6 wbs_dat_i[24]
port 254 nsew signal input
rlabel metal2 s 160834 0 160890 800 6 wbs_dat_i[25]
port 255 nsew signal input
rlabel metal2 s 166630 0 166686 800 6 wbs_dat_i[26]
port 256 nsew signal input
rlabel metal2 s 172426 0 172482 800 6 wbs_dat_i[27]
port 257 nsew signal input
rlabel metal2 s 178222 0 178278 800 6 wbs_dat_i[28]
port 258 nsew signal input
rlabel metal2 s 184018 0 184074 800 6 wbs_dat_i[29]
port 259 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 wbs_dat_i[2]
port 260 nsew signal input
rlabel metal2 s 189814 0 189870 800 6 wbs_dat_i[30]
port 261 nsew signal input
rlabel metal2 s 195610 0 195666 800 6 wbs_dat_i[31]
port 262 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 wbs_dat_i[3]
port 263 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 wbs_dat_i[4]
port 264 nsew signal input
rlabel metal2 s 44914 0 44970 800 6 wbs_dat_i[5]
port 265 nsew signal input
rlabel metal2 s 50710 0 50766 800 6 wbs_dat_i[6]
port 266 nsew signal input
rlabel metal2 s 56506 0 56562 800 6 wbs_dat_i[7]
port 267 nsew signal input
rlabel metal2 s 62302 0 62358 800 6 wbs_dat_i[8]
port 268 nsew signal input
rlabel metal2 s 68098 0 68154 800 6 wbs_dat_i[9]
port 269 nsew signal input
rlabel metal2 s 17866 0 17922 800 6 wbs_dat_o[0]
port 270 nsew signal output
rlabel metal2 s 75826 0 75882 800 6 wbs_dat_o[10]
port 271 nsew signal output
rlabel metal2 s 81622 0 81678 800 6 wbs_dat_o[11]
port 272 nsew signal output
rlabel metal2 s 87418 0 87474 800 6 wbs_dat_o[12]
port 273 nsew signal output
rlabel metal2 s 93214 0 93270 800 6 wbs_dat_o[13]
port 274 nsew signal output
rlabel metal2 s 99010 0 99066 800 6 wbs_dat_o[14]
port 275 nsew signal output
rlabel metal2 s 104806 0 104862 800 6 wbs_dat_o[15]
port 276 nsew signal output
rlabel metal2 s 110602 0 110658 800 6 wbs_dat_o[16]
port 277 nsew signal output
rlabel metal2 s 116398 0 116454 800 6 wbs_dat_o[17]
port 278 nsew signal output
rlabel metal2 s 122194 0 122250 800 6 wbs_dat_o[18]
port 279 nsew signal output
rlabel metal2 s 127990 0 128046 800 6 wbs_dat_o[19]
port 280 nsew signal output
rlabel metal2 s 23662 0 23718 800 6 wbs_dat_o[1]
port 281 nsew signal output
rlabel metal2 s 133786 0 133842 800 6 wbs_dat_o[20]
port 282 nsew signal output
rlabel metal2 s 139582 0 139638 800 6 wbs_dat_o[21]
port 283 nsew signal output
rlabel metal2 s 145378 0 145434 800 6 wbs_dat_o[22]
port 284 nsew signal output
rlabel metal2 s 151174 0 151230 800 6 wbs_dat_o[23]
port 285 nsew signal output
rlabel metal2 s 156970 0 157026 800 6 wbs_dat_o[24]
port 286 nsew signal output
rlabel metal2 s 162766 0 162822 800 6 wbs_dat_o[25]
port 287 nsew signal output
rlabel metal2 s 168562 0 168618 800 6 wbs_dat_o[26]
port 288 nsew signal output
rlabel metal2 s 174358 0 174414 800 6 wbs_dat_o[27]
port 289 nsew signal output
rlabel metal2 s 180154 0 180210 800 6 wbs_dat_o[28]
port 290 nsew signal output
rlabel metal2 s 185950 0 186006 800 6 wbs_dat_o[29]
port 291 nsew signal output
rlabel metal2 s 29458 0 29514 800 6 wbs_dat_o[2]
port 292 nsew signal output
rlabel metal2 s 191746 0 191802 800 6 wbs_dat_o[30]
port 293 nsew signal output
rlabel metal2 s 197542 0 197598 800 6 wbs_dat_o[31]
port 294 nsew signal output
rlabel metal2 s 35254 0 35310 800 6 wbs_dat_o[3]
port 295 nsew signal output
rlabel metal2 s 41050 0 41106 800 6 wbs_dat_o[4]
port 296 nsew signal output
rlabel metal2 s 46846 0 46902 800 6 wbs_dat_o[5]
port 297 nsew signal output
rlabel metal2 s 52642 0 52698 800 6 wbs_dat_o[6]
port 298 nsew signal output
rlabel metal2 s 58438 0 58494 800 6 wbs_dat_o[7]
port 299 nsew signal output
rlabel metal2 s 64234 0 64290 800 6 wbs_dat_o[8]
port 300 nsew signal output
rlabel metal2 s 70030 0 70086 800 6 wbs_dat_o[9]
port 301 nsew signal output
rlabel metal2 s 10138 0 10194 800 6 wbs_stb_i
port 302 nsew signal input
rlabel metal2 s 12070 0 12126 800 6 wbs_we_i
port 303 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 200000 200000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 63695888
string GDS_FILE /home/tholin/mpw-8-as1x00/openlane/wrapped_tms1x00/runs/22_12_30_19_52/results/signoff/wrapped_tms1x00.magic.gds
string GDS_START 901654
<< end >>

