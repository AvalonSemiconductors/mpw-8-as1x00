magic
tech sky130B
magscale 1 2
timestamp 1674150506
<< obsli1 >>
rect 1104 2159 148856 137649
<< obsm1 >>
rect 566 8 148856 137680
<< metal2 >>
rect 2134 139200 2190 140000
rect 3422 139200 3478 140000
rect 4710 139200 4766 140000
rect 5998 139200 6054 140000
rect 7286 139200 7342 140000
rect 8574 139200 8630 140000
rect 9862 139200 9918 140000
rect 11150 139200 11206 140000
rect 12438 139200 12494 140000
rect 13726 139200 13782 140000
rect 15014 139200 15070 140000
rect 16302 139200 16358 140000
rect 17590 139200 17646 140000
rect 18878 139200 18934 140000
rect 20166 139200 20222 140000
rect 21454 139200 21510 140000
rect 22742 139200 22798 140000
rect 24030 139200 24086 140000
rect 25318 139200 25374 140000
rect 26606 139200 26662 140000
rect 27894 139200 27950 140000
rect 29182 139200 29238 140000
rect 30470 139200 30526 140000
rect 31758 139200 31814 140000
rect 33046 139200 33102 140000
rect 34334 139200 34390 140000
rect 35622 139200 35678 140000
rect 36910 139200 36966 140000
rect 38198 139200 38254 140000
rect 39486 139200 39542 140000
rect 40774 139200 40830 140000
rect 42062 139200 42118 140000
rect 43350 139200 43406 140000
rect 44638 139200 44694 140000
rect 45926 139200 45982 140000
rect 47214 139200 47270 140000
rect 48502 139200 48558 140000
rect 49790 139200 49846 140000
rect 51078 139200 51134 140000
rect 52366 139200 52422 140000
rect 53654 139200 53710 140000
rect 54942 139200 54998 140000
rect 56230 139200 56286 140000
rect 57518 139200 57574 140000
rect 58806 139200 58862 140000
rect 60094 139200 60150 140000
rect 61382 139200 61438 140000
rect 62670 139200 62726 140000
rect 63958 139200 64014 140000
rect 65246 139200 65302 140000
rect 66534 139200 66590 140000
rect 67822 139200 67878 140000
rect 69110 139200 69166 140000
rect 70398 139200 70454 140000
rect 71686 139200 71742 140000
rect 72974 139200 73030 140000
rect 74262 139200 74318 140000
rect 75550 139200 75606 140000
rect 76838 139200 76894 140000
rect 78126 139200 78182 140000
rect 79414 139200 79470 140000
rect 80702 139200 80758 140000
rect 81990 139200 82046 140000
rect 83278 139200 83334 140000
rect 84566 139200 84622 140000
rect 85854 139200 85910 140000
rect 87142 139200 87198 140000
rect 88430 139200 88486 140000
rect 89718 139200 89774 140000
rect 91006 139200 91062 140000
rect 92294 139200 92350 140000
rect 93582 139200 93638 140000
rect 94870 139200 94926 140000
rect 96158 139200 96214 140000
rect 97446 139200 97502 140000
rect 98734 139200 98790 140000
rect 100022 139200 100078 140000
rect 101310 139200 101366 140000
rect 102598 139200 102654 140000
rect 103886 139200 103942 140000
rect 105174 139200 105230 140000
rect 106462 139200 106518 140000
rect 107750 139200 107806 140000
rect 109038 139200 109094 140000
rect 110326 139200 110382 140000
rect 111614 139200 111670 140000
rect 112902 139200 112958 140000
rect 114190 139200 114246 140000
rect 115478 139200 115534 140000
rect 116766 139200 116822 140000
rect 118054 139200 118110 140000
rect 119342 139200 119398 140000
rect 120630 139200 120686 140000
rect 121918 139200 121974 140000
rect 123206 139200 123262 140000
rect 124494 139200 124550 140000
rect 125782 139200 125838 140000
rect 127070 139200 127126 140000
rect 128358 139200 128414 140000
rect 129646 139200 129702 140000
rect 130934 139200 130990 140000
rect 132222 139200 132278 140000
rect 133510 139200 133566 140000
rect 134798 139200 134854 140000
rect 136086 139200 136142 140000
rect 137374 139200 137430 140000
rect 138662 139200 138718 140000
rect 139950 139200 140006 140000
rect 141238 139200 141294 140000
rect 142526 139200 142582 140000
rect 143814 139200 143870 140000
rect 145102 139200 145158 140000
rect 146390 139200 146446 140000
rect 147678 139200 147734 140000
rect 2042 0 2098 800
rect 3054 0 3110 800
rect 4066 0 4122 800
rect 5078 0 5134 800
rect 6090 0 6146 800
rect 7102 0 7158 800
rect 8114 0 8170 800
rect 9126 0 9182 800
rect 10138 0 10194 800
rect 11150 0 11206 800
rect 12162 0 12218 800
rect 13174 0 13230 800
rect 14186 0 14242 800
rect 15198 0 15254 800
rect 16210 0 16266 800
rect 17222 0 17278 800
rect 18234 0 18290 800
rect 19246 0 19302 800
rect 20258 0 20314 800
rect 21270 0 21326 800
rect 22282 0 22338 800
rect 23294 0 23350 800
rect 24306 0 24362 800
rect 25318 0 25374 800
rect 26330 0 26386 800
rect 27342 0 27398 800
rect 28354 0 28410 800
rect 29366 0 29422 800
rect 30378 0 30434 800
rect 31390 0 31446 800
rect 32402 0 32458 800
rect 33414 0 33470 800
rect 34426 0 34482 800
rect 35438 0 35494 800
rect 36450 0 36506 800
rect 37462 0 37518 800
rect 38474 0 38530 800
rect 39486 0 39542 800
rect 40498 0 40554 800
rect 41510 0 41566 800
rect 42522 0 42578 800
rect 43534 0 43590 800
rect 44546 0 44602 800
rect 45558 0 45614 800
rect 46570 0 46626 800
rect 47582 0 47638 800
rect 48594 0 48650 800
rect 49606 0 49662 800
rect 50618 0 50674 800
rect 51630 0 51686 800
rect 52642 0 52698 800
rect 53654 0 53710 800
rect 54666 0 54722 800
rect 55678 0 55734 800
rect 56690 0 56746 800
rect 57702 0 57758 800
rect 58714 0 58770 800
rect 59726 0 59782 800
rect 60738 0 60794 800
rect 61750 0 61806 800
rect 62762 0 62818 800
rect 63774 0 63830 800
rect 64786 0 64842 800
rect 65798 0 65854 800
rect 66810 0 66866 800
rect 67822 0 67878 800
rect 68834 0 68890 800
rect 69846 0 69902 800
rect 70858 0 70914 800
rect 71870 0 71926 800
rect 72882 0 72938 800
rect 73894 0 73950 800
rect 74906 0 74962 800
rect 75918 0 75974 800
rect 76930 0 76986 800
rect 77942 0 77998 800
rect 78954 0 79010 800
rect 79966 0 80022 800
rect 80978 0 81034 800
rect 81990 0 82046 800
rect 83002 0 83058 800
rect 84014 0 84070 800
rect 85026 0 85082 800
rect 86038 0 86094 800
rect 87050 0 87106 800
rect 88062 0 88118 800
rect 89074 0 89130 800
rect 90086 0 90142 800
rect 91098 0 91154 800
rect 92110 0 92166 800
rect 93122 0 93178 800
rect 94134 0 94190 800
rect 95146 0 95202 800
rect 96158 0 96214 800
rect 97170 0 97226 800
rect 98182 0 98238 800
rect 99194 0 99250 800
rect 100206 0 100262 800
rect 101218 0 101274 800
rect 102230 0 102286 800
rect 103242 0 103298 800
rect 104254 0 104310 800
rect 105266 0 105322 800
rect 106278 0 106334 800
rect 107290 0 107346 800
rect 108302 0 108358 800
rect 109314 0 109370 800
rect 110326 0 110382 800
rect 111338 0 111394 800
rect 112350 0 112406 800
rect 113362 0 113418 800
rect 114374 0 114430 800
rect 115386 0 115442 800
rect 116398 0 116454 800
rect 117410 0 117466 800
rect 118422 0 118478 800
rect 119434 0 119490 800
rect 120446 0 120502 800
rect 121458 0 121514 800
rect 122470 0 122526 800
rect 123482 0 123538 800
rect 124494 0 124550 800
rect 125506 0 125562 800
rect 126518 0 126574 800
rect 127530 0 127586 800
rect 128542 0 128598 800
rect 129554 0 129610 800
rect 130566 0 130622 800
rect 131578 0 131634 800
rect 132590 0 132646 800
rect 133602 0 133658 800
rect 134614 0 134670 800
rect 135626 0 135682 800
rect 136638 0 136694 800
rect 137650 0 137706 800
rect 138662 0 138718 800
rect 139674 0 139730 800
rect 140686 0 140742 800
rect 141698 0 141754 800
rect 142710 0 142766 800
rect 143722 0 143778 800
rect 144734 0 144790 800
rect 145746 0 145802 800
rect 146758 0 146814 800
rect 147770 0 147826 800
<< obsm2 >>
rect 478 139144 2078 139346
rect 2246 139144 3366 139346
rect 3534 139144 4654 139346
rect 4822 139144 5942 139346
rect 6110 139144 7230 139346
rect 7398 139144 8518 139346
rect 8686 139144 9806 139346
rect 9974 139144 11094 139346
rect 11262 139144 12382 139346
rect 12550 139144 13670 139346
rect 13838 139144 14958 139346
rect 15126 139144 16246 139346
rect 16414 139144 17534 139346
rect 17702 139144 18822 139346
rect 18990 139144 20110 139346
rect 20278 139144 21398 139346
rect 21566 139144 22686 139346
rect 22854 139144 23974 139346
rect 24142 139144 25262 139346
rect 25430 139144 26550 139346
rect 26718 139144 27838 139346
rect 28006 139144 29126 139346
rect 29294 139144 30414 139346
rect 30582 139144 31702 139346
rect 31870 139144 32990 139346
rect 33158 139144 34278 139346
rect 34446 139144 35566 139346
rect 35734 139144 36854 139346
rect 37022 139144 38142 139346
rect 38310 139144 39430 139346
rect 39598 139144 40718 139346
rect 40886 139144 42006 139346
rect 42174 139144 43294 139346
rect 43462 139144 44582 139346
rect 44750 139144 45870 139346
rect 46038 139144 47158 139346
rect 47326 139144 48446 139346
rect 48614 139144 49734 139346
rect 49902 139144 51022 139346
rect 51190 139144 52310 139346
rect 52478 139144 53598 139346
rect 53766 139144 54886 139346
rect 55054 139144 56174 139346
rect 56342 139144 57462 139346
rect 57630 139144 58750 139346
rect 58918 139144 60038 139346
rect 60206 139144 61326 139346
rect 61494 139144 62614 139346
rect 62782 139144 63902 139346
rect 64070 139144 65190 139346
rect 65358 139144 66478 139346
rect 66646 139144 67766 139346
rect 67934 139144 69054 139346
rect 69222 139144 70342 139346
rect 70510 139144 71630 139346
rect 71798 139144 72918 139346
rect 73086 139144 74206 139346
rect 74374 139144 75494 139346
rect 75662 139144 76782 139346
rect 76950 139144 78070 139346
rect 78238 139144 79358 139346
rect 79526 139144 80646 139346
rect 80814 139144 81934 139346
rect 82102 139144 83222 139346
rect 83390 139144 84510 139346
rect 84678 139144 85798 139346
rect 85966 139144 87086 139346
rect 87254 139144 88374 139346
rect 88542 139144 89662 139346
rect 89830 139144 90950 139346
rect 91118 139144 92238 139346
rect 92406 139144 93526 139346
rect 93694 139144 94814 139346
rect 94982 139144 96102 139346
rect 96270 139144 97390 139346
rect 97558 139144 98678 139346
rect 98846 139144 99966 139346
rect 100134 139144 101254 139346
rect 101422 139144 102542 139346
rect 102710 139144 103830 139346
rect 103998 139144 105118 139346
rect 105286 139144 106406 139346
rect 106574 139144 107694 139346
rect 107862 139144 108982 139346
rect 109150 139144 110270 139346
rect 110438 139144 111558 139346
rect 111726 139144 112846 139346
rect 113014 139144 114134 139346
rect 114302 139144 115422 139346
rect 115590 139144 116710 139346
rect 116878 139144 117998 139346
rect 118166 139144 119286 139346
rect 119454 139144 120574 139346
rect 120742 139144 121862 139346
rect 122030 139144 123150 139346
rect 123318 139144 124438 139346
rect 124606 139144 125726 139346
rect 125894 139144 127014 139346
rect 127182 139144 128302 139346
rect 128470 139144 129590 139346
rect 129758 139144 130878 139346
rect 131046 139144 132166 139346
rect 132334 139144 133454 139346
rect 133622 139144 134742 139346
rect 134910 139144 136030 139346
rect 136198 139144 137318 139346
rect 137486 139144 138606 139346
rect 138774 139144 139894 139346
rect 140062 139144 141182 139346
rect 141350 139144 142470 139346
rect 142638 139144 143758 139346
rect 143926 139144 145046 139346
rect 145214 139144 146334 139346
rect 146502 139144 147622 139346
rect 147790 139144 148378 139346
rect 478 856 148378 139144
rect 478 2 1986 856
rect 2154 2 2998 856
rect 3166 2 4010 856
rect 4178 2 5022 856
rect 5190 2 6034 856
rect 6202 2 7046 856
rect 7214 2 8058 856
rect 8226 2 9070 856
rect 9238 2 10082 856
rect 10250 2 11094 856
rect 11262 2 12106 856
rect 12274 2 13118 856
rect 13286 2 14130 856
rect 14298 2 15142 856
rect 15310 2 16154 856
rect 16322 2 17166 856
rect 17334 2 18178 856
rect 18346 2 19190 856
rect 19358 2 20202 856
rect 20370 2 21214 856
rect 21382 2 22226 856
rect 22394 2 23238 856
rect 23406 2 24250 856
rect 24418 2 25262 856
rect 25430 2 26274 856
rect 26442 2 27286 856
rect 27454 2 28298 856
rect 28466 2 29310 856
rect 29478 2 30322 856
rect 30490 2 31334 856
rect 31502 2 32346 856
rect 32514 2 33358 856
rect 33526 2 34370 856
rect 34538 2 35382 856
rect 35550 2 36394 856
rect 36562 2 37406 856
rect 37574 2 38418 856
rect 38586 2 39430 856
rect 39598 2 40442 856
rect 40610 2 41454 856
rect 41622 2 42466 856
rect 42634 2 43478 856
rect 43646 2 44490 856
rect 44658 2 45502 856
rect 45670 2 46514 856
rect 46682 2 47526 856
rect 47694 2 48538 856
rect 48706 2 49550 856
rect 49718 2 50562 856
rect 50730 2 51574 856
rect 51742 2 52586 856
rect 52754 2 53598 856
rect 53766 2 54610 856
rect 54778 2 55622 856
rect 55790 2 56634 856
rect 56802 2 57646 856
rect 57814 2 58658 856
rect 58826 2 59670 856
rect 59838 2 60682 856
rect 60850 2 61694 856
rect 61862 2 62706 856
rect 62874 2 63718 856
rect 63886 2 64730 856
rect 64898 2 65742 856
rect 65910 2 66754 856
rect 66922 2 67766 856
rect 67934 2 68778 856
rect 68946 2 69790 856
rect 69958 2 70802 856
rect 70970 2 71814 856
rect 71982 2 72826 856
rect 72994 2 73838 856
rect 74006 2 74850 856
rect 75018 2 75862 856
rect 76030 2 76874 856
rect 77042 2 77886 856
rect 78054 2 78898 856
rect 79066 2 79910 856
rect 80078 2 80922 856
rect 81090 2 81934 856
rect 82102 2 82946 856
rect 83114 2 83958 856
rect 84126 2 84970 856
rect 85138 2 85982 856
rect 86150 2 86994 856
rect 87162 2 88006 856
rect 88174 2 89018 856
rect 89186 2 90030 856
rect 90198 2 91042 856
rect 91210 2 92054 856
rect 92222 2 93066 856
rect 93234 2 94078 856
rect 94246 2 95090 856
rect 95258 2 96102 856
rect 96270 2 97114 856
rect 97282 2 98126 856
rect 98294 2 99138 856
rect 99306 2 100150 856
rect 100318 2 101162 856
rect 101330 2 102174 856
rect 102342 2 103186 856
rect 103354 2 104198 856
rect 104366 2 105210 856
rect 105378 2 106222 856
rect 106390 2 107234 856
rect 107402 2 108246 856
rect 108414 2 109258 856
rect 109426 2 110270 856
rect 110438 2 111282 856
rect 111450 2 112294 856
rect 112462 2 113306 856
rect 113474 2 114318 856
rect 114486 2 115330 856
rect 115498 2 116342 856
rect 116510 2 117354 856
rect 117522 2 118366 856
rect 118534 2 119378 856
rect 119546 2 120390 856
rect 120558 2 121402 856
rect 121570 2 122414 856
rect 122582 2 123426 856
rect 123594 2 124438 856
rect 124606 2 125450 856
rect 125618 2 126462 856
rect 126630 2 127474 856
rect 127642 2 128486 856
rect 128654 2 129498 856
rect 129666 2 130510 856
rect 130678 2 131522 856
rect 131690 2 132534 856
rect 132702 2 133546 856
rect 133714 2 134558 856
rect 134726 2 135570 856
rect 135738 2 136582 856
rect 136750 2 137594 856
rect 137762 2 138606 856
rect 138774 2 139618 856
rect 139786 2 140630 856
rect 140798 2 141642 856
rect 141810 2 142654 856
rect 142822 2 143666 856
rect 143834 2 144678 856
rect 144846 2 145690 856
rect 145858 2 146702 856
rect 146870 2 147714 856
rect 147882 2 148378 856
<< metal3 >>
rect 0 136824 800 136944
rect 149200 135192 150000 135312
rect 0 133560 800 133680
rect 0 130296 800 130416
rect 0 127032 800 127152
rect 149200 126488 150000 126608
rect 0 123768 800 123888
rect 0 120504 800 120624
rect 149200 117784 150000 117904
rect 0 117240 800 117360
rect 0 113976 800 114096
rect 0 110712 800 110832
rect 149200 109080 150000 109200
rect 0 107448 800 107568
rect 0 104184 800 104304
rect 0 100920 800 101040
rect 149200 100376 150000 100496
rect 0 97656 800 97776
rect 0 94392 800 94512
rect 149200 91672 150000 91792
rect 0 91128 800 91248
rect 0 87864 800 87984
rect 0 84600 800 84720
rect 149200 82968 150000 83088
rect 0 81336 800 81456
rect 0 78072 800 78192
rect 0 74808 800 74928
rect 149200 74264 150000 74384
rect 0 71544 800 71664
rect 0 68280 800 68400
rect 149200 65560 150000 65680
rect 0 65016 800 65136
rect 0 61752 800 61872
rect 0 58488 800 58608
rect 149200 56856 150000 56976
rect 0 55224 800 55344
rect 0 51960 800 52080
rect 0 48696 800 48816
rect 149200 48152 150000 48272
rect 0 45432 800 45552
rect 0 42168 800 42288
rect 149200 39448 150000 39568
rect 0 38904 800 39024
rect 0 35640 800 35760
rect 0 32376 800 32496
rect 149200 30744 150000 30864
rect 0 29112 800 29232
rect 0 25848 800 25968
rect 0 22584 800 22704
rect 149200 22040 150000 22160
rect 0 19320 800 19440
rect 0 16056 800 16176
rect 149200 13336 150000 13456
rect 0 12792 800 12912
rect 0 9528 800 9648
rect 0 6264 800 6384
rect 149200 4632 150000 4752
rect 0 3000 800 3120
<< obsm3 >>
rect 473 137024 149200 137665
rect 880 136744 149200 137024
rect 473 135392 149200 136744
rect 473 135112 149120 135392
rect 473 133760 149200 135112
rect 880 133480 149200 133760
rect 473 130496 149200 133480
rect 880 130216 149200 130496
rect 473 127232 149200 130216
rect 880 126952 149200 127232
rect 473 126688 149200 126952
rect 473 126408 149120 126688
rect 473 123968 149200 126408
rect 880 123688 149200 123968
rect 473 120704 149200 123688
rect 880 120424 149200 120704
rect 473 117984 149200 120424
rect 473 117704 149120 117984
rect 473 117440 149200 117704
rect 880 117160 149200 117440
rect 473 114176 149200 117160
rect 880 113896 149200 114176
rect 473 110912 149200 113896
rect 880 110632 149200 110912
rect 473 109280 149200 110632
rect 473 109000 149120 109280
rect 473 107648 149200 109000
rect 880 107368 149200 107648
rect 473 104384 149200 107368
rect 880 104104 149200 104384
rect 473 101120 149200 104104
rect 880 100840 149200 101120
rect 473 100576 149200 100840
rect 473 100296 149120 100576
rect 473 97856 149200 100296
rect 880 97576 149200 97856
rect 473 94592 149200 97576
rect 880 94312 149200 94592
rect 473 91872 149200 94312
rect 473 91592 149120 91872
rect 473 91328 149200 91592
rect 880 91048 149200 91328
rect 473 88064 149200 91048
rect 880 87784 149200 88064
rect 473 84800 149200 87784
rect 880 84520 149200 84800
rect 473 83168 149200 84520
rect 473 82888 149120 83168
rect 473 81536 149200 82888
rect 880 81256 149200 81536
rect 473 78272 149200 81256
rect 880 77992 149200 78272
rect 473 75008 149200 77992
rect 880 74728 149200 75008
rect 473 74464 149200 74728
rect 473 74184 149120 74464
rect 473 71744 149200 74184
rect 880 71464 149200 71744
rect 473 68480 149200 71464
rect 880 68200 149200 68480
rect 473 65760 149200 68200
rect 473 65480 149120 65760
rect 473 65216 149200 65480
rect 880 64936 149200 65216
rect 473 61952 149200 64936
rect 880 61672 149200 61952
rect 473 58688 149200 61672
rect 880 58408 149200 58688
rect 473 57056 149200 58408
rect 473 56776 149120 57056
rect 473 55424 149200 56776
rect 880 55144 149200 55424
rect 473 52160 149200 55144
rect 880 51880 149200 52160
rect 473 48896 149200 51880
rect 880 48616 149200 48896
rect 473 48352 149200 48616
rect 473 48072 149120 48352
rect 473 45632 149200 48072
rect 880 45352 149200 45632
rect 473 42368 149200 45352
rect 880 42088 149200 42368
rect 473 39648 149200 42088
rect 473 39368 149120 39648
rect 473 39104 149200 39368
rect 880 38824 149200 39104
rect 473 35840 149200 38824
rect 880 35560 149200 35840
rect 473 32576 149200 35560
rect 880 32296 149200 32576
rect 473 30944 149200 32296
rect 473 30664 149120 30944
rect 473 29312 149200 30664
rect 880 29032 149200 29312
rect 473 26048 149200 29032
rect 880 25768 149200 26048
rect 473 22784 149200 25768
rect 880 22504 149200 22784
rect 473 22240 149200 22504
rect 473 21960 149120 22240
rect 473 19520 149200 21960
rect 880 19240 149200 19520
rect 473 16256 149200 19240
rect 880 15976 149200 16256
rect 473 13536 149200 15976
rect 473 13256 149120 13536
rect 473 12992 149200 13256
rect 880 12712 149200 12992
rect 473 9728 149200 12712
rect 880 9448 149200 9728
rect 473 6464 149200 9448
rect 880 6184 149200 6464
rect 473 4832 149200 6184
rect 473 4552 149120 4832
rect 473 3200 149200 4552
rect 880 2920 149200 3200
rect 473 35 149200 2920
<< metal4 >>
rect 4208 2128 4528 137680
rect 19568 2128 19888 137680
rect 34928 2128 35248 137680
rect 50288 2128 50608 137680
rect 65648 2128 65968 137680
rect 81008 2128 81328 137680
rect 96368 2128 96688 137680
rect 111728 2128 112048 137680
rect 127088 2128 127408 137680
rect 142448 2128 142768 137680
<< obsm4 >>
rect 795 2048 4128 137325
rect 4608 2048 19488 137325
rect 19968 2048 34848 137325
rect 35328 2048 50208 137325
rect 50688 2048 65568 137325
rect 66048 2048 80928 137325
rect 81408 2048 96288 137325
rect 96768 2048 111648 137325
rect 112128 2048 127008 137325
rect 127488 2048 128370 137325
rect 795 715 128370 2048
<< labels >>
rlabel metal2 s 2134 139200 2190 140000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 40774 139200 40830 140000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 44638 139200 44694 140000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 48502 139200 48558 140000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 52366 139200 52422 140000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 56230 139200 56286 140000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 60094 139200 60150 140000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 63958 139200 64014 140000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 67822 139200 67878 140000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 71686 139200 71742 140000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 75550 139200 75606 140000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 5998 139200 6054 140000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 79414 139200 79470 140000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 83278 139200 83334 140000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 87142 139200 87198 140000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 91006 139200 91062 140000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 94870 139200 94926 140000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 98734 139200 98790 140000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 102598 139200 102654 140000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 106462 139200 106518 140000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 110326 139200 110382 140000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 114190 139200 114246 140000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 9862 139200 9918 140000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 118054 139200 118110 140000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 121918 139200 121974 140000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 125782 139200 125838 140000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 129646 139200 129702 140000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 133510 139200 133566 140000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 137374 139200 137430 140000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 141238 139200 141294 140000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 145102 139200 145158 140000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 13726 139200 13782 140000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 17590 139200 17646 140000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 21454 139200 21510 140000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 25318 139200 25374 140000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 29182 139200 29238 140000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 33046 139200 33102 140000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 36910 139200 36966 140000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 3422 139200 3478 140000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 42062 139200 42118 140000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 45926 139200 45982 140000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 49790 139200 49846 140000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 53654 139200 53710 140000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 57518 139200 57574 140000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 61382 139200 61438 140000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 65246 139200 65302 140000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 69110 139200 69166 140000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 72974 139200 73030 140000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 76838 139200 76894 140000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 7286 139200 7342 140000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 80702 139200 80758 140000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 84566 139200 84622 140000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 88430 139200 88486 140000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 92294 139200 92350 140000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 96158 139200 96214 140000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 100022 139200 100078 140000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 103886 139200 103942 140000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 107750 139200 107806 140000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 111614 139200 111670 140000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 115478 139200 115534 140000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 11150 139200 11206 140000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 119342 139200 119398 140000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 123206 139200 123262 140000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 127070 139200 127126 140000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 130934 139200 130990 140000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 134798 139200 134854 140000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 138662 139200 138718 140000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 142526 139200 142582 140000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 146390 139200 146446 140000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 15014 139200 15070 140000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 18878 139200 18934 140000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 22742 139200 22798 140000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 26606 139200 26662 140000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 30470 139200 30526 140000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 34334 139200 34390 140000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 38198 139200 38254 140000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 4710 139200 4766 140000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 43350 139200 43406 140000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 47214 139200 47270 140000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 51078 139200 51134 140000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 54942 139200 54998 140000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 58806 139200 58862 140000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 62670 139200 62726 140000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 66534 139200 66590 140000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 70398 139200 70454 140000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 74262 139200 74318 140000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 78126 139200 78182 140000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 8574 139200 8630 140000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 81990 139200 82046 140000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 85854 139200 85910 140000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 89718 139200 89774 140000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 93582 139200 93638 140000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 97446 139200 97502 140000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 101310 139200 101366 140000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 105174 139200 105230 140000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 109038 139200 109094 140000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 112902 139200 112958 140000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 116766 139200 116822 140000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 12438 139200 12494 140000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 120630 139200 120686 140000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 124494 139200 124550 140000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 128358 139200 128414 140000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 132222 139200 132278 140000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 136086 139200 136142 140000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 139950 139200 140006 140000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 143814 139200 143870 140000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 147678 139200 147734 140000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 16302 139200 16358 140000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 20166 139200 20222 140000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 24030 139200 24086 140000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 27894 139200 27950 140000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 31758 139200 31814 140000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 35622 139200 35678 140000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 39486 139200 39542 140000 6 io_out[9]
port 114 nsew signal output
rlabel metal3 s 149200 13336 150000 13456 6 ram_addr[0]
port 115 nsew signal output
rlabel metal3 s 149200 39448 150000 39568 6 ram_addr[1]
port 116 nsew signal output
rlabel metal3 s 149200 65560 150000 65680 6 ram_addr[2]
port 117 nsew signal output
rlabel metal3 s 149200 91672 150000 91792 6 ram_addr[3]
port 118 nsew signal output
rlabel metal3 s 149200 117784 150000 117904 6 ram_addr[4]
port 119 nsew signal output
rlabel metal3 s 149200 126488 150000 126608 6 ram_addr[5]
port 120 nsew signal output
rlabel metal3 s 149200 135192 150000 135312 6 ram_addr[6]
port 121 nsew signal output
rlabel metal3 s 149200 22040 150000 22160 6 ram_val_in[0]
port 122 nsew signal input
rlabel metal3 s 149200 48152 150000 48272 6 ram_val_in[1]
port 123 nsew signal input
rlabel metal3 s 149200 74264 150000 74384 6 ram_val_in[2]
port 124 nsew signal input
rlabel metal3 s 149200 100376 150000 100496 6 ram_val_in[3]
port 125 nsew signal input
rlabel metal3 s 149200 30744 150000 30864 6 ram_val_out[0]
port 126 nsew signal output
rlabel metal3 s 149200 56856 150000 56976 6 ram_val_out[1]
port 127 nsew signal output
rlabel metal3 s 149200 82968 150000 83088 6 ram_val_out[2]
port 128 nsew signal output
rlabel metal3 s 149200 109080 150000 109200 6 ram_val_out[3]
port 129 nsew signal output
rlabel metal3 s 149200 4632 150000 4752 6 ram_we
port 130 nsew signal output
rlabel metal3 s 0 6264 800 6384 6 rom_addr[0]
port 131 nsew signal output
rlabel metal3 s 0 12792 800 12912 6 rom_addr[1]
port 132 nsew signal output
rlabel metal3 s 0 19320 800 19440 6 rom_addr[2]
port 133 nsew signal output
rlabel metal3 s 0 25848 800 25968 6 rom_addr[3]
port 134 nsew signal output
rlabel metal3 s 0 32376 800 32496 6 rom_addr[4]
port 135 nsew signal output
rlabel metal3 s 0 38904 800 39024 6 rom_addr[5]
port 136 nsew signal output
rlabel metal3 s 0 45432 800 45552 6 rom_addr[6]
port 137 nsew signal output
rlabel metal3 s 0 51960 800 52080 6 rom_addr[7]
port 138 nsew signal output
rlabel metal3 s 0 58488 800 58608 6 rom_addr[8]
port 139 nsew signal output
rlabel metal3 s 0 3000 800 3120 6 rom_csb
port 140 nsew signal output
rlabel metal3 s 0 9528 800 9648 6 rom_value[0]
port 141 nsew signal input
rlabel metal3 s 0 68280 800 68400 6 rom_value[10]
port 142 nsew signal input
rlabel metal3 s 0 71544 800 71664 6 rom_value[11]
port 143 nsew signal input
rlabel metal3 s 0 74808 800 74928 6 rom_value[12]
port 144 nsew signal input
rlabel metal3 s 0 78072 800 78192 6 rom_value[13]
port 145 nsew signal input
rlabel metal3 s 0 81336 800 81456 6 rom_value[14]
port 146 nsew signal input
rlabel metal3 s 0 84600 800 84720 6 rom_value[15]
port 147 nsew signal input
rlabel metal3 s 0 87864 800 87984 6 rom_value[16]
port 148 nsew signal input
rlabel metal3 s 0 91128 800 91248 6 rom_value[17]
port 149 nsew signal input
rlabel metal3 s 0 94392 800 94512 6 rom_value[18]
port 150 nsew signal input
rlabel metal3 s 0 97656 800 97776 6 rom_value[19]
port 151 nsew signal input
rlabel metal3 s 0 16056 800 16176 6 rom_value[1]
port 152 nsew signal input
rlabel metal3 s 0 100920 800 101040 6 rom_value[20]
port 153 nsew signal input
rlabel metal3 s 0 104184 800 104304 6 rom_value[21]
port 154 nsew signal input
rlabel metal3 s 0 107448 800 107568 6 rom_value[22]
port 155 nsew signal input
rlabel metal3 s 0 110712 800 110832 6 rom_value[23]
port 156 nsew signal input
rlabel metal3 s 0 113976 800 114096 6 rom_value[24]
port 157 nsew signal input
rlabel metal3 s 0 117240 800 117360 6 rom_value[25]
port 158 nsew signal input
rlabel metal3 s 0 120504 800 120624 6 rom_value[26]
port 159 nsew signal input
rlabel metal3 s 0 123768 800 123888 6 rom_value[27]
port 160 nsew signal input
rlabel metal3 s 0 127032 800 127152 6 rom_value[28]
port 161 nsew signal input
rlabel metal3 s 0 130296 800 130416 6 rom_value[29]
port 162 nsew signal input
rlabel metal3 s 0 22584 800 22704 6 rom_value[2]
port 163 nsew signal input
rlabel metal3 s 0 133560 800 133680 6 rom_value[30]
port 164 nsew signal input
rlabel metal3 s 0 136824 800 136944 6 rom_value[31]
port 165 nsew signal input
rlabel metal3 s 0 29112 800 29232 6 rom_value[3]
port 166 nsew signal input
rlabel metal3 s 0 35640 800 35760 6 rom_value[4]
port 167 nsew signal input
rlabel metal3 s 0 42168 800 42288 6 rom_value[5]
port 168 nsew signal input
rlabel metal3 s 0 48696 800 48816 6 rom_value[6]
port 169 nsew signal input
rlabel metal3 s 0 55224 800 55344 6 rom_value[7]
port 170 nsew signal input
rlabel metal3 s 0 61752 800 61872 6 rom_value[8]
port 171 nsew signal input
rlabel metal3 s 0 65016 800 65136 6 rom_value[9]
port 172 nsew signal input
rlabel metal4 s 4208 2128 4528 137680 6 vccd1
port 173 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 137680 6 vccd1
port 173 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 137680 6 vccd1
port 173 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 137680 6 vccd1
port 173 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 137680 6 vccd1
port 173 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 137680 6 vssd1
port 174 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 137680 6 vssd1
port 174 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 137680 6 vssd1
port 174 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 137680 6 vssd1
port 174 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 137680 6 vssd1
port 174 nsew ground bidirectional
rlabel metal2 s 2042 0 2098 800 6 wb_clk_i
port 175 nsew signal input
rlabel metal2 s 6090 0 6146 800 6 wb_rom_adrb[0]
port 176 nsew signal output
rlabel metal2 s 8114 0 8170 800 6 wb_rom_adrb[1]
port 177 nsew signal output
rlabel metal2 s 10138 0 10194 800 6 wb_rom_adrb[2]
port 178 nsew signal output
rlabel metal2 s 12162 0 12218 800 6 wb_rom_adrb[3]
port 179 nsew signal output
rlabel metal2 s 14186 0 14242 800 6 wb_rom_adrb[4]
port 180 nsew signal output
rlabel metal2 s 16210 0 16266 800 6 wb_rom_adrb[5]
port 181 nsew signal output
rlabel metal2 s 18234 0 18290 800 6 wb_rom_adrb[6]
port 182 nsew signal output
rlabel metal2 s 20258 0 20314 800 6 wb_rom_adrb[7]
port 183 nsew signal output
rlabel metal2 s 22282 0 22338 800 6 wb_rom_adrb[8]
port 184 nsew signal output
rlabel metal2 s 3054 0 3110 800 6 wb_rom_csb
port 185 nsew signal output
rlabel metal2 s 7102 0 7158 800 6 wb_rom_val[0]
port 186 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 wb_rom_val[10]
port 187 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 wb_rom_val[11]
port 188 nsew signal input
rlabel metal2 s 27342 0 27398 800 6 wb_rom_val[12]
port 189 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 wb_rom_val[13]
port 190 nsew signal input
rlabel metal2 s 29366 0 29422 800 6 wb_rom_val[14]
port 191 nsew signal input
rlabel metal2 s 30378 0 30434 800 6 wb_rom_val[15]
port 192 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 wb_rom_val[16]
port 193 nsew signal input
rlabel metal2 s 32402 0 32458 800 6 wb_rom_val[17]
port 194 nsew signal input
rlabel metal2 s 33414 0 33470 800 6 wb_rom_val[18]
port 195 nsew signal input
rlabel metal2 s 34426 0 34482 800 6 wb_rom_val[19]
port 196 nsew signal input
rlabel metal2 s 9126 0 9182 800 6 wb_rom_val[1]
port 197 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 wb_rom_val[20]
port 198 nsew signal input
rlabel metal2 s 36450 0 36506 800 6 wb_rom_val[21]
port 199 nsew signal input
rlabel metal2 s 37462 0 37518 800 6 wb_rom_val[22]
port 200 nsew signal input
rlabel metal2 s 38474 0 38530 800 6 wb_rom_val[23]
port 201 nsew signal input
rlabel metal2 s 39486 0 39542 800 6 wb_rom_val[24]
port 202 nsew signal input
rlabel metal2 s 40498 0 40554 800 6 wb_rom_val[25]
port 203 nsew signal input
rlabel metal2 s 41510 0 41566 800 6 wb_rom_val[26]
port 204 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 wb_rom_val[27]
port 205 nsew signal input
rlabel metal2 s 43534 0 43590 800 6 wb_rom_val[28]
port 206 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 wb_rom_val[29]
port 207 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 wb_rom_val[2]
port 208 nsew signal input
rlabel metal2 s 45558 0 45614 800 6 wb_rom_val[30]
port 209 nsew signal input
rlabel metal2 s 46570 0 46626 800 6 wb_rom_val[31]
port 210 nsew signal input
rlabel metal2 s 13174 0 13230 800 6 wb_rom_val[3]
port 211 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 wb_rom_val[4]
port 212 nsew signal input
rlabel metal2 s 17222 0 17278 800 6 wb_rom_val[5]
port 213 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 wb_rom_val[6]
port 214 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 wb_rom_val[7]
port 215 nsew signal input
rlabel metal2 s 23294 0 23350 800 6 wb_rom_val[8]
port 216 nsew signal input
rlabel metal2 s 24306 0 24362 800 6 wb_rom_val[9]
port 217 nsew signal input
rlabel metal2 s 4066 0 4122 800 6 wb_rom_web
port 218 nsew signal output
rlabel metal2 s 5078 0 5134 800 6 wb_rst_i
port 219 nsew signal input
rlabel metal2 s 47582 0 47638 800 6 wbs_ack_o
port 220 nsew signal output
rlabel metal2 s 51630 0 51686 800 6 wbs_adr_i[0]
port 221 nsew signal input
rlabel metal2 s 81990 0 82046 800 6 wbs_adr_i[10]
port 222 nsew signal input
rlabel metal2 s 85026 0 85082 800 6 wbs_adr_i[11]
port 223 nsew signal input
rlabel metal2 s 88062 0 88118 800 6 wbs_adr_i[12]
port 224 nsew signal input
rlabel metal2 s 91098 0 91154 800 6 wbs_adr_i[13]
port 225 nsew signal input
rlabel metal2 s 94134 0 94190 800 6 wbs_adr_i[14]
port 226 nsew signal input
rlabel metal2 s 97170 0 97226 800 6 wbs_adr_i[15]
port 227 nsew signal input
rlabel metal2 s 100206 0 100262 800 6 wbs_adr_i[16]
port 228 nsew signal input
rlabel metal2 s 103242 0 103298 800 6 wbs_adr_i[17]
port 229 nsew signal input
rlabel metal2 s 106278 0 106334 800 6 wbs_adr_i[18]
port 230 nsew signal input
rlabel metal2 s 109314 0 109370 800 6 wbs_adr_i[19]
port 231 nsew signal input
rlabel metal2 s 54666 0 54722 800 6 wbs_adr_i[1]
port 232 nsew signal input
rlabel metal2 s 112350 0 112406 800 6 wbs_adr_i[20]
port 233 nsew signal input
rlabel metal2 s 115386 0 115442 800 6 wbs_adr_i[21]
port 234 nsew signal input
rlabel metal2 s 118422 0 118478 800 6 wbs_adr_i[22]
port 235 nsew signal input
rlabel metal2 s 121458 0 121514 800 6 wbs_adr_i[23]
port 236 nsew signal input
rlabel metal2 s 124494 0 124550 800 6 wbs_adr_i[24]
port 237 nsew signal input
rlabel metal2 s 127530 0 127586 800 6 wbs_adr_i[25]
port 238 nsew signal input
rlabel metal2 s 130566 0 130622 800 6 wbs_adr_i[26]
port 239 nsew signal input
rlabel metal2 s 133602 0 133658 800 6 wbs_adr_i[27]
port 240 nsew signal input
rlabel metal2 s 136638 0 136694 800 6 wbs_adr_i[28]
port 241 nsew signal input
rlabel metal2 s 139674 0 139730 800 6 wbs_adr_i[29]
port 242 nsew signal input
rlabel metal2 s 57702 0 57758 800 6 wbs_adr_i[2]
port 243 nsew signal input
rlabel metal2 s 142710 0 142766 800 6 wbs_adr_i[30]
port 244 nsew signal input
rlabel metal2 s 145746 0 145802 800 6 wbs_adr_i[31]
port 245 nsew signal input
rlabel metal2 s 60738 0 60794 800 6 wbs_adr_i[3]
port 246 nsew signal input
rlabel metal2 s 63774 0 63830 800 6 wbs_adr_i[4]
port 247 nsew signal input
rlabel metal2 s 66810 0 66866 800 6 wbs_adr_i[5]
port 248 nsew signal input
rlabel metal2 s 69846 0 69902 800 6 wbs_adr_i[6]
port 249 nsew signal input
rlabel metal2 s 72882 0 72938 800 6 wbs_adr_i[7]
port 250 nsew signal input
rlabel metal2 s 75918 0 75974 800 6 wbs_adr_i[8]
port 251 nsew signal input
rlabel metal2 s 78954 0 79010 800 6 wbs_adr_i[9]
port 252 nsew signal input
rlabel metal2 s 48594 0 48650 800 6 wbs_cyc_i
port 253 nsew signal input
rlabel metal2 s 52642 0 52698 800 6 wbs_dat_i[0]
port 254 nsew signal input
rlabel metal2 s 83002 0 83058 800 6 wbs_dat_i[10]
port 255 nsew signal input
rlabel metal2 s 86038 0 86094 800 6 wbs_dat_i[11]
port 256 nsew signal input
rlabel metal2 s 89074 0 89130 800 6 wbs_dat_i[12]
port 257 nsew signal input
rlabel metal2 s 92110 0 92166 800 6 wbs_dat_i[13]
port 258 nsew signal input
rlabel metal2 s 95146 0 95202 800 6 wbs_dat_i[14]
port 259 nsew signal input
rlabel metal2 s 98182 0 98238 800 6 wbs_dat_i[15]
port 260 nsew signal input
rlabel metal2 s 101218 0 101274 800 6 wbs_dat_i[16]
port 261 nsew signal input
rlabel metal2 s 104254 0 104310 800 6 wbs_dat_i[17]
port 262 nsew signal input
rlabel metal2 s 107290 0 107346 800 6 wbs_dat_i[18]
port 263 nsew signal input
rlabel metal2 s 110326 0 110382 800 6 wbs_dat_i[19]
port 264 nsew signal input
rlabel metal2 s 55678 0 55734 800 6 wbs_dat_i[1]
port 265 nsew signal input
rlabel metal2 s 113362 0 113418 800 6 wbs_dat_i[20]
port 266 nsew signal input
rlabel metal2 s 116398 0 116454 800 6 wbs_dat_i[21]
port 267 nsew signal input
rlabel metal2 s 119434 0 119490 800 6 wbs_dat_i[22]
port 268 nsew signal input
rlabel metal2 s 122470 0 122526 800 6 wbs_dat_i[23]
port 269 nsew signal input
rlabel metal2 s 125506 0 125562 800 6 wbs_dat_i[24]
port 270 nsew signal input
rlabel metal2 s 128542 0 128598 800 6 wbs_dat_i[25]
port 271 nsew signal input
rlabel metal2 s 131578 0 131634 800 6 wbs_dat_i[26]
port 272 nsew signal input
rlabel metal2 s 134614 0 134670 800 6 wbs_dat_i[27]
port 273 nsew signal input
rlabel metal2 s 137650 0 137706 800 6 wbs_dat_i[28]
port 274 nsew signal input
rlabel metal2 s 140686 0 140742 800 6 wbs_dat_i[29]
port 275 nsew signal input
rlabel metal2 s 58714 0 58770 800 6 wbs_dat_i[2]
port 276 nsew signal input
rlabel metal2 s 143722 0 143778 800 6 wbs_dat_i[30]
port 277 nsew signal input
rlabel metal2 s 146758 0 146814 800 6 wbs_dat_i[31]
port 278 nsew signal input
rlabel metal2 s 61750 0 61806 800 6 wbs_dat_i[3]
port 279 nsew signal input
rlabel metal2 s 64786 0 64842 800 6 wbs_dat_i[4]
port 280 nsew signal input
rlabel metal2 s 67822 0 67878 800 6 wbs_dat_i[5]
port 281 nsew signal input
rlabel metal2 s 70858 0 70914 800 6 wbs_dat_i[6]
port 282 nsew signal input
rlabel metal2 s 73894 0 73950 800 6 wbs_dat_i[7]
port 283 nsew signal input
rlabel metal2 s 76930 0 76986 800 6 wbs_dat_i[8]
port 284 nsew signal input
rlabel metal2 s 79966 0 80022 800 6 wbs_dat_i[9]
port 285 nsew signal input
rlabel metal2 s 53654 0 53710 800 6 wbs_dat_o[0]
port 286 nsew signal output
rlabel metal2 s 84014 0 84070 800 6 wbs_dat_o[10]
port 287 nsew signal output
rlabel metal2 s 87050 0 87106 800 6 wbs_dat_o[11]
port 288 nsew signal output
rlabel metal2 s 90086 0 90142 800 6 wbs_dat_o[12]
port 289 nsew signal output
rlabel metal2 s 93122 0 93178 800 6 wbs_dat_o[13]
port 290 nsew signal output
rlabel metal2 s 96158 0 96214 800 6 wbs_dat_o[14]
port 291 nsew signal output
rlabel metal2 s 99194 0 99250 800 6 wbs_dat_o[15]
port 292 nsew signal output
rlabel metal2 s 102230 0 102286 800 6 wbs_dat_o[16]
port 293 nsew signal output
rlabel metal2 s 105266 0 105322 800 6 wbs_dat_o[17]
port 294 nsew signal output
rlabel metal2 s 108302 0 108358 800 6 wbs_dat_o[18]
port 295 nsew signal output
rlabel metal2 s 111338 0 111394 800 6 wbs_dat_o[19]
port 296 nsew signal output
rlabel metal2 s 56690 0 56746 800 6 wbs_dat_o[1]
port 297 nsew signal output
rlabel metal2 s 114374 0 114430 800 6 wbs_dat_o[20]
port 298 nsew signal output
rlabel metal2 s 117410 0 117466 800 6 wbs_dat_o[21]
port 299 nsew signal output
rlabel metal2 s 120446 0 120502 800 6 wbs_dat_o[22]
port 300 nsew signal output
rlabel metal2 s 123482 0 123538 800 6 wbs_dat_o[23]
port 301 nsew signal output
rlabel metal2 s 126518 0 126574 800 6 wbs_dat_o[24]
port 302 nsew signal output
rlabel metal2 s 129554 0 129610 800 6 wbs_dat_o[25]
port 303 nsew signal output
rlabel metal2 s 132590 0 132646 800 6 wbs_dat_o[26]
port 304 nsew signal output
rlabel metal2 s 135626 0 135682 800 6 wbs_dat_o[27]
port 305 nsew signal output
rlabel metal2 s 138662 0 138718 800 6 wbs_dat_o[28]
port 306 nsew signal output
rlabel metal2 s 141698 0 141754 800 6 wbs_dat_o[29]
port 307 nsew signal output
rlabel metal2 s 59726 0 59782 800 6 wbs_dat_o[2]
port 308 nsew signal output
rlabel metal2 s 144734 0 144790 800 6 wbs_dat_o[30]
port 309 nsew signal output
rlabel metal2 s 147770 0 147826 800 6 wbs_dat_o[31]
port 310 nsew signal output
rlabel metal2 s 62762 0 62818 800 6 wbs_dat_o[3]
port 311 nsew signal output
rlabel metal2 s 65798 0 65854 800 6 wbs_dat_o[4]
port 312 nsew signal output
rlabel metal2 s 68834 0 68890 800 6 wbs_dat_o[5]
port 313 nsew signal output
rlabel metal2 s 71870 0 71926 800 6 wbs_dat_o[6]
port 314 nsew signal output
rlabel metal2 s 74906 0 74962 800 6 wbs_dat_o[7]
port 315 nsew signal output
rlabel metal2 s 77942 0 77998 800 6 wbs_dat_o[8]
port 316 nsew signal output
rlabel metal2 s 80978 0 81034 800 6 wbs_dat_o[9]
port 317 nsew signal output
rlabel metal2 s 49606 0 49662 800 6 wbs_stb_i
port 318 nsew signal input
rlabel metal2 s 50618 0 50674 800 6 wbs_we_i
port 319 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 150000 140000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 47901890
string GDS_FILE /home/lucah/Videos/mpw-8-as1x00/openlane/wrapped_tms1x00/runs/23_01_19_17_45/results/signoff/wrapped_tms1x00.magic.gds
string GDS_START 790528
<< end >>

