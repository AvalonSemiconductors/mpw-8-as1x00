magic
tech sky130B
magscale 1 2
timestamp 1674061931
<< obsli1 >>
rect 1104 2159 50048 48977
<< obsm1 >>
rect 1104 1980 50048 49292
<< metal2 >>
rect 12714 50400 12770 51200
rect 38290 50400 38346 51200
<< obsm2 >>
rect 1400 50344 12658 50538
rect 12826 50344 38234 50538
rect 38402 50344 49476 50538
rect 1400 1663 49476 50344
<< metal3 >>
rect 0 49240 800 49360
rect 0 45840 800 45960
rect 0 42440 800 42560
rect 0 39040 800 39160
rect 0 35640 800 35760
rect 0 32240 800 32360
rect 0 28840 800 28960
rect 0 25440 800 25560
rect 0 22040 800 22160
rect 0 18640 800 18760
rect 0 15240 800 15360
rect 0 11840 800 11960
rect 0 8440 800 8560
rect 0 5040 800 5160
rect 0 1640 800 1760
<< obsm3 >>
rect 880 49160 49115 49333
rect 800 46040 49115 49160
rect 880 45760 49115 46040
rect 800 42640 49115 45760
rect 880 42360 49115 42640
rect 800 39240 49115 42360
rect 880 38960 49115 39240
rect 800 35840 49115 38960
rect 880 35560 49115 35840
rect 800 32440 49115 35560
rect 880 32160 49115 32440
rect 800 29040 49115 32160
rect 880 28760 49115 29040
rect 800 25640 49115 28760
rect 880 25360 49115 25640
rect 800 22240 49115 25360
rect 880 21960 49115 22240
rect 800 18840 49115 21960
rect 880 18560 49115 18840
rect 800 15440 49115 18560
rect 880 15160 49115 15440
rect 800 12040 49115 15160
rect 880 11760 49115 12040
rect 800 8640 49115 11760
rect 880 8360 49115 8640
rect 800 5240 49115 8360
rect 880 4960 49115 5240
rect 800 1840 49115 4960
rect 880 1667 49115 1840
<< metal4 >>
rect 4208 2128 4528 49008
rect 19568 2128 19888 49008
rect 34928 2128 35248 49008
<< obsm4 >>
rect 4843 2483 19488 48653
rect 19968 2483 34848 48653
rect 35328 2483 45389 48653
<< labels >>
rlabel metal2 s 38290 50400 38346 51200 6 clk
port 1 nsew signal input
rlabel metal3 s 0 39040 800 39160 6 r_val[0]
port 2 nsew signal output
rlabel metal3 s 0 42440 800 42560 6 r_val[1]
port 3 nsew signal output
rlabel metal3 s 0 45840 800 45960 6 r_val[2]
port 4 nsew signal output
rlabel metal3 s 0 49240 800 49360 6 r_val[3]
port 5 nsew signal output
rlabel metal3 s 0 1640 800 1760 6 ram_addr[0]
port 6 nsew signal input
rlabel metal3 s 0 5040 800 5160 6 ram_addr[1]
port 7 nsew signal input
rlabel metal3 s 0 8440 800 8560 6 ram_addr[2]
port 8 nsew signal input
rlabel metal3 s 0 11840 800 11960 6 ram_addr[3]
port 9 nsew signal input
rlabel metal3 s 0 15240 800 15360 6 ram_addr[4]
port 10 nsew signal input
rlabel metal3 s 0 18640 800 18760 6 ram_addr[5]
port 11 nsew signal input
rlabel metal3 s 0 22040 800 22160 6 ram_addr[6]
port 12 nsew signal input
rlabel metal4 s 4208 2128 4528 49008 6 vccd1
port 13 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 49008 6 vccd1
port 13 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 49008 6 vssd1
port 14 nsew ground bidirectional
rlabel metal3 s 0 25440 800 25560 6 w_val[0]
port 15 nsew signal input
rlabel metal3 s 0 28840 800 28960 6 w_val[1]
port 16 nsew signal input
rlabel metal3 s 0 32240 800 32360 6 w_val[2]
port 17 nsew signal input
rlabel metal3 s 0 35640 800 35760 6 w_val[3]
port 18 nsew signal input
rlabel metal2 s 12714 50400 12770 51200 6 wen
port 19 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 51200 51200
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 7964888
string GDS_FILE /home/lucah/Videos/mpw-8-as1x00/openlane/tms1x00_ram/runs/23_01_18_18_08/results/signoff/tms1x00_ram.magic.gds
string GDS_START 389350
<< end >>

