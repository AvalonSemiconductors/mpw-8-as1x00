VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_tms1x00
  CLASS BLOCK ;
  FOREIGN wrapped_tms1x00 ;
  ORIGIN 0.000 0.000 ;
  SIZE 650.000 BY 450.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 446.000 13.250 450.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.570 446.000 178.850 450.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.130 446.000 195.410 450.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.690 446.000 211.970 450.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.250 446.000 228.530 450.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 446.000 245.090 450.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.370 446.000 261.650 450.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.930 446.000 278.210 450.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.490 446.000 294.770 450.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.050 446.000 311.330 450.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.610 446.000 327.890 450.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 446.000 29.810 450.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.170 446.000 344.450 450.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 446.000 361.010 450.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.290 446.000 377.570 450.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.850 446.000 394.130 450.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.410 446.000 410.690 450.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.970 446.000 427.250 450.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.530 446.000 443.810 450.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.090 446.000 460.370 450.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.650 446.000 476.930 450.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.210 446.000 493.490 450.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 446.000 46.370 450.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.770 446.000 510.050 450.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.330 446.000 526.610 450.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.890 446.000 543.170 450.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.450 446.000 559.730 450.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.010 446.000 576.290 450.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.570 446.000 592.850 450.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.130 446.000 609.410 450.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 625.690 446.000 625.970 450.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 446.000 62.930 450.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 446.000 79.490 450.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 446.000 96.050 450.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 446.000 112.610 450.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 446.000 129.170 450.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.450 446.000 145.730 450.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 446.000 162.290 450.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 446.000 18.770 450.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 446.000 184.370 450.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.650 446.000 200.930 450.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.210 446.000 217.490 450.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 446.000 234.050 450.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.330 446.000 250.610 450.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 446.000 267.170 450.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 446.000 283.730 450.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.010 446.000 300.290 450.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.570 446.000 316.850 450.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.130 446.000 333.410 450.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 446.000 35.330 450.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.690 446.000 349.970 450.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.250 446.000 366.530 450.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.810 446.000 383.090 450.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 446.000 399.650 450.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.930 446.000 416.210 450.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.490 446.000 432.770 450.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.050 446.000 449.330 450.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.610 446.000 465.890 450.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.170 446.000 482.450 450.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.730 446.000 499.010 450.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 446.000 51.890 450.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.290 446.000 515.570 450.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.850 446.000 532.130 450.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 548.410 446.000 548.690 450.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.970 446.000 565.250 450.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.530 446.000 581.810 450.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.090 446.000 598.370 450.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.650 446.000 614.930 450.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.210 446.000 631.490 450.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 446.000 68.450 450.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 446.000 85.010 450.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 446.000 101.570 450.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 446.000 118.130 450.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.410 446.000 134.690 450.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 446.000 151.250 450.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 446.000 167.810 450.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 446.000 24.290 450.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.610 446.000 189.890 450.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 446.000 206.450 450.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.730 446.000 223.010 450.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.290 446.000 239.570 450.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.850 446.000 256.130 450.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.410 446.000 272.690 450.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.970 446.000 289.250 450.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.530 446.000 305.810 450.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 446.000 322.370 450.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.650 446.000 338.930 450.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 446.000 40.850 450.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.210 446.000 355.490 450.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.770 446.000 372.050 450.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.330 446.000 388.610 450.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.890 446.000 405.170 450.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.450 446.000 421.730 450.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 446.000 438.290 450.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.570 446.000 454.850 450.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.130 446.000 471.410 450.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.690 446.000 487.970 450.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.250 446.000 504.530 450.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 446.000 57.410 450.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.810 446.000 521.090 450.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.370 446.000 537.650 450.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 446.000 554.210 450.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.490 446.000 570.770 450.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.050 446.000 587.330 450.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.610 446.000 603.890 450.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.170 446.000 620.450 450.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 636.730 446.000 637.010 450.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 446.000 73.970 450.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 446.000 90.530 450.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 446.000 107.090 450.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 446.000 123.650 450.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.930 446.000 140.210 450.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.490 446.000 156.770 450.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.050 446.000 173.330 450.000 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.630 0.000 620.910 4.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.770 0.000 625.050 4.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.910 0.000 629.190 4.000 ;
    END
  END irq[2]
  PIN ram_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 646.000 43.560 650.000 44.160 ;
    END
  END ram_addr[0]
  PIN ram_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 646.000 127.200 650.000 127.800 ;
    END
  END ram_addr[1]
  PIN ram_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 646.000 210.840 650.000 211.440 ;
    END
  END ram_addr[2]
  PIN ram_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 646.000 294.480 650.000 295.080 ;
    END
  END ram_addr[3]
  PIN ram_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 646.000 378.120 650.000 378.720 ;
    END
  END ram_addr[4]
  PIN ram_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 646.000 406.000 650.000 406.600 ;
    END
  END ram_addr[5]
  PIN ram_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 646.000 433.880 650.000 434.480 ;
    END
  END ram_addr[6]
  PIN ram_val_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 646.000 71.440 650.000 72.040 ;
    END
  END ram_val_in[0]
  PIN ram_val_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 646.000 155.080 650.000 155.680 ;
    END
  END ram_val_in[1]
  PIN ram_val_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 646.000 238.720 650.000 239.320 ;
    END
  END ram_val_in[2]
  PIN ram_val_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 646.000 322.360 650.000 322.960 ;
    END
  END ram_val_in[3]
  PIN ram_val_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 646.000 99.320 650.000 99.920 ;
    END
  END ram_val_out[0]
  PIN ram_val_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 646.000 182.960 650.000 183.560 ;
    END
  END ram_val_out[1]
  PIN ram_val_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 646.000 266.600 650.000 267.200 ;
    END
  END ram_val_out[2]
  PIN ram_val_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 646.000 350.240 650.000 350.840 ;
    END
  END ram_val_out[3]
  PIN ram_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 646.000 15.680 650.000 16.280 ;
    END
  END ram_we
  PIN rom_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END rom_addr[0]
  PIN rom_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END rom_addr[1]
  PIN rom_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 4.000 67.280 ;
    END
  END rom_addr[2]
  PIN rom_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END rom_addr[3]
  PIN rom_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 4.000 108.080 ;
    END
  END rom_addr[4]
  PIN rom_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END rom_addr[5]
  PIN rom_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 4.000 148.880 ;
    END
  END rom_addr[6]
  PIN rom_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 4.000 169.280 ;
    END
  END rom_addr[7]
  PIN rom_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 4.000 189.680 ;
    END
  END rom_addr[8]
  PIN rom_csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.680 4.000 16.280 ;
    END
  END rom_csb
  PIN rom_value[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.080 4.000 36.680 ;
    END
  END rom_value[0]
  PIN rom_value[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.680 4.000 220.280 ;
    END
  END rom_value[10]
  PIN rom_value[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.880 4.000 230.480 ;
    END
  END rom_value[11]
  PIN rom_value[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.080 4.000 240.680 ;
    END
  END rom_value[12]
  PIN rom_value[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.280 4.000 250.880 ;
    END
  END rom_value[13]
  PIN rom_value[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 260.480 4.000 261.080 ;
    END
  END rom_value[14]
  PIN rom_value[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.680 4.000 271.280 ;
    END
  END rom_value[15]
  PIN rom_value[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.880 4.000 281.480 ;
    END
  END rom_value[16]
  PIN rom_value[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.080 4.000 291.680 ;
    END
  END rom_value[17]
  PIN rom_value[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.280 4.000 301.880 ;
    END
  END rom_value[18]
  PIN rom_value[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 311.480 4.000 312.080 ;
    END
  END rom_value[19]
  PIN rom_value[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.480 4.000 57.080 ;
    END
  END rom_value[1]
  PIN rom_value[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.680 4.000 322.280 ;
    END
  END rom_value[20]
  PIN rom_value[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.880 4.000 332.480 ;
    END
  END rom_value[21]
  PIN rom_value[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.080 4.000 342.680 ;
    END
  END rom_value[22]
  PIN rom_value[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.280 4.000 352.880 ;
    END
  END rom_value[23]
  PIN rom_value[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 362.480 4.000 363.080 ;
    END
  END rom_value[24]
  PIN rom_value[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 372.680 4.000 373.280 ;
    END
  END rom_value[25]
  PIN rom_value[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 382.880 4.000 383.480 ;
    END
  END rom_value[26]
  PIN rom_value[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.080 4.000 393.680 ;
    END
  END rom_value[27]
  PIN rom_value[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 403.280 4.000 403.880 ;
    END
  END rom_value[28]
  PIN rom_value[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 413.480 4.000 414.080 ;
    END
  END rom_value[29]
  PIN rom_value[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.880 4.000 77.480 ;
    END
  END rom_value[2]
  PIN rom_value[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 423.680 4.000 424.280 ;
    END
  END rom_value[30]
  PIN rom_value[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 433.880 4.000 434.480 ;
    END
  END rom_value[31]
  PIN rom_value[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.280 4.000 97.880 ;
    END
  END rom_value[3]
  PIN rom_value[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.680 4.000 118.280 ;
    END
  END rom_value[4]
  PIN rom_value[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.080 4.000 138.680 ;
    END
  END rom_value[5]
  PIN rom_value[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 158.480 4.000 159.080 ;
    END
  END rom_value[6]
  PIN rom_value[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.880 4.000 179.480 ;
    END
  END rom_value[7]
  PIN rom_value[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.280 4.000 199.880 ;
    END
  END rom_value[8]
  PIN rom_value[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END rom_value[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 438.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 438.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 438.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 438.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 438.160 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 438.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 438.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 438.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 438.160 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 0.000 20.610 4.000 ;
    END
  END wb_clk_i
  PIN wb_rom_adrb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 4.000 ;
    END
  END wb_rom_adrb[0]
  PIN wb_rom_adrb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END wb_rom_adrb[1]
  PIN wb_rom_adrb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 0.000 53.730 4.000 ;
    END
  END wb_rom_adrb[2]
  PIN wb_rom_adrb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 0.000 62.010 4.000 ;
    END
  END wb_rom_adrb[3]
  PIN wb_rom_adrb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 0.000 70.290 4.000 ;
    END
  END wb_rom_adrb[4]
  PIN wb_rom_adrb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 0.000 78.570 4.000 ;
    END
  END wb_rom_adrb[5]
  PIN wb_rom_adrb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.570 0.000 86.850 4.000 ;
    END
  END wb_rom_adrb[6]
  PIN wb_rom_adrb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 0.000 95.130 4.000 ;
    END
  END wb_rom_adrb[7]
  PIN wb_rom_adrb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END wb_rom_adrb[8]
  PIN wb_rom_csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.470 0.000 24.750 4.000 ;
    END
  END wb_rom_csb
  PIN wb_rom_val[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 0.000 41.310 4.000 ;
    END
  END wb_rom_val[0]
  PIN wb_rom_val[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 0.000 115.830 4.000 ;
    END
  END wb_rom_val[10]
  PIN wb_rom_val[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END wb_rom_val[11]
  PIN wb_rom_val[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.830 0.000 124.110 4.000 ;
    END
  END wb_rom_val[12]
  PIN wb_rom_val[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.970 0.000 128.250 4.000 ;
    END
  END wb_rom_val[13]
  PIN wb_rom_val[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END wb_rom_val[14]
  PIN wb_rom_val[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.250 0.000 136.530 4.000 ;
    END
  END wb_rom_val[15]
  PIN wb_rom_val[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 0.000 140.670 4.000 ;
    END
  END wb_rom_val[16]
  PIN wb_rom_val[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 0.000 144.810 4.000 ;
    END
  END wb_rom_val[17]
  PIN wb_rom_val[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.670 0.000 148.950 4.000 ;
    END
  END wb_rom_val[18]
  PIN wb_rom_val[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.810 0.000 153.090 4.000 ;
    END
  END wb_rom_val[19]
  PIN wb_rom_val[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 0.000 49.590 4.000 ;
    END
  END wb_rom_val[1]
  PIN wb_rom_val[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.950 0.000 157.230 4.000 ;
    END
  END wb_rom_val[20]
  PIN wb_rom_val[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END wb_rom_val[21]
  PIN wb_rom_val[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.230 0.000 165.510 4.000 ;
    END
  END wb_rom_val[22]
  PIN wb_rom_val[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.370 0.000 169.650 4.000 ;
    END
  END wb_rom_val[23]
  PIN wb_rom_val[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.510 0.000 173.790 4.000 ;
    END
  END wb_rom_val[24]
  PIN wb_rom_val[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.650 0.000 177.930 4.000 ;
    END
  END wb_rom_val[25]
  PIN wb_rom_val[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.790 0.000 182.070 4.000 ;
    END
  END wb_rom_val[26]
  PIN wb_rom_val[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 0.000 186.210 4.000 ;
    END
  END wb_rom_val[27]
  PIN wb_rom_val[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 4.000 ;
    END
  END wb_rom_val[28]
  PIN wb_rom_val[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.210 0.000 194.490 4.000 ;
    END
  END wb_rom_val[29]
  PIN wb_rom_val[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 0.000 57.870 4.000 ;
    END
  END wb_rom_val[2]
  PIN wb_rom_val[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.350 0.000 198.630 4.000 ;
    END
  END wb_rom_val[30]
  PIN wb_rom_val[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.490 0.000 202.770 4.000 ;
    END
  END wb_rom_val[31]
  PIN wb_rom_val[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 0.000 66.150 4.000 ;
    END
  END wb_rom_val[3]
  PIN wb_rom_val[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END wb_rom_val[4]
  PIN wb_rom_val[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 0.000 82.710 4.000 ;
    END
  END wb_rom_val[5]
  PIN wb_rom_val[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 0.000 90.990 4.000 ;
    END
  END wb_rom_val[6]
  PIN wb_rom_val[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.990 0.000 99.270 4.000 ;
    END
  END wb_rom_val[7]
  PIN wb_rom_val[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.270 0.000 107.550 4.000 ;
    END
  END wb_rom_val[8]
  PIN wb_rom_val[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.410 0.000 111.690 4.000 ;
    END
  END wb_rom_val[9]
  PIN wb_rom_web
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 4.000 ;
    END
  END wb_rom_web
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.750 0.000 33.030 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.630 0.000 206.910 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.190 0.000 223.470 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.390 0.000 347.670 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.810 0.000 360.090 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.230 0.000 372.510 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.650 0.000 384.930 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.070 0.000 397.350 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.490 0.000 409.770 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 0.000 422.190 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.330 0.000 434.610 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.750 0.000 447.030 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.170 0.000 459.450 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.610 0.000 235.890 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.590 0.000 471.870 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.010 0.000 484.290 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.430 0.000 496.710 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 0.000 509.130 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.270 0.000 521.550 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.690 0.000 533.970 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.110 0.000 546.390 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.530 0.000 558.810 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.950 0.000 571.230 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.370 0.000 583.650 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 0.000 248.310 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.790 0.000 596.070 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.210 0.000 608.490 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.450 0.000 260.730 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.870 0.000 273.150 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.290 0.000 285.570 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.710 0.000 297.990 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.130 0.000 310.410 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.550 0.000 322.830 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 0.000 335.250 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.770 0.000 211.050 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.330 0.000 227.610 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.530 0.000 351.810 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 0.000 364.230 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.370 0.000 376.650 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.790 0.000 389.070 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.210 0.000 401.490 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.630 0.000 413.910 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.050 0.000 426.330 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.470 0.000 438.750 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 0.000 451.170 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.310 0.000 463.590 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.750 0.000 240.030 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.730 0.000 476.010 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.150 0.000 488.430 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.570 0.000 500.850 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.990 0.000 513.270 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.410 0.000 525.690 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.830 0.000 538.110 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.250 0.000 550.530 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.670 0.000 562.950 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.090 0.000 575.370 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.510 0.000 587.790 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.170 0.000 252.450 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.930 0.000 600.210 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.350 0.000 612.630 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.590 0.000 264.870 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.430 0.000 289.710 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.850 0.000 302.130 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.270 0.000 314.550 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.690 0.000 326.970 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.110 0.000 339.390 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.470 0.000 231.750 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.670 0.000 355.950 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.090 0.000 368.370 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.510 0.000 380.790 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 0.000 393.210 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.350 0.000 405.630 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.770 0.000 418.050 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.190 0.000 430.470 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.610 0.000 442.890 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.030 0.000 455.310 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.450 0.000 467.730 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.890 0.000 244.170 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 0.000 480.150 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.290 0.000 492.570 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.710 0.000 504.990 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.130 0.000 517.410 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.550 0.000 529.830 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.970 0.000 542.250 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 554.390 0.000 554.670 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.810 0.000 567.090 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.230 0.000 579.510 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.650 0.000 591.930 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.310 0.000 256.590 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.070 0.000 604.350 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.490 0.000 616.770 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.730 0.000 269.010 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.150 0.000 281.430 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 0.000 293.850 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.410 0.000 318.690 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.830 0.000 331.110 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.250 0.000 343.530 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.910 0.000 215.190 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 644.460 438.005 ;
      LAYER met1 ;
        RECT 4.670 0.380 645.310 438.160 ;
      LAYER met2 ;
        RECT 4.690 445.720 12.690 446.490 ;
        RECT 13.530 445.720 18.210 446.490 ;
        RECT 19.050 445.720 23.730 446.490 ;
        RECT 24.570 445.720 29.250 446.490 ;
        RECT 30.090 445.720 34.770 446.490 ;
        RECT 35.610 445.720 40.290 446.490 ;
        RECT 41.130 445.720 45.810 446.490 ;
        RECT 46.650 445.720 51.330 446.490 ;
        RECT 52.170 445.720 56.850 446.490 ;
        RECT 57.690 445.720 62.370 446.490 ;
        RECT 63.210 445.720 67.890 446.490 ;
        RECT 68.730 445.720 73.410 446.490 ;
        RECT 74.250 445.720 78.930 446.490 ;
        RECT 79.770 445.720 84.450 446.490 ;
        RECT 85.290 445.720 89.970 446.490 ;
        RECT 90.810 445.720 95.490 446.490 ;
        RECT 96.330 445.720 101.010 446.490 ;
        RECT 101.850 445.720 106.530 446.490 ;
        RECT 107.370 445.720 112.050 446.490 ;
        RECT 112.890 445.720 117.570 446.490 ;
        RECT 118.410 445.720 123.090 446.490 ;
        RECT 123.930 445.720 128.610 446.490 ;
        RECT 129.450 445.720 134.130 446.490 ;
        RECT 134.970 445.720 139.650 446.490 ;
        RECT 140.490 445.720 145.170 446.490 ;
        RECT 146.010 445.720 150.690 446.490 ;
        RECT 151.530 445.720 156.210 446.490 ;
        RECT 157.050 445.720 161.730 446.490 ;
        RECT 162.570 445.720 167.250 446.490 ;
        RECT 168.090 445.720 172.770 446.490 ;
        RECT 173.610 445.720 178.290 446.490 ;
        RECT 179.130 445.720 183.810 446.490 ;
        RECT 184.650 445.720 189.330 446.490 ;
        RECT 190.170 445.720 194.850 446.490 ;
        RECT 195.690 445.720 200.370 446.490 ;
        RECT 201.210 445.720 205.890 446.490 ;
        RECT 206.730 445.720 211.410 446.490 ;
        RECT 212.250 445.720 216.930 446.490 ;
        RECT 217.770 445.720 222.450 446.490 ;
        RECT 223.290 445.720 227.970 446.490 ;
        RECT 228.810 445.720 233.490 446.490 ;
        RECT 234.330 445.720 239.010 446.490 ;
        RECT 239.850 445.720 244.530 446.490 ;
        RECT 245.370 445.720 250.050 446.490 ;
        RECT 250.890 445.720 255.570 446.490 ;
        RECT 256.410 445.720 261.090 446.490 ;
        RECT 261.930 445.720 266.610 446.490 ;
        RECT 267.450 445.720 272.130 446.490 ;
        RECT 272.970 445.720 277.650 446.490 ;
        RECT 278.490 445.720 283.170 446.490 ;
        RECT 284.010 445.720 288.690 446.490 ;
        RECT 289.530 445.720 294.210 446.490 ;
        RECT 295.050 445.720 299.730 446.490 ;
        RECT 300.570 445.720 305.250 446.490 ;
        RECT 306.090 445.720 310.770 446.490 ;
        RECT 311.610 445.720 316.290 446.490 ;
        RECT 317.130 445.720 321.810 446.490 ;
        RECT 322.650 445.720 327.330 446.490 ;
        RECT 328.170 445.720 332.850 446.490 ;
        RECT 333.690 445.720 338.370 446.490 ;
        RECT 339.210 445.720 343.890 446.490 ;
        RECT 344.730 445.720 349.410 446.490 ;
        RECT 350.250 445.720 354.930 446.490 ;
        RECT 355.770 445.720 360.450 446.490 ;
        RECT 361.290 445.720 365.970 446.490 ;
        RECT 366.810 445.720 371.490 446.490 ;
        RECT 372.330 445.720 377.010 446.490 ;
        RECT 377.850 445.720 382.530 446.490 ;
        RECT 383.370 445.720 388.050 446.490 ;
        RECT 388.890 445.720 393.570 446.490 ;
        RECT 394.410 445.720 399.090 446.490 ;
        RECT 399.930 445.720 404.610 446.490 ;
        RECT 405.450 445.720 410.130 446.490 ;
        RECT 410.970 445.720 415.650 446.490 ;
        RECT 416.490 445.720 421.170 446.490 ;
        RECT 422.010 445.720 426.690 446.490 ;
        RECT 427.530 445.720 432.210 446.490 ;
        RECT 433.050 445.720 437.730 446.490 ;
        RECT 438.570 445.720 443.250 446.490 ;
        RECT 444.090 445.720 448.770 446.490 ;
        RECT 449.610 445.720 454.290 446.490 ;
        RECT 455.130 445.720 459.810 446.490 ;
        RECT 460.650 445.720 465.330 446.490 ;
        RECT 466.170 445.720 470.850 446.490 ;
        RECT 471.690 445.720 476.370 446.490 ;
        RECT 477.210 445.720 481.890 446.490 ;
        RECT 482.730 445.720 487.410 446.490 ;
        RECT 488.250 445.720 492.930 446.490 ;
        RECT 493.770 445.720 498.450 446.490 ;
        RECT 499.290 445.720 503.970 446.490 ;
        RECT 504.810 445.720 509.490 446.490 ;
        RECT 510.330 445.720 515.010 446.490 ;
        RECT 515.850 445.720 520.530 446.490 ;
        RECT 521.370 445.720 526.050 446.490 ;
        RECT 526.890 445.720 531.570 446.490 ;
        RECT 532.410 445.720 537.090 446.490 ;
        RECT 537.930 445.720 542.610 446.490 ;
        RECT 543.450 445.720 548.130 446.490 ;
        RECT 548.970 445.720 553.650 446.490 ;
        RECT 554.490 445.720 559.170 446.490 ;
        RECT 560.010 445.720 564.690 446.490 ;
        RECT 565.530 445.720 570.210 446.490 ;
        RECT 571.050 445.720 575.730 446.490 ;
        RECT 576.570 445.720 581.250 446.490 ;
        RECT 582.090 445.720 586.770 446.490 ;
        RECT 587.610 445.720 592.290 446.490 ;
        RECT 593.130 445.720 597.810 446.490 ;
        RECT 598.650 445.720 603.330 446.490 ;
        RECT 604.170 445.720 608.850 446.490 ;
        RECT 609.690 445.720 614.370 446.490 ;
        RECT 615.210 445.720 619.890 446.490 ;
        RECT 620.730 445.720 625.410 446.490 ;
        RECT 626.250 445.720 630.930 446.490 ;
        RECT 631.770 445.720 636.450 446.490 ;
        RECT 637.290 445.720 645.290 446.490 ;
        RECT 4.690 4.280 645.290 445.720 ;
        RECT 4.690 0.350 20.050 4.280 ;
        RECT 20.890 0.350 24.190 4.280 ;
        RECT 25.030 0.350 28.330 4.280 ;
        RECT 29.170 0.350 32.470 4.280 ;
        RECT 33.310 0.350 36.610 4.280 ;
        RECT 37.450 0.350 40.750 4.280 ;
        RECT 41.590 0.350 44.890 4.280 ;
        RECT 45.730 0.350 49.030 4.280 ;
        RECT 49.870 0.350 53.170 4.280 ;
        RECT 54.010 0.350 57.310 4.280 ;
        RECT 58.150 0.350 61.450 4.280 ;
        RECT 62.290 0.350 65.590 4.280 ;
        RECT 66.430 0.350 69.730 4.280 ;
        RECT 70.570 0.350 73.870 4.280 ;
        RECT 74.710 0.350 78.010 4.280 ;
        RECT 78.850 0.350 82.150 4.280 ;
        RECT 82.990 0.350 86.290 4.280 ;
        RECT 87.130 0.350 90.430 4.280 ;
        RECT 91.270 0.350 94.570 4.280 ;
        RECT 95.410 0.350 98.710 4.280 ;
        RECT 99.550 0.350 102.850 4.280 ;
        RECT 103.690 0.350 106.990 4.280 ;
        RECT 107.830 0.350 111.130 4.280 ;
        RECT 111.970 0.350 115.270 4.280 ;
        RECT 116.110 0.350 119.410 4.280 ;
        RECT 120.250 0.350 123.550 4.280 ;
        RECT 124.390 0.350 127.690 4.280 ;
        RECT 128.530 0.350 131.830 4.280 ;
        RECT 132.670 0.350 135.970 4.280 ;
        RECT 136.810 0.350 140.110 4.280 ;
        RECT 140.950 0.350 144.250 4.280 ;
        RECT 145.090 0.350 148.390 4.280 ;
        RECT 149.230 0.350 152.530 4.280 ;
        RECT 153.370 0.350 156.670 4.280 ;
        RECT 157.510 0.350 160.810 4.280 ;
        RECT 161.650 0.350 164.950 4.280 ;
        RECT 165.790 0.350 169.090 4.280 ;
        RECT 169.930 0.350 173.230 4.280 ;
        RECT 174.070 0.350 177.370 4.280 ;
        RECT 178.210 0.350 181.510 4.280 ;
        RECT 182.350 0.350 185.650 4.280 ;
        RECT 186.490 0.350 189.790 4.280 ;
        RECT 190.630 0.350 193.930 4.280 ;
        RECT 194.770 0.350 198.070 4.280 ;
        RECT 198.910 0.350 202.210 4.280 ;
        RECT 203.050 0.350 206.350 4.280 ;
        RECT 207.190 0.350 210.490 4.280 ;
        RECT 211.330 0.350 214.630 4.280 ;
        RECT 215.470 0.350 218.770 4.280 ;
        RECT 219.610 0.350 222.910 4.280 ;
        RECT 223.750 0.350 227.050 4.280 ;
        RECT 227.890 0.350 231.190 4.280 ;
        RECT 232.030 0.350 235.330 4.280 ;
        RECT 236.170 0.350 239.470 4.280 ;
        RECT 240.310 0.350 243.610 4.280 ;
        RECT 244.450 0.350 247.750 4.280 ;
        RECT 248.590 0.350 251.890 4.280 ;
        RECT 252.730 0.350 256.030 4.280 ;
        RECT 256.870 0.350 260.170 4.280 ;
        RECT 261.010 0.350 264.310 4.280 ;
        RECT 265.150 0.350 268.450 4.280 ;
        RECT 269.290 0.350 272.590 4.280 ;
        RECT 273.430 0.350 276.730 4.280 ;
        RECT 277.570 0.350 280.870 4.280 ;
        RECT 281.710 0.350 285.010 4.280 ;
        RECT 285.850 0.350 289.150 4.280 ;
        RECT 289.990 0.350 293.290 4.280 ;
        RECT 294.130 0.350 297.430 4.280 ;
        RECT 298.270 0.350 301.570 4.280 ;
        RECT 302.410 0.350 305.710 4.280 ;
        RECT 306.550 0.350 309.850 4.280 ;
        RECT 310.690 0.350 313.990 4.280 ;
        RECT 314.830 0.350 318.130 4.280 ;
        RECT 318.970 0.350 322.270 4.280 ;
        RECT 323.110 0.350 326.410 4.280 ;
        RECT 327.250 0.350 330.550 4.280 ;
        RECT 331.390 0.350 334.690 4.280 ;
        RECT 335.530 0.350 338.830 4.280 ;
        RECT 339.670 0.350 342.970 4.280 ;
        RECT 343.810 0.350 347.110 4.280 ;
        RECT 347.950 0.350 351.250 4.280 ;
        RECT 352.090 0.350 355.390 4.280 ;
        RECT 356.230 0.350 359.530 4.280 ;
        RECT 360.370 0.350 363.670 4.280 ;
        RECT 364.510 0.350 367.810 4.280 ;
        RECT 368.650 0.350 371.950 4.280 ;
        RECT 372.790 0.350 376.090 4.280 ;
        RECT 376.930 0.350 380.230 4.280 ;
        RECT 381.070 0.350 384.370 4.280 ;
        RECT 385.210 0.350 388.510 4.280 ;
        RECT 389.350 0.350 392.650 4.280 ;
        RECT 393.490 0.350 396.790 4.280 ;
        RECT 397.630 0.350 400.930 4.280 ;
        RECT 401.770 0.350 405.070 4.280 ;
        RECT 405.910 0.350 409.210 4.280 ;
        RECT 410.050 0.350 413.350 4.280 ;
        RECT 414.190 0.350 417.490 4.280 ;
        RECT 418.330 0.350 421.630 4.280 ;
        RECT 422.470 0.350 425.770 4.280 ;
        RECT 426.610 0.350 429.910 4.280 ;
        RECT 430.750 0.350 434.050 4.280 ;
        RECT 434.890 0.350 438.190 4.280 ;
        RECT 439.030 0.350 442.330 4.280 ;
        RECT 443.170 0.350 446.470 4.280 ;
        RECT 447.310 0.350 450.610 4.280 ;
        RECT 451.450 0.350 454.750 4.280 ;
        RECT 455.590 0.350 458.890 4.280 ;
        RECT 459.730 0.350 463.030 4.280 ;
        RECT 463.870 0.350 467.170 4.280 ;
        RECT 468.010 0.350 471.310 4.280 ;
        RECT 472.150 0.350 475.450 4.280 ;
        RECT 476.290 0.350 479.590 4.280 ;
        RECT 480.430 0.350 483.730 4.280 ;
        RECT 484.570 0.350 487.870 4.280 ;
        RECT 488.710 0.350 492.010 4.280 ;
        RECT 492.850 0.350 496.150 4.280 ;
        RECT 496.990 0.350 500.290 4.280 ;
        RECT 501.130 0.350 504.430 4.280 ;
        RECT 505.270 0.350 508.570 4.280 ;
        RECT 509.410 0.350 512.710 4.280 ;
        RECT 513.550 0.350 516.850 4.280 ;
        RECT 517.690 0.350 520.990 4.280 ;
        RECT 521.830 0.350 525.130 4.280 ;
        RECT 525.970 0.350 529.270 4.280 ;
        RECT 530.110 0.350 533.410 4.280 ;
        RECT 534.250 0.350 537.550 4.280 ;
        RECT 538.390 0.350 541.690 4.280 ;
        RECT 542.530 0.350 545.830 4.280 ;
        RECT 546.670 0.350 549.970 4.280 ;
        RECT 550.810 0.350 554.110 4.280 ;
        RECT 554.950 0.350 558.250 4.280 ;
        RECT 559.090 0.350 562.390 4.280 ;
        RECT 563.230 0.350 566.530 4.280 ;
        RECT 567.370 0.350 570.670 4.280 ;
        RECT 571.510 0.350 574.810 4.280 ;
        RECT 575.650 0.350 578.950 4.280 ;
        RECT 579.790 0.350 583.090 4.280 ;
        RECT 583.930 0.350 587.230 4.280 ;
        RECT 588.070 0.350 591.370 4.280 ;
        RECT 592.210 0.350 595.510 4.280 ;
        RECT 596.350 0.350 599.650 4.280 ;
        RECT 600.490 0.350 603.790 4.280 ;
        RECT 604.630 0.350 607.930 4.280 ;
        RECT 608.770 0.350 612.070 4.280 ;
        RECT 612.910 0.350 616.210 4.280 ;
        RECT 617.050 0.350 620.350 4.280 ;
        RECT 621.190 0.350 624.490 4.280 ;
        RECT 625.330 0.350 628.630 4.280 ;
        RECT 629.470 0.350 645.290 4.280 ;
      LAYER met3 ;
        RECT 4.000 434.880 646.000 438.085 ;
        RECT 4.400 433.480 645.600 434.880 ;
        RECT 4.000 424.680 646.000 433.480 ;
        RECT 4.400 423.280 646.000 424.680 ;
        RECT 4.000 414.480 646.000 423.280 ;
        RECT 4.400 413.080 646.000 414.480 ;
        RECT 4.000 407.000 646.000 413.080 ;
        RECT 4.000 405.600 645.600 407.000 ;
        RECT 4.000 404.280 646.000 405.600 ;
        RECT 4.400 402.880 646.000 404.280 ;
        RECT 4.000 394.080 646.000 402.880 ;
        RECT 4.400 392.680 646.000 394.080 ;
        RECT 4.000 383.880 646.000 392.680 ;
        RECT 4.400 382.480 646.000 383.880 ;
        RECT 4.000 379.120 646.000 382.480 ;
        RECT 4.000 377.720 645.600 379.120 ;
        RECT 4.000 373.680 646.000 377.720 ;
        RECT 4.400 372.280 646.000 373.680 ;
        RECT 4.000 363.480 646.000 372.280 ;
        RECT 4.400 362.080 646.000 363.480 ;
        RECT 4.000 353.280 646.000 362.080 ;
        RECT 4.400 351.880 646.000 353.280 ;
        RECT 4.000 351.240 646.000 351.880 ;
        RECT 4.000 349.840 645.600 351.240 ;
        RECT 4.000 343.080 646.000 349.840 ;
        RECT 4.400 341.680 646.000 343.080 ;
        RECT 4.000 332.880 646.000 341.680 ;
        RECT 4.400 331.480 646.000 332.880 ;
        RECT 4.000 323.360 646.000 331.480 ;
        RECT 4.000 322.680 645.600 323.360 ;
        RECT 4.400 321.960 645.600 322.680 ;
        RECT 4.400 321.280 646.000 321.960 ;
        RECT 4.000 312.480 646.000 321.280 ;
        RECT 4.400 311.080 646.000 312.480 ;
        RECT 4.000 302.280 646.000 311.080 ;
        RECT 4.400 300.880 646.000 302.280 ;
        RECT 4.000 295.480 646.000 300.880 ;
        RECT 4.000 294.080 645.600 295.480 ;
        RECT 4.000 292.080 646.000 294.080 ;
        RECT 4.400 290.680 646.000 292.080 ;
        RECT 4.000 281.880 646.000 290.680 ;
        RECT 4.400 280.480 646.000 281.880 ;
        RECT 4.000 271.680 646.000 280.480 ;
        RECT 4.400 270.280 646.000 271.680 ;
        RECT 4.000 267.600 646.000 270.280 ;
        RECT 4.000 266.200 645.600 267.600 ;
        RECT 4.000 261.480 646.000 266.200 ;
        RECT 4.400 260.080 646.000 261.480 ;
        RECT 4.000 251.280 646.000 260.080 ;
        RECT 4.400 249.880 646.000 251.280 ;
        RECT 4.000 241.080 646.000 249.880 ;
        RECT 4.400 239.720 646.000 241.080 ;
        RECT 4.400 239.680 645.600 239.720 ;
        RECT 4.000 238.320 645.600 239.680 ;
        RECT 4.000 230.880 646.000 238.320 ;
        RECT 4.400 229.480 646.000 230.880 ;
        RECT 4.000 220.680 646.000 229.480 ;
        RECT 4.400 219.280 646.000 220.680 ;
        RECT 4.000 211.840 646.000 219.280 ;
        RECT 4.000 210.480 645.600 211.840 ;
        RECT 4.400 210.440 645.600 210.480 ;
        RECT 4.400 209.080 646.000 210.440 ;
        RECT 4.000 200.280 646.000 209.080 ;
        RECT 4.400 198.880 646.000 200.280 ;
        RECT 4.000 190.080 646.000 198.880 ;
        RECT 4.400 188.680 646.000 190.080 ;
        RECT 4.000 183.960 646.000 188.680 ;
        RECT 4.000 182.560 645.600 183.960 ;
        RECT 4.000 179.880 646.000 182.560 ;
        RECT 4.400 178.480 646.000 179.880 ;
        RECT 4.000 169.680 646.000 178.480 ;
        RECT 4.400 168.280 646.000 169.680 ;
        RECT 4.000 159.480 646.000 168.280 ;
        RECT 4.400 158.080 646.000 159.480 ;
        RECT 4.000 156.080 646.000 158.080 ;
        RECT 4.000 154.680 645.600 156.080 ;
        RECT 4.000 149.280 646.000 154.680 ;
        RECT 4.400 147.880 646.000 149.280 ;
        RECT 4.000 139.080 646.000 147.880 ;
        RECT 4.400 137.680 646.000 139.080 ;
        RECT 4.000 128.880 646.000 137.680 ;
        RECT 4.400 128.200 646.000 128.880 ;
        RECT 4.400 127.480 645.600 128.200 ;
        RECT 4.000 126.800 645.600 127.480 ;
        RECT 4.000 118.680 646.000 126.800 ;
        RECT 4.400 117.280 646.000 118.680 ;
        RECT 4.000 108.480 646.000 117.280 ;
        RECT 4.400 107.080 646.000 108.480 ;
        RECT 4.000 100.320 646.000 107.080 ;
        RECT 4.000 98.920 645.600 100.320 ;
        RECT 4.000 98.280 646.000 98.920 ;
        RECT 4.400 96.880 646.000 98.280 ;
        RECT 4.000 88.080 646.000 96.880 ;
        RECT 4.400 86.680 646.000 88.080 ;
        RECT 4.000 77.880 646.000 86.680 ;
        RECT 4.400 76.480 646.000 77.880 ;
        RECT 4.000 72.440 646.000 76.480 ;
        RECT 4.000 71.040 645.600 72.440 ;
        RECT 4.000 67.680 646.000 71.040 ;
        RECT 4.400 66.280 646.000 67.680 ;
        RECT 4.000 57.480 646.000 66.280 ;
        RECT 4.400 56.080 646.000 57.480 ;
        RECT 4.000 47.280 646.000 56.080 ;
        RECT 4.400 45.880 646.000 47.280 ;
        RECT 4.000 44.560 646.000 45.880 ;
        RECT 4.000 43.160 645.600 44.560 ;
        RECT 4.000 37.080 646.000 43.160 ;
        RECT 4.400 35.680 646.000 37.080 ;
        RECT 4.000 26.880 646.000 35.680 ;
        RECT 4.400 25.480 646.000 26.880 ;
        RECT 4.000 16.680 646.000 25.480 ;
        RECT 4.400 15.280 645.600 16.680 ;
        RECT 4.000 8.335 646.000 15.280 ;
      LAYER met4 ;
        RECT 9.495 13.095 20.640 437.065 ;
        RECT 23.040 13.095 97.440 437.065 ;
        RECT 99.840 13.095 174.240 437.065 ;
        RECT 176.640 13.095 251.040 437.065 ;
        RECT 253.440 13.095 327.840 437.065 ;
        RECT 330.240 13.095 404.640 437.065 ;
        RECT 407.040 13.095 481.440 437.065 ;
        RECT 483.840 13.095 558.240 437.065 ;
        RECT 560.640 13.095 589.425 437.065 ;
  END
END wrapped_tms1x00
END LIBRARY

