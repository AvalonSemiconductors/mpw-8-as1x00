magic
tech sky130B
magscale 1 2
timestamp 1671698854
<< obsli1 >>
rect 1104 2159 88872 47345
<< obsm1 >>
rect 1104 416 88872 47456
<< metal2 >>
rect 3330 49200 3386 50000
rect 4066 49200 4122 50000
rect 4802 49200 4858 50000
rect 5538 49200 5594 50000
rect 6274 49200 6330 50000
rect 7010 49200 7066 50000
rect 7746 49200 7802 50000
rect 8482 49200 8538 50000
rect 9218 49200 9274 50000
rect 9954 49200 10010 50000
rect 10690 49200 10746 50000
rect 11426 49200 11482 50000
rect 12162 49200 12218 50000
rect 12898 49200 12954 50000
rect 13634 49200 13690 50000
rect 14370 49200 14426 50000
rect 15106 49200 15162 50000
rect 15842 49200 15898 50000
rect 16578 49200 16634 50000
rect 17314 49200 17370 50000
rect 18050 49200 18106 50000
rect 18786 49200 18842 50000
rect 19522 49200 19578 50000
rect 20258 49200 20314 50000
rect 20994 49200 21050 50000
rect 21730 49200 21786 50000
rect 22466 49200 22522 50000
rect 23202 49200 23258 50000
rect 23938 49200 23994 50000
rect 24674 49200 24730 50000
rect 25410 49200 25466 50000
rect 26146 49200 26202 50000
rect 26882 49200 26938 50000
rect 27618 49200 27674 50000
rect 28354 49200 28410 50000
rect 29090 49200 29146 50000
rect 29826 49200 29882 50000
rect 30562 49200 30618 50000
rect 31298 49200 31354 50000
rect 32034 49200 32090 50000
rect 32770 49200 32826 50000
rect 33506 49200 33562 50000
rect 34242 49200 34298 50000
rect 34978 49200 35034 50000
rect 35714 49200 35770 50000
rect 36450 49200 36506 50000
rect 37186 49200 37242 50000
rect 37922 49200 37978 50000
rect 38658 49200 38714 50000
rect 39394 49200 39450 50000
rect 40130 49200 40186 50000
rect 40866 49200 40922 50000
rect 41602 49200 41658 50000
rect 42338 49200 42394 50000
rect 43074 49200 43130 50000
rect 43810 49200 43866 50000
rect 44546 49200 44602 50000
rect 45282 49200 45338 50000
rect 46018 49200 46074 50000
rect 46754 49200 46810 50000
rect 47490 49200 47546 50000
rect 48226 49200 48282 50000
rect 48962 49200 49018 50000
rect 49698 49200 49754 50000
rect 50434 49200 50490 50000
rect 51170 49200 51226 50000
rect 51906 49200 51962 50000
rect 52642 49200 52698 50000
rect 53378 49200 53434 50000
rect 54114 49200 54170 50000
rect 54850 49200 54906 50000
rect 55586 49200 55642 50000
rect 56322 49200 56378 50000
rect 57058 49200 57114 50000
rect 57794 49200 57850 50000
rect 58530 49200 58586 50000
rect 59266 49200 59322 50000
rect 60002 49200 60058 50000
rect 60738 49200 60794 50000
rect 61474 49200 61530 50000
rect 62210 49200 62266 50000
rect 62946 49200 63002 50000
rect 63682 49200 63738 50000
rect 64418 49200 64474 50000
rect 65154 49200 65210 50000
rect 65890 49200 65946 50000
rect 66626 49200 66682 50000
rect 67362 49200 67418 50000
rect 68098 49200 68154 50000
rect 68834 49200 68890 50000
rect 69570 49200 69626 50000
rect 70306 49200 70362 50000
rect 71042 49200 71098 50000
rect 71778 49200 71834 50000
rect 72514 49200 72570 50000
rect 73250 49200 73306 50000
rect 73986 49200 74042 50000
rect 74722 49200 74778 50000
rect 75458 49200 75514 50000
rect 76194 49200 76250 50000
rect 76930 49200 76986 50000
rect 77666 49200 77722 50000
rect 78402 49200 78458 50000
rect 79138 49200 79194 50000
rect 79874 49200 79930 50000
rect 80610 49200 80666 50000
rect 81346 49200 81402 50000
rect 82082 49200 82138 50000
rect 82818 49200 82874 50000
rect 83554 49200 83610 50000
rect 84290 49200 84346 50000
rect 85026 49200 85082 50000
rect 85762 49200 85818 50000
rect 86498 49200 86554 50000
rect 5170 0 5226 800
rect 5722 0 5778 800
rect 6274 0 6330 800
rect 6826 0 6882 800
rect 7378 0 7434 800
rect 7930 0 7986 800
rect 8482 0 8538 800
rect 9034 0 9090 800
rect 9586 0 9642 800
rect 10138 0 10194 800
rect 10690 0 10746 800
rect 11242 0 11298 800
rect 11794 0 11850 800
rect 12346 0 12402 800
rect 12898 0 12954 800
rect 13450 0 13506 800
rect 14002 0 14058 800
rect 14554 0 14610 800
rect 15106 0 15162 800
rect 15658 0 15714 800
rect 16210 0 16266 800
rect 16762 0 16818 800
rect 17314 0 17370 800
rect 17866 0 17922 800
rect 18418 0 18474 800
rect 18970 0 19026 800
rect 19522 0 19578 800
rect 20074 0 20130 800
rect 20626 0 20682 800
rect 21178 0 21234 800
rect 21730 0 21786 800
rect 22282 0 22338 800
rect 22834 0 22890 800
rect 23386 0 23442 800
rect 23938 0 23994 800
rect 24490 0 24546 800
rect 25042 0 25098 800
rect 25594 0 25650 800
rect 26146 0 26202 800
rect 26698 0 26754 800
rect 27250 0 27306 800
rect 27802 0 27858 800
rect 28354 0 28410 800
rect 28906 0 28962 800
rect 29458 0 29514 800
rect 30010 0 30066 800
rect 30562 0 30618 800
rect 31114 0 31170 800
rect 31666 0 31722 800
rect 32218 0 32274 800
rect 32770 0 32826 800
rect 33322 0 33378 800
rect 33874 0 33930 800
rect 34426 0 34482 800
rect 34978 0 35034 800
rect 35530 0 35586 800
rect 36082 0 36138 800
rect 36634 0 36690 800
rect 37186 0 37242 800
rect 37738 0 37794 800
rect 38290 0 38346 800
rect 38842 0 38898 800
rect 39394 0 39450 800
rect 39946 0 40002 800
rect 40498 0 40554 800
rect 41050 0 41106 800
rect 41602 0 41658 800
rect 42154 0 42210 800
rect 42706 0 42762 800
rect 43258 0 43314 800
rect 43810 0 43866 800
rect 44362 0 44418 800
rect 44914 0 44970 800
rect 45466 0 45522 800
rect 46018 0 46074 800
rect 46570 0 46626 800
rect 47122 0 47178 800
rect 47674 0 47730 800
rect 48226 0 48282 800
rect 48778 0 48834 800
rect 49330 0 49386 800
rect 49882 0 49938 800
rect 50434 0 50490 800
rect 50986 0 51042 800
rect 51538 0 51594 800
rect 52090 0 52146 800
rect 52642 0 52698 800
rect 53194 0 53250 800
rect 53746 0 53802 800
rect 54298 0 54354 800
rect 54850 0 54906 800
rect 55402 0 55458 800
rect 55954 0 56010 800
rect 56506 0 56562 800
rect 57058 0 57114 800
rect 57610 0 57666 800
rect 58162 0 58218 800
rect 58714 0 58770 800
rect 59266 0 59322 800
rect 59818 0 59874 800
rect 60370 0 60426 800
rect 60922 0 60978 800
rect 61474 0 61530 800
rect 62026 0 62082 800
rect 62578 0 62634 800
rect 63130 0 63186 800
rect 63682 0 63738 800
rect 64234 0 64290 800
rect 64786 0 64842 800
rect 65338 0 65394 800
rect 65890 0 65946 800
rect 66442 0 66498 800
rect 66994 0 67050 800
rect 67546 0 67602 800
rect 68098 0 68154 800
rect 68650 0 68706 800
rect 69202 0 69258 800
rect 69754 0 69810 800
rect 70306 0 70362 800
rect 70858 0 70914 800
rect 71410 0 71466 800
rect 71962 0 72018 800
rect 72514 0 72570 800
rect 73066 0 73122 800
rect 73618 0 73674 800
rect 74170 0 74226 800
rect 74722 0 74778 800
rect 75274 0 75330 800
rect 75826 0 75882 800
rect 76378 0 76434 800
rect 76930 0 76986 800
rect 77482 0 77538 800
rect 78034 0 78090 800
rect 78586 0 78642 800
rect 79138 0 79194 800
rect 79690 0 79746 800
rect 80242 0 80298 800
rect 80794 0 80850 800
rect 81346 0 81402 800
rect 81898 0 81954 800
rect 82450 0 82506 800
rect 83002 0 83058 800
rect 83554 0 83610 800
rect 84106 0 84162 800
rect 84658 0 84714 800
<< obsm2 >>
rect 1400 49144 3274 49314
rect 3442 49144 4010 49314
rect 4178 49144 4746 49314
rect 4914 49144 5482 49314
rect 5650 49144 6218 49314
rect 6386 49144 6954 49314
rect 7122 49144 7690 49314
rect 7858 49144 8426 49314
rect 8594 49144 9162 49314
rect 9330 49144 9898 49314
rect 10066 49144 10634 49314
rect 10802 49144 11370 49314
rect 11538 49144 12106 49314
rect 12274 49144 12842 49314
rect 13010 49144 13578 49314
rect 13746 49144 14314 49314
rect 14482 49144 15050 49314
rect 15218 49144 15786 49314
rect 15954 49144 16522 49314
rect 16690 49144 17258 49314
rect 17426 49144 17994 49314
rect 18162 49144 18730 49314
rect 18898 49144 19466 49314
rect 19634 49144 20202 49314
rect 20370 49144 20938 49314
rect 21106 49144 21674 49314
rect 21842 49144 22410 49314
rect 22578 49144 23146 49314
rect 23314 49144 23882 49314
rect 24050 49144 24618 49314
rect 24786 49144 25354 49314
rect 25522 49144 26090 49314
rect 26258 49144 26826 49314
rect 26994 49144 27562 49314
rect 27730 49144 28298 49314
rect 28466 49144 29034 49314
rect 29202 49144 29770 49314
rect 29938 49144 30506 49314
rect 30674 49144 31242 49314
rect 31410 49144 31978 49314
rect 32146 49144 32714 49314
rect 32882 49144 33450 49314
rect 33618 49144 34186 49314
rect 34354 49144 34922 49314
rect 35090 49144 35658 49314
rect 35826 49144 36394 49314
rect 36562 49144 37130 49314
rect 37298 49144 37866 49314
rect 38034 49144 38602 49314
rect 38770 49144 39338 49314
rect 39506 49144 40074 49314
rect 40242 49144 40810 49314
rect 40978 49144 41546 49314
rect 41714 49144 42282 49314
rect 42450 49144 43018 49314
rect 43186 49144 43754 49314
rect 43922 49144 44490 49314
rect 44658 49144 45226 49314
rect 45394 49144 45962 49314
rect 46130 49144 46698 49314
rect 46866 49144 47434 49314
rect 47602 49144 48170 49314
rect 48338 49144 48906 49314
rect 49074 49144 49642 49314
rect 49810 49144 50378 49314
rect 50546 49144 51114 49314
rect 51282 49144 51850 49314
rect 52018 49144 52586 49314
rect 52754 49144 53322 49314
rect 53490 49144 54058 49314
rect 54226 49144 54794 49314
rect 54962 49144 55530 49314
rect 55698 49144 56266 49314
rect 56434 49144 57002 49314
rect 57170 49144 57738 49314
rect 57906 49144 58474 49314
rect 58642 49144 59210 49314
rect 59378 49144 59946 49314
rect 60114 49144 60682 49314
rect 60850 49144 61418 49314
rect 61586 49144 62154 49314
rect 62322 49144 62890 49314
rect 63058 49144 63626 49314
rect 63794 49144 64362 49314
rect 64530 49144 65098 49314
rect 65266 49144 65834 49314
rect 66002 49144 66570 49314
rect 66738 49144 67306 49314
rect 67474 49144 68042 49314
rect 68210 49144 68778 49314
rect 68946 49144 69514 49314
rect 69682 49144 70250 49314
rect 70418 49144 70986 49314
rect 71154 49144 71722 49314
rect 71890 49144 72458 49314
rect 72626 49144 73194 49314
rect 73362 49144 73930 49314
rect 74098 49144 74666 49314
rect 74834 49144 75402 49314
rect 75570 49144 76138 49314
rect 76306 49144 76874 49314
rect 77042 49144 77610 49314
rect 77778 49144 78346 49314
rect 78514 49144 79082 49314
rect 79250 49144 79818 49314
rect 79986 49144 80554 49314
rect 80722 49144 81290 49314
rect 81458 49144 82026 49314
rect 82194 49144 82762 49314
rect 82930 49144 83498 49314
rect 83666 49144 84234 49314
rect 84402 49144 84970 49314
rect 85138 49144 85706 49314
rect 85874 49144 86442 49314
rect 86610 49144 88392 49314
rect 1400 856 88392 49144
rect 1400 410 5114 856
rect 5282 410 5666 856
rect 5834 410 6218 856
rect 6386 410 6770 856
rect 6938 410 7322 856
rect 7490 410 7874 856
rect 8042 410 8426 856
rect 8594 410 8978 856
rect 9146 410 9530 856
rect 9698 410 10082 856
rect 10250 410 10634 856
rect 10802 410 11186 856
rect 11354 410 11738 856
rect 11906 410 12290 856
rect 12458 410 12842 856
rect 13010 410 13394 856
rect 13562 410 13946 856
rect 14114 410 14498 856
rect 14666 410 15050 856
rect 15218 410 15602 856
rect 15770 410 16154 856
rect 16322 410 16706 856
rect 16874 410 17258 856
rect 17426 410 17810 856
rect 17978 410 18362 856
rect 18530 410 18914 856
rect 19082 410 19466 856
rect 19634 410 20018 856
rect 20186 410 20570 856
rect 20738 410 21122 856
rect 21290 410 21674 856
rect 21842 410 22226 856
rect 22394 410 22778 856
rect 22946 410 23330 856
rect 23498 410 23882 856
rect 24050 410 24434 856
rect 24602 410 24986 856
rect 25154 410 25538 856
rect 25706 410 26090 856
rect 26258 410 26642 856
rect 26810 410 27194 856
rect 27362 410 27746 856
rect 27914 410 28298 856
rect 28466 410 28850 856
rect 29018 410 29402 856
rect 29570 410 29954 856
rect 30122 410 30506 856
rect 30674 410 31058 856
rect 31226 410 31610 856
rect 31778 410 32162 856
rect 32330 410 32714 856
rect 32882 410 33266 856
rect 33434 410 33818 856
rect 33986 410 34370 856
rect 34538 410 34922 856
rect 35090 410 35474 856
rect 35642 410 36026 856
rect 36194 410 36578 856
rect 36746 410 37130 856
rect 37298 410 37682 856
rect 37850 410 38234 856
rect 38402 410 38786 856
rect 38954 410 39338 856
rect 39506 410 39890 856
rect 40058 410 40442 856
rect 40610 410 40994 856
rect 41162 410 41546 856
rect 41714 410 42098 856
rect 42266 410 42650 856
rect 42818 410 43202 856
rect 43370 410 43754 856
rect 43922 410 44306 856
rect 44474 410 44858 856
rect 45026 410 45410 856
rect 45578 410 45962 856
rect 46130 410 46514 856
rect 46682 410 47066 856
rect 47234 410 47618 856
rect 47786 410 48170 856
rect 48338 410 48722 856
rect 48890 410 49274 856
rect 49442 410 49826 856
rect 49994 410 50378 856
rect 50546 410 50930 856
rect 51098 410 51482 856
rect 51650 410 52034 856
rect 52202 410 52586 856
rect 52754 410 53138 856
rect 53306 410 53690 856
rect 53858 410 54242 856
rect 54410 410 54794 856
rect 54962 410 55346 856
rect 55514 410 55898 856
rect 56066 410 56450 856
rect 56618 410 57002 856
rect 57170 410 57554 856
rect 57722 410 58106 856
rect 58274 410 58658 856
rect 58826 410 59210 856
rect 59378 410 59762 856
rect 59930 410 60314 856
rect 60482 410 60866 856
rect 61034 410 61418 856
rect 61586 410 61970 856
rect 62138 410 62522 856
rect 62690 410 63074 856
rect 63242 410 63626 856
rect 63794 410 64178 856
rect 64346 410 64730 856
rect 64898 410 65282 856
rect 65450 410 65834 856
rect 66002 410 66386 856
rect 66554 410 66938 856
rect 67106 410 67490 856
rect 67658 410 68042 856
rect 68210 410 68594 856
rect 68762 410 69146 856
rect 69314 410 69698 856
rect 69866 410 70250 856
rect 70418 410 70802 856
rect 70970 410 71354 856
rect 71522 410 71906 856
rect 72074 410 72458 856
rect 72626 410 73010 856
rect 73178 410 73562 856
rect 73730 410 74114 856
rect 74282 410 74666 856
rect 74834 410 75218 856
rect 75386 410 75770 856
rect 75938 410 76322 856
rect 76490 410 76874 856
rect 77042 410 77426 856
rect 77594 410 77978 856
rect 78146 410 78530 856
rect 78698 410 79082 856
rect 79250 410 79634 856
rect 79802 410 80186 856
rect 80354 410 80738 856
rect 80906 410 81290 856
rect 81458 410 81842 856
rect 82010 410 82394 856
rect 82562 410 82946 856
rect 83114 410 83498 856
rect 83666 410 84050 856
rect 84218 410 84602 856
rect 84770 410 88392 856
<< metal3 >>
rect 0 47200 800 47320
rect 0 46112 800 46232
rect 0 45024 800 45144
rect 0 43936 800 44056
rect 0 42848 800 42968
rect 0 41760 800 41880
rect 0 40672 800 40792
rect 0 39584 800 39704
rect 0 38496 800 38616
rect 0 37408 800 37528
rect 0 36320 800 36440
rect 0 35232 800 35352
rect 0 34144 800 34264
rect 0 33056 800 33176
rect 0 31968 800 32088
rect 0 30880 800 31000
rect 0 29792 800 29912
rect 0 28704 800 28824
rect 0 27616 800 27736
rect 0 26528 800 26648
rect 0 25440 800 25560
rect 0 24352 800 24472
rect 0 23264 800 23384
rect 0 22176 800 22296
rect 0 21088 800 21208
rect 0 20000 800 20120
rect 0 18912 800 19032
rect 0 17824 800 17944
rect 0 16736 800 16856
rect 0 15648 800 15768
rect 0 14560 800 14680
rect 0 13472 800 13592
rect 0 12384 800 12504
rect 0 11296 800 11416
rect 0 10208 800 10328
rect 0 9120 800 9240
rect 0 8032 800 8152
rect 0 6944 800 7064
rect 0 5856 800 5976
rect 0 4768 800 4888
rect 0 3680 800 3800
rect 0 2592 800 2712
<< obsm3 >>
rect 880 47120 88215 47361
rect 800 46312 88215 47120
rect 880 46032 88215 46312
rect 800 45224 88215 46032
rect 880 44944 88215 45224
rect 800 44136 88215 44944
rect 880 43856 88215 44136
rect 800 43048 88215 43856
rect 880 42768 88215 43048
rect 800 41960 88215 42768
rect 880 41680 88215 41960
rect 800 40872 88215 41680
rect 880 40592 88215 40872
rect 800 39784 88215 40592
rect 880 39504 88215 39784
rect 800 38696 88215 39504
rect 880 38416 88215 38696
rect 800 37608 88215 38416
rect 880 37328 88215 37608
rect 800 36520 88215 37328
rect 880 36240 88215 36520
rect 800 35432 88215 36240
rect 880 35152 88215 35432
rect 800 34344 88215 35152
rect 880 34064 88215 34344
rect 800 33256 88215 34064
rect 880 32976 88215 33256
rect 800 32168 88215 32976
rect 880 31888 88215 32168
rect 800 31080 88215 31888
rect 880 30800 88215 31080
rect 800 29992 88215 30800
rect 880 29712 88215 29992
rect 800 28904 88215 29712
rect 880 28624 88215 28904
rect 800 27816 88215 28624
rect 880 27536 88215 27816
rect 800 26728 88215 27536
rect 880 26448 88215 26728
rect 800 25640 88215 26448
rect 880 25360 88215 25640
rect 800 24552 88215 25360
rect 880 24272 88215 24552
rect 800 23464 88215 24272
rect 880 23184 88215 23464
rect 800 22376 88215 23184
rect 880 22096 88215 22376
rect 800 21288 88215 22096
rect 880 21008 88215 21288
rect 800 20200 88215 21008
rect 880 19920 88215 20200
rect 800 19112 88215 19920
rect 880 18832 88215 19112
rect 800 18024 88215 18832
rect 880 17744 88215 18024
rect 800 16936 88215 17744
rect 880 16656 88215 16936
rect 800 15848 88215 16656
rect 880 15568 88215 15848
rect 800 14760 88215 15568
rect 880 14480 88215 14760
rect 800 13672 88215 14480
rect 880 13392 88215 13672
rect 800 12584 88215 13392
rect 880 12304 88215 12584
rect 800 11496 88215 12304
rect 880 11216 88215 11496
rect 800 10408 88215 11216
rect 880 10128 88215 10408
rect 800 9320 88215 10128
rect 880 9040 88215 9320
rect 800 8232 88215 9040
rect 880 7952 88215 8232
rect 800 7144 88215 7952
rect 880 6864 88215 7144
rect 800 6056 88215 6864
rect 880 5776 88215 6056
rect 800 4968 88215 5776
rect 880 4688 88215 4968
rect 800 3880 88215 4688
rect 880 3600 88215 3880
rect 800 2792 88215 3600
rect 880 2512 88215 2792
rect 800 1395 88215 2512
<< metal4 >>
rect 4208 2128 4528 47376
rect 19568 2128 19888 47376
rect 34928 2128 35248 47376
rect 50288 2128 50608 47376
rect 65648 2128 65968 47376
rect 81008 2128 81328 47376
<< obsm4 >>
rect 4659 3571 19488 45661
rect 19968 3571 34848 45661
rect 35328 3571 50208 45661
rect 50688 3571 65568 45661
rect 66048 3571 78509 45661
<< labels >>
rlabel metal2 s 3330 49200 3386 50000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 25410 49200 25466 50000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 27618 49200 27674 50000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 29826 49200 29882 50000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 32034 49200 32090 50000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 34242 49200 34298 50000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 36450 49200 36506 50000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 38658 49200 38714 50000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 40866 49200 40922 50000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 43074 49200 43130 50000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 45282 49200 45338 50000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 5538 49200 5594 50000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 47490 49200 47546 50000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 49698 49200 49754 50000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 51906 49200 51962 50000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 54114 49200 54170 50000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 56322 49200 56378 50000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 58530 49200 58586 50000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 60738 49200 60794 50000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 62946 49200 63002 50000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 65154 49200 65210 50000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 67362 49200 67418 50000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 7746 49200 7802 50000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 69570 49200 69626 50000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 71778 49200 71834 50000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 73986 49200 74042 50000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 76194 49200 76250 50000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 78402 49200 78458 50000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 80610 49200 80666 50000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 82818 49200 82874 50000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 85026 49200 85082 50000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 9954 49200 10010 50000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 12162 49200 12218 50000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 14370 49200 14426 50000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 16578 49200 16634 50000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 18786 49200 18842 50000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 20994 49200 21050 50000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 23202 49200 23258 50000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 4066 49200 4122 50000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 26146 49200 26202 50000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 28354 49200 28410 50000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 30562 49200 30618 50000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 32770 49200 32826 50000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 34978 49200 35034 50000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 37186 49200 37242 50000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 39394 49200 39450 50000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 41602 49200 41658 50000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 43810 49200 43866 50000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 46018 49200 46074 50000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 6274 49200 6330 50000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 48226 49200 48282 50000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 50434 49200 50490 50000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 52642 49200 52698 50000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 54850 49200 54906 50000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 57058 49200 57114 50000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 59266 49200 59322 50000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 61474 49200 61530 50000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 63682 49200 63738 50000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 65890 49200 65946 50000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 68098 49200 68154 50000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 8482 49200 8538 50000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 70306 49200 70362 50000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 72514 49200 72570 50000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 74722 49200 74778 50000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 76930 49200 76986 50000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 79138 49200 79194 50000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 81346 49200 81402 50000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 83554 49200 83610 50000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 85762 49200 85818 50000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 10690 49200 10746 50000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 12898 49200 12954 50000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 15106 49200 15162 50000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 17314 49200 17370 50000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 19522 49200 19578 50000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 21730 49200 21786 50000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 23938 49200 23994 50000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 4802 49200 4858 50000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 26882 49200 26938 50000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 29090 49200 29146 50000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 31298 49200 31354 50000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 33506 49200 33562 50000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 35714 49200 35770 50000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 37922 49200 37978 50000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 40130 49200 40186 50000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 42338 49200 42394 50000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 44546 49200 44602 50000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 46754 49200 46810 50000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 7010 49200 7066 50000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 48962 49200 49018 50000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 51170 49200 51226 50000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 53378 49200 53434 50000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 55586 49200 55642 50000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 57794 49200 57850 50000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 60002 49200 60058 50000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 62210 49200 62266 50000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 64418 49200 64474 50000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 66626 49200 66682 50000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 68834 49200 68890 50000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 9218 49200 9274 50000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 71042 49200 71098 50000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 73250 49200 73306 50000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 75458 49200 75514 50000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 77666 49200 77722 50000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 79874 49200 79930 50000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 82082 49200 82138 50000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 84290 49200 84346 50000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 86498 49200 86554 50000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 11426 49200 11482 50000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 13634 49200 13690 50000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 15842 49200 15898 50000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 18050 49200 18106 50000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 20258 49200 20314 50000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 22466 49200 22522 50000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 24674 49200 24730 50000 6 io_out[9]
port 114 nsew signal output
rlabel metal3 s 0 3680 800 3800 6 oram_addr[0]
port 115 nsew signal output
rlabel metal3 s 0 5856 800 5976 6 oram_addr[1]
port 116 nsew signal output
rlabel metal3 s 0 8032 800 8152 6 oram_addr[2]
port 117 nsew signal output
rlabel metal3 s 0 10208 800 10328 6 oram_addr[3]
port 118 nsew signal output
rlabel metal3 s 0 12384 800 12504 6 oram_addr[4]
port 119 nsew signal output
rlabel metal3 s 0 14560 800 14680 6 oram_addr[5]
port 120 nsew signal output
rlabel metal3 s 0 16736 800 16856 6 oram_addr[6]
port 121 nsew signal output
rlabel metal3 s 0 18912 800 19032 6 oram_addr[7]
port 122 nsew signal output
rlabel metal3 s 0 21088 800 21208 6 oram_addr[8]
port 123 nsew signal output
rlabel metal3 s 0 2592 800 2712 6 oram_csb
port 124 nsew signal output
rlabel metal3 s 0 4768 800 4888 6 oram_value[0]
port 125 nsew signal input
rlabel metal3 s 0 24352 800 24472 6 oram_value[10]
port 126 nsew signal input
rlabel metal3 s 0 25440 800 25560 6 oram_value[11]
port 127 nsew signal input
rlabel metal3 s 0 26528 800 26648 6 oram_value[12]
port 128 nsew signal input
rlabel metal3 s 0 27616 800 27736 6 oram_value[13]
port 129 nsew signal input
rlabel metal3 s 0 28704 800 28824 6 oram_value[14]
port 130 nsew signal input
rlabel metal3 s 0 29792 800 29912 6 oram_value[15]
port 131 nsew signal input
rlabel metal3 s 0 30880 800 31000 6 oram_value[16]
port 132 nsew signal input
rlabel metal3 s 0 31968 800 32088 6 oram_value[17]
port 133 nsew signal input
rlabel metal3 s 0 33056 800 33176 6 oram_value[18]
port 134 nsew signal input
rlabel metal3 s 0 34144 800 34264 6 oram_value[19]
port 135 nsew signal input
rlabel metal3 s 0 6944 800 7064 6 oram_value[1]
port 136 nsew signal input
rlabel metal3 s 0 35232 800 35352 6 oram_value[20]
port 137 nsew signal input
rlabel metal3 s 0 36320 800 36440 6 oram_value[21]
port 138 nsew signal input
rlabel metal3 s 0 37408 800 37528 6 oram_value[22]
port 139 nsew signal input
rlabel metal3 s 0 38496 800 38616 6 oram_value[23]
port 140 nsew signal input
rlabel metal3 s 0 39584 800 39704 6 oram_value[24]
port 141 nsew signal input
rlabel metal3 s 0 40672 800 40792 6 oram_value[25]
port 142 nsew signal input
rlabel metal3 s 0 41760 800 41880 6 oram_value[26]
port 143 nsew signal input
rlabel metal3 s 0 42848 800 42968 6 oram_value[27]
port 144 nsew signal input
rlabel metal3 s 0 43936 800 44056 6 oram_value[28]
port 145 nsew signal input
rlabel metal3 s 0 45024 800 45144 6 oram_value[29]
port 146 nsew signal input
rlabel metal3 s 0 9120 800 9240 6 oram_value[2]
port 147 nsew signal input
rlabel metal3 s 0 46112 800 46232 6 oram_value[30]
port 148 nsew signal input
rlabel metal3 s 0 47200 800 47320 6 oram_value[31]
port 149 nsew signal input
rlabel metal3 s 0 11296 800 11416 6 oram_value[3]
port 150 nsew signal input
rlabel metal3 s 0 13472 800 13592 6 oram_value[4]
port 151 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 oram_value[5]
port 152 nsew signal input
rlabel metal3 s 0 17824 800 17944 6 oram_value[6]
port 153 nsew signal input
rlabel metal3 s 0 20000 800 20120 6 oram_value[7]
port 154 nsew signal input
rlabel metal3 s 0 22176 800 22296 6 oram_value[8]
port 155 nsew signal input
rlabel metal3 s 0 23264 800 23384 6 oram_value[9]
port 156 nsew signal input
rlabel metal2 s 62578 0 62634 800 6 ram_adrb[0]
port 157 nsew signal output
rlabel metal2 s 63682 0 63738 800 6 ram_adrb[1]
port 158 nsew signal output
rlabel metal2 s 64786 0 64842 800 6 ram_adrb[2]
port 159 nsew signal output
rlabel metal2 s 65890 0 65946 800 6 ram_adrb[3]
port 160 nsew signal output
rlabel metal2 s 66994 0 67050 800 6 ram_adrb[4]
port 161 nsew signal output
rlabel metal2 s 68098 0 68154 800 6 ram_adrb[5]
port 162 nsew signal output
rlabel metal2 s 69202 0 69258 800 6 ram_adrb[6]
port 163 nsew signal output
rlabel metal2 s 70306 0 70362 800 6 ram_adrb[7]
port 164 nsew signal output
rlabel metal2 s 71410 0 71466 800 6 ram_adrb[8]
port 165 nsew signal output
rlabel metal2 s 61474 0 61530 800 6 ram_csb
port 166 nsew signal output
rlabel metal2 s 63130 0 63186 800 6 ram_val[0]
port 167 nsew signal input
rlabel metal2 s 73066 0 73122 800 6 ram_val[10]
port 168 nsew signal input
rlabel metal2 s 73618 0 73674 800 6 ram_val[11]
port 169 nsew signal input
rlabel metal2 s 74170 0 74226 800 6 ram_val[12]
port 170 nsew signal input
rlabel metal2 s 74722 0 74778 800 6 ram_val[13]
port 171 nsew signal input
rlabel metal2 s 75274 0 75330 800 6 ram_val[14]
port 172 nsew signal input
rlabel metal2 s 75826 0 75882 800 6 ram_val[15]
port 173 nsew signal input
rlabel metal2 s 76378 0 76434 800 6 ram_val[16]
port 174 nsew signal input
rlabel metal2 s 76930 0 76986 800 6 ram_val[17]
port 175 nsew signal input
rlabel metal2 s 77482 0 77538 800 6 ram_val[18]
port 176 nsew signal input
rlabel metal2 s 78034 0 78090 800 6 ram_val[19]
port 177 nsew signal input
rlabel metal2 s 64234 0 64290 800 6 ram_val[1]
port 178 nsew signal input
rlabel metal2 s 78586 0 78642 800 6 ram_val[20]
port 179 nsew signal input
rlabel metal2 s 79138 0 79194 800 6 ram_val[21]
port 180 nsew signal input
rlabel metal2 s 79690 0 79746 800 6 ram_val[22]
port 181 nsew signal input
rlabel metal2 s 80242 0 80298 800 6 ram_val[23]
port 182 nsew signal input
rlabel metal2 s 80794 0 80850 800 6 ram_val[24]
port 183 nsew signal input
rlabel metal2 s 81346 0 81402 800 6 ram_val[25]
port 184 nsew signal input
rlabel metal2 s 81898 0 81954 800 6 ram_val[26]
port 185 nsew signal input
rlabel metal2 s 82450 0 82506 800 6 ram_val[27]
port 186 nsew signal input
rlabel metal2 s 83002 0 83058 800 6 ram_val[28]
port 187 nsew signal input
rlabel metal2 s 83554 0 83610 800 6 ram_val[29]
port 188 nsew signal input
rlabel metal2 s 65338 0 65394 800 6 ram_val[2]
port 189 nsew signal input
rlabel metal2 s 84106 0 84162 800 6 ram_val[30]
port 190 nsew signal input
rlabel metal2 s 84658 0 84714 800 6 ram_val[31]
port 191 nsew signal input
rlabel metal2 s 66442 0 66498 800 6 ram_val[3]
port 192 nsew signal input
rlabel metal2 s 67546 0 67602 800 6 ram_val[4]
port 193 nsew signal input
rlabel metal2 s 68650 0 68706 800 6 ram_val[5]
port 194 nsew signal input
rlabel metal2 s 69754 0 69810 800 6 ram_val[6]
port 195 nsew signal input
rlabel metal2 s 70858 0 70914 800 6 ram_val[7]
port 196 nsew signal input
rlabel metal2 s 71962 0 72018 800 6 ram_val[8]
port 197 nsew signal input
rlabel metal2 s 72514 0 72570 800 6 ram_val[9]
port 198 nsew signal input
rlabel metal2 s 62026 0 62082 800 6 ram_web
port 199 nsew signal output
rlabel metal4 s 4208 2128 4528 47376 6 vccd1
port 200 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 47376 6 vccd1
port 200 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 47376 6 vccd1
port 200 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 47376 6 vssd1
port 201 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 47376 6 vssd1
port 201 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 47376 6 vssd1
port 201 nsew ground bidirectional
rlabel metal2 s 5170 0 5226 800 6 wb_clk_i
port 202 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 wb_rst_i
port 203 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 wbs_ack_o
port 204 nsew signal output
rlabel metal2 s 8482 0 8538 800 6 wbs_adr_i[0]
port 205 nsew signal input
rlabel metal2 s 25042 0 25098 800 6 wbs_adr_i[10]
port 206 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 wbs_adr_i[11]
port 207 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 wbs_adr_i[12]
port 208 nsew signal input
rlabel metal2 s 30010 0 30066 800 6 wbs_adr_i[13]
port 209 nsew signal input
rlabel metal2 s 31666 0 31722 800 6 wbs_adr_i[14]
port 210 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 wbs_adr_i[15]
port 211 nsew signal input
rlabel metal2 s 34978 0 35034 800 6 wbs_adr_i[16]
port 212 nsew signal input
rlabel metal2 s 36634 0 36690 800 6 wbs_adr_i[17]
port 213 nsew signal input
rlabel metal2 s 38290 0 38346 800 6 wbs_adr_i[18]
port 214 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 wbs_adr_i[19]
port 215 nsew signal input
rlabel metal2 s 10138 0 10194 800 6 wbs_adr_i[1]
port 216 nsew signal input
rlabel metal2 s 41602 0 41658 800 6 wbs_adr_i[20]
port 217 nsew signal input
rlabel metal2 s 43258 0 43314 800 6 wbs_adr_i[21]
port 218 nsew signal input
rlabel metal2 s 44914 0 44970 800 6 wbs_adr_i[22]
port 219 nsew signal input
rlabel metal2 s 46570 0 46626 800 6 wbs_adr_i[23]
port 220 nsew signal input
rlabel metal2 s 48226 0 48282 800 6 wbs_adr_i[24]
port 221 nsew signal input
rlabel metal2 s 49882 0 49938 800 6 wbs_adr_i[25]
port 222 nsew signal input
rlabel metal2 s 51538 0 51594 800 6 wbs_adr_i[26]
port 223 nsew signal input
rlabel metal2 s 53194 0 53250 800 6 wbs_adr_i[27]
port 224 nsew signal input
rlabel metal2 s 54850 0 54906 800 6 wbs_adr_i[28]
port 225 nsew signal input
rlabel metal2 s 56506 0 56562 800 6 wbs_adr_i[29]
port 226 nsew signal input
rlabel metal2 s 11794 0 11850 800 6 wbs_adr_i[2]
port 227 nsew signal input
rlabel metal2 s 58162 0 58218 800 6 wbs_adr_i[30]
port 228 nsew signal input
rlabel metal2 s 59818 0 59874 800 6 wbs_adr_i[31]
port 229 nsew signal input
rlabel metal2 s 13450 0 13506 800 6 wbs_adr_i[3]
port 230 nsew signal input
rlabel metal2 s 15106 0 15162 800 6 wbs_adr_i[4]
port 231 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 wbs_adr_i[5]
port 232 nsew signal input
rlabel metal2 s 18418 0 18474 800 6 wbs_adr_i[6]
port 233 nsew signal input
rlabel metal2 s 20074 0 20130 800 6 wbs_adr_i[7]
port 234 nsew signal input
rlabel metal2 s 21730 0 21786 800 6 wbs_adr_i[8]
port 235 nsew signal input
rlabel metal2 s 23386 0 23442 800 6 wbs_adr_i[9]
port 236 nsew signal input
rlabel metal2 s 6826 0 6882 800 6 wbs_cyc_i
port 237 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 wbs_dat_i[0]
port 238 nsew signal input
rlabel metal2 s 25594 0 25650 800 6 wbs_dat_i[10]
port 239 nsew signal input
rlabel metal2 s 27250 0 27306 800 6 wbs_dat_i[11]
port 240 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 wbs_dat_i[12]
port 241 nsew signal input
rlabel metal2 s 30562 0 30618 800 6 wbs_dat_i[13]
port 242 nsew signal input
rlabel metal2 s 32218 0 32274 800 6 wbs_dat_i[14]
port 243 nsew signal input
rlabel metal2 s 33874 0 33930 800 6 wbs_dat_i[15]
port 244 nsew signal input
rlabel metal2 s 35530 0 35586 800 6 wbs_dat_i[16]
port 245 nsew signal input
rlabel metal2 s 37186 0 37242 800 6 wbs_dat_i[17]
port 246 nsew signal input
rlabel metal2 s 38842 0 38898 800 6 wbs_dat_i[18]
port 247 nsew signal input
rlabel metal2 s 40498 0 40554 800 6 wbs_dat_i[19]
port 248 nsew signal input
rlabel metal2 s 10690 0 10746 800 6 wbs_dat_i[1]
port 249 nsew signal input
rlabel metal2 s 42154 0 42210 800 6 wbs_dat_i[20]
port 250 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 wbs_dat_i[21]
port 251 nsew signal input
rlabel metal2 s 45466 0 45522 800 6 wbs_dat_i[22]
port 252 nsew signal input
rlabel metal2 s 47122 0 47178 800 6 wbs_dat_i[23]
port 253 nsew signal input
rlabel metal2 s 48778 0 48834 800 6 wbs_dat_i[24]
port 254 nsew signal input
rlabel metal2 s 50434 0 50490 800 6 wbs_dat_i[25]
port 255 nsew signal input
rlabel metal2 s 52090 0 52146 800 6 wbs_dat_i[26]
port 256 nsew signal input
rlabel metal2 s 53746 0 53802 800 6 wbs_dat_i[27]
port 257 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 wbs_dat_i[28]
port 258 nsew signal input
rlabel metal2 s 57058 0 57114 800 6 wbs_dat_i[29]
port 259 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 wbs_dat_i[2]
port 260 nsew signal input
rlabel metal2 s 58714 0 58770 800 6 wbs_dat_i[30]
port 261 nsew signal input
rlabel metal2 s 60370 0 60426 800 6 wbs_dat_i[31]
port 262 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 wbs_dat_i[3]
port 263 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 wbs_dat_i[4]
port 264 nsew signal input
rlabel metal2 s 17314 0 17370 800 6 wbs_dat_i[5]
port 265 nsew signal input
rlabel metal2 s 18970 0 19026 800 6 wbs_dat_i[6]
port 266 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 wbs_dat_i[7]
port 267 nsew signal input
rlabel metal2 s 22282 0 22338 800 6 wbs_dat_i[8]
port 268 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 wbs_dat_i[9]
port 269 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 wbs_dat_o[0]
port 270 nsew signal output
rlabel metal2 s 26146 0 26202 800 6 wbs_dat_o[10]
port 271 nsew signal output
rlabel metal2 s 27802 0 27858 800 6 wbs_dat_o[11]
port 272 nsew signal output
rlabel metal2 s 29458 0 29514 800 6 wbs_dat_o[12]
port 273 nsew signal output
rlabel metal2 s 31114 0 31170 800 6 wbs_dat_o[13]
port 274 nsew signal output
rlabel metal2 s 32770 0 32826 800 6 wbs_dat_o[14]
port 275 nsew signal output
rlabel metal2 s 34426 0 34482 800 6 wbs_dat_o[15]
port 276 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 wbs_dat_o[16]
port 277 nsew signal output
rlabel metal2 s 37738 0 37794 800 6 wbs_dat_o[17]
port 278 nsew signal output
rlabel metal2 s 39394 0 39450 800 6 wbs_dat_o[18]
port 279 nsew signal output
rlabel metal2 s 41050 0 41106 800 6 wbs_dat_o[19]
port 280 nsew signal output
rlabel metal2 s 11242 0 11298 800 6 wbs_dat_o[1]
port 281 nsew signal output
rlabel metal2 s 42706 0 42762 800 6 wbs_dat_o[20]
port 282 nsew signal output
rlabel metal2 s 44362 0 44418 800 6 wbs_dat_o[21]
port 283 nsew signal output
rlabel metal2 s 46018 0 46074 800 6 wbs_dat_o[22]
port 284 nsew signal output
rlabel metal2 s 47674 0 47730 800 6 wbs_dat_o[23]
port 285 nsew signal output
rlabel metal2 s 49330 0 49386 800 6 wbs_dat_o[24]
port 286 nsew signal output
rlabel metal2 s 50986 0 51042 800 6 wbs_dat_o[25]
port 287 nsew signal output
rlabel metal2 s 52642 0 52698 800 6 wbs_dat_o[26]
port 288 nsew signal output
rlabel metal2 s 54298 0 54354 800 6 wbs_dat_o[27]
port 289 nsew signal output
rlabel metal2 s 55954 0 56010 800 6 wbs_dat_o[28]
port 290 nsew signal output
rlabel metal2 s 57610 0 57666 800 6 wbs_dat_o[29]
port 291 nsew signal output
rlabel metal2 s 12898 0 12954 800 6 wbs_dat_o[2]
port 292 nsew signal output
rlabel metal2 s 59266 0 59322 800 6 wbs_dat_o[30]
port 293 nsew signal output
rlabel metal2 s 60922 0 60978 800 6 wbs_dat_o[31]
port 294 nsew signal output
rlabel metal2 s 14554 0 14610 800 6 wbs_dat_o[3]
port 295 nsew signal output
rlabel metal2 s 16210 0 16266 800 6 wbs_dat_o[4]
port 296 nsew signal output
rlabel metal2 s 17866 0 17922 800 6 wbs_dat_o[5]
port 297 nsew signal output
rlabel metal2 s 19522 0 19578 800 6 wbs_dat_o[6]
port 298 nsew signal output
rlabel metal2 s 21178 0 21234 800 6 wbs_dat_o[7]
port 299 nsew signal output
rlabel metal2 s 22834 0 22890 800 6 wbs_dat_o[8]
port 300 nsew signal output
rlabel metal2 s 24490 0 24546 800 6 wbs_dat_o[9]
port 301 nsew signal output
rlabel metal2 s 7378 0 7434 800 6 wbs_stb_i
port 302 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 wbs_we_i
port 303 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 90000 50000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 12173056
string GDS_FILE /home/lucah/Videos/mpw-8-as1x00/openlane/wrapped_tms1x00/runs/22_12_22_09_38/results/signoff/wrapped_tms1x00.magic.gds
string GDS_START 662648
<< end >>

