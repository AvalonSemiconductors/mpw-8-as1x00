// This is the unpowered netlist.
module tms1x00_ram (clk,
    wen,
    r_val,
    ram_addr,
    w_val);
 input clk;
 input wen;
 output [3:0] r_val;
 input [6:0] ram_addr;
 input [3:0] w_val;

 wire \RAM[0][0] ;
 wire \RAM[0][1] ;
 wire \RAM[0][2] ;
 wire \RAM[0][3] ;
 wire \RAM[100][0] ;
 wire \RAM[100][1] ;
 wire \RAM[100][2] ;
 wire \RAM[100][3] ;
 wire \RAM[101][0] ;
 wire \RAM[101][1] ;
 wire \RAM[101][2] ;
 wire \RAM[101][3] ;
 wire \RAM[102][0] ;
 wire \RAM[102][1] ;
 wire \RAM[102][2] ;
 wire \RAM[102][3] ;
 wire \RAM[103][0] ;
 wire \RAM[103][1] ;
 wire \RAM[103][2] ;
 wire \RAM[103][3] ;
 wire \RAM[104][0] ;
 wire \RAM[104][1] ;
 wire \RAM[104][2] ;
 wire \RAM[104][3] ;
 wire \RAM[105][0] ;
 wire \RAM[105][1] ;
 wire \RAM[105][2] ;
 wire \RAM[105][3] ;
 wire \RAM[106][0] ;
 wire \RAM[106][1] ;
 wire \RAM[106][2] ;
 wire \RAM[106][3] ;
 wire \RAM[107][0] ;
 wire \RAM[107][1] ;
 wire \RAM[107][2] ;
 wire \RAM[107][3] ;
 wire \RAM[108][0] ;
 wire \RAM[108][1] ;
 wire \RAM[108][2] ;
 wire \RAM[108][3] ;
 wire \RAM[109][0] ;
 wire \RAM[109][1] ;
 wire \RAM[109][2] ;
 wire \RAM[109][3] ;
 wire \RAM[10][0] ;
 wire \RAM[10][1] ;
 wire \RAM[10][2] ;
 wire \RAM[10][3] ;
 wire \RAM[110][0] ;
 wire \RAM[110][1] ;
 wire \RAM[110][2] ;
 wire \RAM[110][3] ;
 wire \RAM[111][0] ;
 wire \RAM[111][1] ;
 wire \RAM[111][2] ;
 wire \RAM[111][3] ;
 wire \RAM[112][0] ;
 wire \RAM[112][1] ;
 wire \RAM[112][2] ;
 wire \RAM[112][3] ;
 wire \RAM[113][0] ;
 wire \RAM[113][1] ;
 wire \RAM[113][2] ;
 wire \RAM[113][3] ;
 wire \RAM[114][0] ;
 wire \RAM[114][1] ;
 wire \RAM[114][2] ;
 wire \RAM[114][3] ;
 wire \RAM[115][0] ;
 wire \RAM[115][1] ;
 wire \RAM[115][2] ;
 wire \RAM[115][3] ;
 wire \RAM[116][0] ;
 wire \RAM[116][1] ;
 wire \RAM[116][2] ;
 wire \RAM[116][3] ;
 wire \RAM[117][0] ;
 wire \RAM[117][1] ;
 wire \RAM[117][2] ;
 wire \RAM[117][3] ;
 wire \RAM[118][0] ;
 wire \RAM[118][1] ;
 wire \RAM[118][2] ;
 wire \RAM[118][3] ;
 wire \RAM[119][0] ;
 wire \RAM[119][1] ;
 wire \RAM[119][2] ;
 wire \RAM[119][3] ;
 wire \RAM[11][0] ;
 wire \RAM[11][1] ;
 wire \RAM[11][2] ;
 wire \RAM[11][3] ;
 wire \RAM[120][0] ;
 wire \RAM[120][1] ;
 wire \RAM[120][2] ;
 wire \RAM[120][3] ;
 wire \RAM[121][0] ;
 wire \RAM[121][1] ;
 wire \RAM[121][2] ;
 wire \RAM[121][3] ;
 wire \RAM[122][0] ;
 wire \RAM[122][1] ;
 wire \RAM[122][2] ;
 wire \RAM[122][3] ;
 wire \RAM[123][0] ;
 wire \RAM[123][1] ;
 wire \RAM[123][2] ;
 wire \RAM[123][3] ;
 wire \RAM[124][0] ;
 wire \RAM[124][1] ;
 wire \RAM[124][2] ;
 wire \RAM[124][3] ;
 wire \RAM[125][0] ;
 wire \RAM[125][1] ;
 wire \RAM[125][2] ;
 wire \RAM[125][3] ;
 wire \RAM[126][0] ;
 wire \RAM[126][1] ;
 wire \RAM[126][2] ;
 wire \RAM[126][3] ;
 wire \RAM[127][0] ;
 wire \RAM[127][1] ;
 wire \RAM[127][2] ;
 wire \RAM[127][3] ;
 wire \RAM[12][0] ;
 wire \RAM[12][1] ;
 wire \RAM[12][2] ;
 wire \RAM[12][3] ;
 wire \RAM[13][0] ;
 wire \RAM[13][1] ;
 wire \RAM[13][2] ;
 wire \RAM[13][3] ;
 wire \RAM[14][0] ;
 wire \RAM[14][1] ;
 wire \RAM[14][2] ;
 wire \RAM[14][3] ;
 wire \RAM[15][0] ;
 wire \RAM[15][1] ;
 wire \RAM[15][2] ;
 wire \RAM[15][3] ;
 wire \RAM[16][0] ;
 wire \RAM[16][1] ;
 wire \RAM[16][2] ;
 wire \RAM[16][3] ;
 wire \RAM[17][0] ;
 wire \RAM[17][1] ;
 wire \RAM[17][2] ;
 wire \RAM[17][3] ;
 wire \RAM[18][0] ;
 wire \RAM[18][1] ;
 wire \RAM[18][2] ;
 wire \RAM[18][3] ;
 wire \RAM[19][0] ;
 wire \RAM[19][1] ;
 wire \RAM[19][2] ;
 wire \RAM[19][3] ;
 wire \RAM[1][0] ;
 wire \RAM[1][1] ;
 wire \RAM[1][2] ;
 wire \RAM[1][3] ;
 wire \RAM[20][0] ;
 wire \RAM[20][1] ;
 wire \RAM[20][2] ;
 wire \RAM[20][3] ;
 wire \RAM[21][0] ;
 wire \RAM[21][1] ;
 wire \RAM[21][2] ;
 wire \RAM[21][3] ;
 wire \RAM[22][0] ;
 wire \RAM[22][1] ;
 wire \RAM[22][2] ;
 wire \RAM[22][3] ;
 wire \RAM[23][0] ;
 wire \RAM[23][1] ;
 wire \RAM[23][2] ;
 wire \RAM[23][3] ;
 wire \RAM[24][0] ;
 wire \RAM[24][1] ;
 wire \RAM[24][2] ;
 wire \RAM[24][3] ;
 wire \RAM[25][0] ;
 wire \RAM[25][1] ;
 wire \RAM[25][2] ;
 wire \RAM[25][3] ;
 wire \RAM[26][0] ;
 wire \RAM[26][1] ;
 wire \RAM[26][2] ;
 wire \RAM[26][3] ;
 wire \RAM[27][0] ;
 wire \RAM[27][1] ;
 wire \RAM[27][2] ;
 wire \RAM[27][3] ;
 wire \RAM[28][0] ;
 wire \RAM[28][1] ;
 wire \RAM[28][2] ;
 wire \RAM[28][3] ;
 wire \RAM[29][0] ;
 wire \RAM[29][1] ;
 wire \RAM[29][2] ;
 wire \RAM[29][3] ;
 wire \RAM[2][0] ;
 wire \RAM[2][1] ;
 wire \RAM[2][2] ;
 wire \RAM[2][3] ;
 wire \RAM[30][0] ;
 wire \RAM[30][1] ;
 wire \RAM[30][2] ;
 wire \RAM[30][3] ;
 wire \RAM[31][0] ;
 wire \RAM[31][1] ;
 wire \RAM[31][2] ;
 wire \RAM[31][3] ;
 wire \RAM[32][0] ;
 wire \RAM[32][1] ;
 wire \RAM[32][2] ;
 wire \RAM[32][3] ;
 wire \RAM[33][0] ;
 wire \RAM[33][1] ;
 wire \RAM[33][2] ;
 wire \RAM[33][3] ;
 wire \RAM[34][0] ;
 wire \RAM[34][1] ;
 wire \RAM[34][2] ;
 wire \RAM[34][3] ;
 wire \RAM[35][0] ;
 wire \RAM[35][1] ;
 wire \RAM[35][2] ;
 wire \RAM[35][3] ;
 wire \RAM[36][0] ;
 wire \RAM[36][1] ;
 wire \RAM[36][2] ;
 wire \RAM[36][3] ;
 wire \RAM[37][0] ;
 wire \RAM[37][1] ;
 wire \RAM[37][2] ;
 wire \RAM[37][3] ;
 wire \RAM[38][0] ;
 wire \RAM[38][1] ;
 wire \RAM[38][2] ;
 wire \RAM[38][3] ;
 wire \RAM[39][0] ;
 wire \RAM[39][1] ;
 wire \RAM[39][2] ;
 wire \RAM[39][3] ;
 wire \RAM[3][0] ;
 wire \RAM[3][1] ;
 wire \RAM[3][2] ;
 wire \RAM[3][3] ;
 wire \RAM[40][0] ;
 wire \RAM[40][1] ;
 wire \RAM[40][2] ;
 wire \RAM[40][3] ;
 wire \RAM[41][0] ;
 wire \RAM[41][1] ;
 wire \RAM[41][2] ;
 wire \RAM[41][3] ;
 wire \RAM[42][0] ;
 wire \RAM[42][1] ;
 wire \RAM[42][2] ;
 wire \RAM[42][3] ;
 wire \RAM[43][0] ;
 wire \RAM[43][1] ;
 wire \RAM[43][2] ;
 wire \RAM[43][3] ;
 wire \RAM[44][0] ;
 wire \RAM[44][1] ;
 wire \RAM[44][2] ;
 wire \RAM[44][3] ;
 wire \RAM[45][0] ;
 wire \RAM[45][1] ;
 wire \RAM[45][2] ;
 wire \RAM[45][3] ;
 wire \RAM[46][0] ;
 wire \RAM[46][1] ;
 wire \RAM[46][2] ;
 wire \RAM[46][3] ;
 wire \RAM[47][0] ;
 wire \RAM[47][1] ;
 wire \RAM[47][2] ;
 wire \RAM[47][3] ;
 wire \RAM[48][0] ;
 wire \RAM[48][1] ;
 wire \RAM[48][2] ;
 wire \RAM[48][3] ;
 wire \RAM[49][0] ;
 wire \RAM[49][1] ;
 wire \RAM[49][2] ;
 wire \RAM[49][3] ;
 wire \RAM[4][0] ;
 wire \RAM[4][1] ;
 wire \RAM[4][2] ;
 wire \RAM[4][3] ;
 wire \RAM[50][0] ;
 wire \RAM[50][1] ;
 wire \RAM[50][2] ;
 wire \RAM[50][3] ;
 wire \RAM[51][0] ;
 wire \RAM[51][1] ;
 wire \RAM[51][2] ;
 wire \RAM[51][3] ;
 wire \RAM[52][0] ;
 wire \RAM[52][1] ;
 wire \RAM[52][2] ;
 wire \RAM[52][3] ;
 wire \RAM[53][0] ;
 wire \RAM[53][1] ;
 wire \RAM[53][2] ;
 wire \RAM[53][3] ;
 wire \RAM[54][0] ;
 wire \RAM[54][1] ;
 wire \RAM[54][2] ;
 wire \RAM[54][3] ;
 wire \RAM[55][0] ;
 wire \RAM[55][1] ;
 wire \RAM[55][2] ;
 wire \RAM[55][3] ;
 wire \RAM[56][0] ;
 wire \RAM[56][1] ;
 wire \RAM[56][2] ;
 wire \RAM[56][3] ;
 wire \RAM[57][0] ;
 wire \RAM[57][1] ;
 wire \RAM[57][2] ;
 wire \RAM[57][3] ;
 wire \RAM[58][0] ;
 wire \RAM[58][1] ;
 wire \RAM[58][2] ;
 wire \RAM[58][3] ;
 wire \RAM[59][0] ;
 wire \RAM[59][1] ;
 wire \RAM[59][2] ;
 wire \RAM[59][3] ;
 wire \RAM[5][0] ;
 wire \RAM[5][1] ;
 wire \RAM[5][2] ;
 wire \RAM[5][3] ;
 wire \RAM[60][0] ;
 wire \RAM[60][1] ;
 wire \RAM[60][2] ;
 wire \RAM[60][3] ;
 wire \RAM[61][0] ;
 wire \RAM[61][1] ;
 wire \RAM[61][2] ;
 wire \RAM[61][3] ;
 wire \RAM[62][0] ;
 wire \RAM[62][1] ;
 wire \RAM[62][2] ;
 wire \RAM[62][3] ;
 wire \RAM[63][0] ;
 wire \RAM[63][1] ;
 wire \RAM[63][2] ;
 wire \RAM[63][3] ;
 wire \RAM[64][0] ;
 wire \RAM[64][1] ;
 wire \RAM[64][2] ;
 wire \RAM[64][3] ;
 wire \RAM[65][0] ;
 wire \RAM[65][1] ;
 wire \RAM[65][2] ;
 wire \RAM[65][3] ;
 wire \RAM[66][0] ;
 wire \RAM[66][1] ;
 wire \RAM[66][2] ;
 wire \RAM[66][3] ;
 wire \RAM[67][0] ;
 wire \RAM[67][1] ;
 wire \RAM[67][2] ;
 wire \RAM[67][3] ;
 wire \RAM[68][0] ;
 wire \RAM[68][1] ;
 wire \RAM[68][2] ;
 wire \RAM[68][3] ;
 wire \RAM[69][0] ;
 wire \RAM[69][1] ;
 wire \RAM[69][2] ;
 wire \RAM[69][3] ;
 wire \RAM[6][0] ;
 wire \RAM[6][1] ;
 wire \RAM[6][2] ;
 wire \RAM[6][3] ;
 wire \RAM[70][0] ;
 wire \RAM[70][1] ;
 wire \RAM[70][2] ;
 wire \RAM[70][3] ;
 wire \RAM[71][0] ;
 wire \RAM[71][1] ;
 wire \RAM[71][2] ;
 wire \RAM[71][3] ;
 wire \RAM[72][0] ;
 wire \RAM[72][1] ;
 wire \RAM[72][2] ;
 wire \RAM[72][3] ;
 wire \RAM[73][0] ;
 wire \RAM[73][1] ;
 wire \RAM[73][2] ;
 wire \RAM[73][3] ;
 wire \RAM[74][0] ;
 wire \RAM[74][1] ;
 wire \RAM[74][2] ;
 wire \RAM[74][3] ;
 wire \RAM[75][0] ;
 wire \RAM[75][1] ;
 wire \RAM[75][2] ;
 wire \RAM[75][3] ;
 wire \RAM[76][0] ;
 wire \RAM[76][1] ;
 wire \RAM[76][2] ;
 wire \RAM[76][3] ;
 wire \RAM[77][0] ;
 wire \RAM[77][1] ;
 wire \RAM[77][2] ;
 wire \RAM[77][3] ;
 wire \RAM[78][0] ;
 wire \RAM[78][1] ;
 wire \RAM[78][2] ;
 wire \RAM[78][3] ;
 wire \RAM[79][0] ;
 wire \RAM[79][1] ;
 wire \RAM[79][2] ;
 wire \RAM[79][3] ;
 wire \RAM[7][0] ;
 wire \RAM[7][1] ;
 wire \RAM[7][2] ;
 wire \RAM[7][3] ;
 wire \RAM[80][0] ;
 wire \RAM[80][1] ;
 wire \RAM[80][2] ;
 wire \RAM[80][3] ;
 wire \RAM[81][0] ;
 wire \RAM[81][1] ;
 wire \RAM[81][2] ;
 wire \RAM[81][3] ;
 wire \RAM[82][0] ;
 wire \RAM[82][1] ;
 wire \RAM[82][2] ;
 wire \RAM[82][3] ;
 wire \RAM[83][0] ;
 wire \RAM[83][1] ;
 wire \RAM[83][2] ;
 wire \RAM[83][3] ;
 wire \RAM[84][0] ;
 wire \RAM[84][1] ;
 wire \RAM[84][2] ;
 wire \RAM[84][3] ;
 wire \RAM[85][0] ;
 wire \RAM[85][1] ;
 wire \RAM[85][2] ;
 wire \RAM[85][3] ;
 wire \RAM[86][0] ;
 wire \RAM[86][1] ;
 wire \RAM[86][2] ;
 wire \RAM[86][3] ;
 wire \RAM[87][0] ;
 wire \RAM[87][1] ;
 wire \RAM[87][2] ;
 wire \RAM[87][3] ;
 wire \RAM[88][0] ;
 wire \RAM[88][1] ;
 wire \RAM[88][2] ;
 wire \RAM[88][3] ;
 wire \RAM[89][0] ;
 wire \RAM[89][1] ;
 wire \RAM[89][2] ;
 wire \RAM[89][3] ;
 wire \RAM[8][0] ;
 wire \RAM[8][1] ;
 wire \RAM[8][2] ;
 wire \RAM[8][3] ;
 wire \RAM[90][0] ;
 wire \RAM[90][1] ;
 wire \RAM[90][2] ;
 wire \RAM[90][3] ;
 wire \RAM[91][0] ;
 wire \RAM[91][1] ;
 wire \RAM[91][2] ;
 wire \RAM[91][3] ;
 wire \RAM[92][0] ;
 wire \RAM[92][1] ;
 wire \RAM[92][2] ;
 wire \RAM[92][3] ;
 wire \RAM[93][0] ;
 wire \RAM[93][1] ;
 wire \RAM[93][2] ;
 wire \RAM[93][3] ;
 wire \RAM[94][0] ;
 wire \RAM[94][1] ;
 wire \RAM[94][2] ;
 wire \RAM[94][3] ;
 wire \RAM[95][0] ;
 wire \RAM[95][1] ;
 wire \RAM[95][2] ;
 wire \RAM[95][3] ;
 wire \RAM[96][0] ;
 wire \RAM[96][1] ;
 wire \RAM[96][2] ;
 wire \RAM[96][3] ;
 wire \RAM[97][0] ;
 wire \RAM[97][1] ;
 wire \RAM[97][2] ;
 wire \RAM[97][3] ;
 wire \RAM[98][0] ;
 wire \RAM[98][1] ;
 wire \RAM[98][2] ;
 wire \RAM[98][3] ;
 wire \RAM[99][0] ;
 wire \RAM[99][1] ;
 wire \RAM[99][2] ;
 wire \RAM[99][3] ;
 wire \RAM[9][0] ;
 wire \RAM[9][1] ;
 wire \RAM[9][2] ;
 wire \RAM[9][3] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net73));
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_30 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_83 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__inv_2 _0991_ (.A(net7),
    .Y(_0512_));
 sky130_fd_sc_hd__clkinv_4 _0992_ (.A(net84),
    .Y(_0513_));
 sky130_fd_sc_hd__inv_2 _0993_ (.A(net75),
    .Y(_0514_));
 sky130_fd_sc_hd__nor2_1 _0994_ (.A(net69),
    .B(net6),
    .Y(_0515_));
 sky130_fd_sc_hd__or2_4 _0995_ (.A(net69),
    .B(net6),
    .X(_0516_));
 sky130_fd_sc_hd__mux2_1 _0996_ (.A0(\RAM[70][0] ),
    .A1(\RAM[71][0] ),
    .S(net142),
    .X(_0517_));
 sky130_fd_sc_hd__mux2_1 _0997_ (.A0(\RAM[68][0] ),
    .A1(\RAM[69][0] ),
    .S(net142),
    .X(_0518_));
 sky130_fd_sc_hd__a21o_1 _0998_ (.A1(net34),
    .A2(_0518_),
    .B1(net31),
    .X(_0519_));
 sky130_fd_sc_hd__a21oi_1 _0999_ (.A1(net90),
    .A2(_0517_),
    .B1(_0519_),
    .Y(_0520_));
 sky130_fd_sc_hd__mux4_1 _1000_ (.A0(\RAM[64][0] ),
    .A1(\RAM[65][0] ),
    .A2(\RAM[66][0] ),
    .A3(\RAM[67][0] ),
    .S0(net143),
    .S1(net90),
    .X(_0521_));
 sky130_fd_sc_hd__nor2_1 _1001_ (.A(net74),
    .B(_0521_),
    .Y(_0522_));
 sky130_fd_sc_hd__mux4_1 _1002_ (.A0(\RAM[72][0] ),
    .A1(\RAM[73][0] ),
    .A2(\RAM[74][0] ),
    .A3(\RAM[75][0] ),
    .S0(net135),
    .S1(net84),
    .X(_0523_));
 sky130_fd_sc_hd__mux2_1 _1003_ (.A0(\RAM[76][0] ),
    .A1(\RAM[77][0] ),
    .S(net142),
    .X(_0524_));
 sky130_fd_sc_hd__mux2_1 _1004_ (.A0(\RAM[78][0] ),
    .A1(\RAM[79][0] ),
    .S(net142),
    .X(_0525_));
 sky130_fd_sc_hd__a21o_1 _1005_ (.A1(net35),
    .A2(_0524_),
    .B1(net31),
    .X(_0526_));
 sky130_fd_sc_hd__a21oi_1 _1006_ (.A1(net91),
    .A2(_0525_),
    .B1(_0526_),
    .Y(_0527_));
 sky130_fd_sc_hd__o21ai_1 _1007_ (.A1(net73),
    .A2(_0523_),
    .B1(net70),
    .Y(_0528_));
 sky130_fd_sc_hd__o32a_1 _1008_ (.A1(net71),
    .A2(_0520_),
    .A3(_0522_),
    .B1(_0527_),
    .B2(_0528_),
    .X(_0529_));
 sky130_fd_sc_hd__nor2_1 _1009_ (.A(_0516_),
    .B(_0529_),
    .Y(_0530_));
 sky130_fd_sc_hd__nand2_8 _1010_ (.A(net69),
    .B(net6),
    .Y(_0531_));
 sky130_fd_sc_hd__and2b_2 _1011_ (.A_N(net71),
    .B(net74),
    .X(_0532_));
 sky130_fd_sc_hd__nand2b_4 _1012_ (.A_N(net72),
    .B(net73),
    .Y(_0533_));
 sky130_fd_sc_hd__nand2_8 _1013_ (.A(net130),
    .B(net79),
    .Y(_0534_));
 sky130_fd_sc_hd__nand2_8 _1014_ (.A(net130),
    .B(net35),
    .Y(_0535_));
 sky130_fd_sc_hd__mux4_1 _1015_ (.A0(\RAM[116][0] ),
    .A1(\RAM[117][0] ),
    .A2(\RAM[118][0] ),
    .A3(\RAM[119][0] ),
    .S0(net143),
    .S1(net90),
    .X(_0536_));
 sky130_fd_sc_hd__o21ba_1 _1016_ (.A1(net28),
    .A2(_0536_),
    .B1_N(_0531_),
    .X(_0537_));
 sky130_fd_sc_hd__nor2_1 _1017_ (.A(net75),
    .B(net72),
    .Y(_0538_));
 sky130_fd_sc_hd__or2_4 _1018_ (.A(net73),
    .B(net72),
    .X(_0539_));
 sky130_fd_sc_hd__mux4_1 _1019_ (.A0(\RAM[112][0] ),
    .A1(\RAM[113][0] ),
    .A2(\RAM[114][0] ),
    .A3(\RAM[115][0] ),
    .S0(net130),
    .S1(net83),
    .X(_0540_));
 sky130_fd_sc_hd__and2_4 _1020_ (.A(net32),
    .B(net72),
    .X(_0541_));
 sky130_fd_sc_hd__nand2b_4 _1021_ (.A_N(net73),
    .B(net70),
    .Y(_0542_));
 sky130_fd_sc_hd__mux4_1 _1022_ (.A0(\RAM[120][0] ),
    .A1(\RAM[121][0] ),
    .A2(\RAM[122][0] ),
    .A3(\RAM[123][0] ),
    .S0(net136),
    .S1(net83),
    .X(_0543_));
 sky130_fd_sc_hd__and2_2 _1023_ (.A(net75),
    .B(net72),
    .X(_0544_));
 sky130_fd_sc_hd__nand2_4 _1024_ (.A(net73),
    .B(net70),
    .Y(_0545_));
 sky130_fd_sc_hd__mux4_2 _1025_ (.A0(\RAM[124][0] ),
    .A1(\RAM[125][0] ),
    .A2(\RAM[126][0] ),
    .A3(\RAM[127][0] ),
    .S0(net129),
    .S1(net81),
    .X(_0546_));
 sky130_fd_sc_hd__o22a_1 _1026_ (.A1(net24),
    .A2(_0543_),
    .B1(net22),
    .B2(_0546_),
    .X(_0547_));
 sky130_fd_sc_hd__o211a_1 _1027_ (.A1(net25),
    .A2(_0540_),
    .B1(_0547_),
    .C1(_0537_),
    .X(_0548_));
 sky130_fd_sc_hd__mux2_1 _1028_ (.A0(\RAM[104][0] ),
    .A1(\RAM[105][0] ),
    .S(net135),
    .X(_0549_));
 sky130_fd_sc_hd__or2_1 _1029_ (.A(net83),
    .B(_0549_),
    .X(_0550_));
 sky130_fd_sc_hd__mux2_1 _1030_ (.A0(\RAM[106][0] ),
    .A1(\RAM[107][0] ),
    .S(net135),
    .X(_0551_));
 sky130_fd_sc_hd__or2_1 _1031_ (.A(net35),
    .B(_0551_),
    .X(_0552_));
 sky130_fd_sc_hd__mux4_1 _1032_ (.A0(\RAM[96][0] ),
    .A1(\RAM[97][0] ),
    .A2(\RAM[98][0] ),
    .A3(\RAM[99][0] ),
    .S0(net133),
    .S1(net81),
    .X(_0553_));
 sky130_fd_sc_hd__a32o_1 _1033_ (.A1(_0541_),
    .A2(_0550_),
    .A3(_0552_),
    .B1(_0553_),
    .B2(net26),
    .X(_0554_));
 sky130_fd_sc_hd__mux4_2 _1034_ (.A0(\RAM[108][0] ),
    .A1(\RAM[109][0] ),
    .A2(\RAM[110][0] ),
    .A3(\RAM[111][0] ),
    .S0(net134),
    .S1(net81),
    .X(_0555_));
 sky130_fd_sc_hd__mux4_1 _1035_ (.A0(\RAM[100][0] ),
    .A1(\RAM[101][0] ),
    .A2(\RAM[102][0] ),
    .A3(\RAM[103][0] ),
    .S0(net133),
    .S1(net82),
    .X(_0556_));
 sky130_fd_sc_hd__a22o_1 _1036_ (.A1(net23),
    .A2(_0555_),
    .B1(_0556_),
    .B2(net29),
    .X(_0557_));
 sky130_fd_sc_hd__and2b_4 _1037_ (.A_N(net69),
    .B(net6),
    .X(_0558_));
 sky130_fd_sc_hd__nand2b_4 _1038_ (.A_N(net69),
    .B(net6),
    .Y(_0559_));
 sky130_fd_sc_hd__o21a_1 _1039_ (.A1(_0554_),
    .A2(_0557_),
    .B1(_0558_),
    .X(_0560_));
 sky130_fd_sc_hd__nand2b_4 _1040_ (.A_N(net6),
    .B(net69),
    .Y(_0561_));
 sky130_fd_sc_hd__mux4_2 _1041_ (.A0(\RAM[84][0] ),
    .A1(\RAM[85][0] ),
    .A2(\RAM[86][0] ),
    .A3(\RAM[87][0] ),
    .S0(net146),
    .S1(net92),
    .X(_0562_));
 sky130_fd_sc_hd__mux4_1 _1042_ (.A0(\RAM[88][0] ),
    .A1(\RAM[89][0] ),
    .A2(\RAM[90][0] ),
    .A3(\RAM[91][0] ),
    .S0(net138),
    .S1(net90),
    .X(_0563_));
 sky130_fd_sc_hd__a22o_1 _1043_ (.A1(net29),
    .A2(_0562_),
    .B1(_0563_),
    .B2(_0541_),
    .X(_0564_));
 sky130_fd_sc_hd__mux4_1 _1044_ (.A0(\RAM[92][0] ),
    .A1(\RAM[93][0] ),
    .A2(\RAM[94][0] ),
    .A3(\RAM[95][0] ),
    .S0(net138),
    .S1(net86),
    .X(_0565_));
 sky130_fd_sc_hd__mux4_2 _1045_ (.A0(\RAM[80][0] ),
    .A1(\RAM[81][0] ),
    .A2(\RAM[82][0] ),
    .A3(\RAM[83][0] ),
    .S0(net138),
    .S1(net86),
    .X(_0566_));
 sky130_fd_sc_hd__a22o_1 _1046_ (.A1(net23),
    .A2(_0565_),
    .B1(_0566_),
    .B2(net26),
    .X(_0567_));
 sky130_fd_sc_hd__o21ba_1 _1047_ (.A1(_0564_),
    .A2(_0567_),
    .B1_N(net21),
    .X(_0568_));
 sky130_fd_sc_hd__or4_1 _1048_ (.A(_0512_),
    .B(_0548_),
    .C(_0560_),
    .D(_0568_),
    .X(_0569_));
 sky130_fd_sc_hd__mux4_1 _1049_ (.A0(\RAM[32][0] ),
    .A1(\RAM[33][0] ),
    .A2(\RAM[34][0] ),
    .A3(\RAM[35][0] ),
    .S0(net131),
    .S1(net79),
    .X(_0570_));
 sky130_fd_sc_hd__mux4_2 _1050_ (.A0(\RAM[44][0] ),
    .A1(\RAM[45][0] ),
    .A2(\RAM[46][0] ),
    .A3(\RAM[47][0] ),
    .S0(net128),
    .S1(net77),
    .X(_0571_));
 sky130_fd_sc_hd__mux4_1 _1051_ (.A0(\RAM[40][0] ),
    .A1(\RAM[41][0] ),
    .A2(\RAM[42][0] ),
    .A3(\RAM[43][0] ),
    .S0(net129),
    .S1(net77),
    .X(_0572_));
 sky130_fd_sc_hd__or2_1 _1052_ (.A(net73),
    .B(_0572_),
    .X(_0573_));
 sky130_fd_sc_hd__o211a_1 _1053_ (.A1(net33),
    .A2(_0571_),
    .B1(_0573_),
    .C1(net70),
    .X(_0574_));
 sky130_fd_sc_hd__mux4_1 _1054_ (.A0(\RAM[36][0] ),
    .A1(\RAM[37][0] ),
    .A2(\RAM[38][0] ),
    .A3(\RAM[39][0] ),
    .S0(net131),
    .S1(net79),
    .X(_0575_));
 sky130_fd_sc_hd__a22o_1 _1055_ (.A1(net26),
    .A2(_0570_),
    .B1(_0575_),
    .B2(net29),
    .X(_0576_));
 sky130_fd_sc_hd__mux4_1 _1056_ (.A0(\RAM[52][0] ),
    .A1(\RAM[53][0] ),
    .A2(\RAM[54][0] ),
    .A3(\RAM[55][0] ),
    .S0(net130),
    .S1(net79),
    .X(_0577_));
 sky130_fd_sc_hd__mux4_1 _1057_ (.A0(\RAM[56][0] ),
    .A1(\RAM[57][0] ),
    .A2(\RAM[58][0] ),
    .A3(\RAM[59][0] ),
    .S0(net130),
    .S1(net80),
    .X(_0578_));
 sky130_fd_sc_hd__o22a_1 _1058_ (.A1(net28),
    .A2(_0577_),
    .B1(_0578_),
    .B2(net24),
    .X(_0579_));
 sky130_fd_sc_hd__mux4_2 _1059_ (.A0(\RAM[60][0] ),
    .A1(\RAM[61][0] ),
    .A2(\RAM[62][0] ),
    .A3(\RAM[63][0] ),
    .S0(net131),
    .S1(net79),
    .X(_0580_));
 sky130_fd_sc_hd__mux4_2 _1060_ (.A0(\RAM[48][0] ),
    .A1(\RAM[49][0] ),
    .A2(\RAM[50][0] ),
    .A3(\RAM[51][0] ),
    .S0(net131),
    .S1(net79),
    .X(_0581_));
 sky130_fd_sc_hd__o22a_1 _1061_ (.A1(net22),
    .A2(_0580_),
    .B1(_0581_),
    .B2(net25),
    .X(_0582_));
 sky130_fd_sc_hd__a21bo_1 _1062_ (.A1(_0579_),
    .A2(_0582_),
    .B1_N(net69),
    .X(_0583_));
 sky130_fd_sc_hd__o311a_2 _1063_ (.A1(net69),
    .A2(_0574_),
    .A3(_0576_),
    .B1(_0583_),
    .C1(net6),
    .X(_0584_));
 sky130_fd_sc_hd__mux2_1 _1064_ (.A0(\RAM[6][0] ),
    .A1(\RAM[7][0] ),
    .S(net144),
    .X(_0585_));
 sky130_fd_sc_hd__and2_1 _1065_ (.A(net92),
    .B(_0585_),
    .X(_0586_));
 sky130_fd_sc_hd__mux2_1 _1066_ (.A0(\RAM[4][0] ),
    .A1(\RAM[5][0] ),
    .S(net144),
    .X(_0587_));
 sky130_fd_sc_hd__a211o_1 _1067_ (.A1(net34),
    .A2(_0587_),
    .B1(_0586_),
    .C1(net31),
    .X(_0588_));
 sky130_fd_sc_hd__mux4_1 _1068_ (.A0(\RAM[0][0] ),
    .A1(\RAM[1][0] ),
    .A2(\RAM[2][0] ),
    .A3(\RAM[3][0] ),
    .S0(net146),
    .S1(net92),
    .X(_0589_));
 sky130_fd_sc_hd__o21ba_1 _1069_ (.A1(net74),
    .A2(_0589_),
    .B1_N(net71),
    .X(_0590_));
 sky130_fd_sc_hd__mux4_1 _1070_ (.A0(\RAM[8][0] ),
    .A1(\RAM[9][0] ),
    .A2(\RAM[10][0] ),
    .A3(\RAM[11][0] ),
    .S0(net143),
    .S1(net90),
    .X(_0591_));
 sky130_fd_sc_hd__or2_1 _1071_ (.A(net74),
    .B(_0591_),
    .X(_0592_));
 sky130_fd_sc_hd__mux2_1 _1072_ (.A0(\RAM[12][0] ),
    .A1(\RAM[13][0] ),
    .S(net144),
    .X(_0593_));
 sky130_fd_sc_hd__mux2_1 _1073_ (.A0(\RAM[14][0] ),
    .A1(\RAM[15][0] ),
    .S(net144),
    .X(_0594_));
 sky130_fd_sc_hd__a21o_1 _1074_ (.A1(net34),
    .A2(_0593_),
    .B1(net31),
    .X(_0595_));
 sky130_fd_sc_hd__a21o_1 _1075_ (.A1(net92),
    .A2(_0594_),
    .B1(_0595_),
    .X(_0596_));
 sky130_fd_sc_hd__a32o_2 _1076_ (.A1(net71),
    .A2(_0592_),
    .A3(_0596_),
    .B1(_0588_),
    .B2(_0590_),
    .X(_0597_));
 sky130_fd_sc_hd__mux4_1 _1077_ (.A0(\RAM[20][0] ),
    .A1(\RAM[21][0] ),
    .A2(\RAM[22][0] ),
    .A3(\RAM[23][0] ),
    .S0(net141),
    .S1(net87),
    .X(_0598_));
 sky130_fd_sc_hd__mux4_1 _1078_ (.A0(\RAM[24][0] ),
    .A1(\RAM[25][0] ),
    .A2(\RAM[26][0] ),
    .A3(\RAM[27][0] ),
    .S0(net140),
    .S1(net87),
    .X(_0599_));
 sky130_fd_sc_hd__a22o_1 _1079_ (.A1(net29),
    .A2(_0598_),
    .B1(_0599_),
    .B2(_0541_),
    .X(_0600_));
 sky130_fd_sc_hd__mux4_1 _1080_ (.A0(\RAM[28][0] ),
    .A1(\RAM[29][0] ),
    .A2(\RAM[30][0] ),
    .A3(\RAM[31][0] ),
    .S0(net140),
    .S1(net87),
    .X(_0601_));
 sky130_fd_sc_hd__mux4_1 _1081_ (.A0(\RAM[16][0] ),
    .A1(\RAM[17][0] ),
    .A2(\RAM[18][0] ),
    .A3(\RAM[19][0] ),
    .S0(net140),
    .S1(net87),
    .X(_0602_));
 sky130_fd_sc_hd__a22o_1 _1082_ (.A1(net23),
    .A2(_0601_),
    .B1(_0602_),
    .B2(net26),
    .X(_0603_));
 sky130_fd_sc_hd__o21ba_1 _1083_ (.A1(_0600_),
    .A2(_0603_),
    .B1_N(net21),
    .X(_0604_));
 sky130_fd_sc_hd__a211o_1 _1084_ (.A1(_0515_),
    .A2(_0597_),
    .B1(_0604_),
    .C1(_0584_),
    .X(_0605_));
 sky130_fd_sc_hd__o22a_2 _1085_ (.A1(_0530_),
    .A2(_0569_),
    .B1(_0605_),
    .B2(net7),
    .X(net13));
 sky130_fd_sc_hd__mux4_1 _1086_ (.A0(\RAM[44][1] ),
    .A1(\RAM[45][1] ),
    .A2(\RAM[46][1] ),
    .A3(\RAM[47][1] ),
    .S0(net128),
    .S1(net77),
    .X(_0606_));
 sky130_fd_sc_hd__mux4_2 _1087_ (.A0(\RAM[36][1] ),
    .A1(\RAM[37][1] ),
    .A2(\RAM[38][1] ),
    .A3(\RAM[39][1] ),
    .S0(net128),
    .S1(net77),
    .X(_0607_));
 sky130_fd_sc_hd__mux4_1 _1088_ (.A0(\RAM[32][1] ),
    .A1(\RAM[33][1] ),
    .A2(\RAM[34][1] ),
    .A3(\RAM[35][1] ),
    .S0(net128),
    .S1(net77),
    .X(_0608_));
 sky130_fd_sc_hd__mux4_1 _1089_ (.A0(\RAM[40][1] ),
    .A1(\RAM[41][1] ),
    .A2(\RAM[42][1] ),
    .A3(\RAM[43][1] ),
    .S0(net129),
    .S1(net78),
    .X(_0609_));
 sky130_fd_sc_hd__mux4_2 _1090_ (.A0(_0607_),
    .A1(_0608_),
    .A2(_0606_),
    .A3(_0609_),
    .S0(net33),
    .S1(net70),
    .X(_0610_));
 sky130_fd_sc_hd__mux4_1 _1091_ (.A0(\RAM[52][1] ),
    .A1(\RAM[53][1] ),
    .A2(\RAM[54][1] ),
    .A3(\RAM[55][1] ),
    .S0(net139),
    .S1(net86),
    .X(_0611_));
 sky130_fd_sc_hd__mux4_1 _1092_ (.A0(\RAM[56][1] ),
    .A1(\RAM[57][1] ),
    .A2(\RAM[58][1] ),
    .A3(\RAM[59][1] ),
    .S0(net130),
    .S1(net80),
    .X(_0612_));
 sky130_fd_sc_hd__o22a_2 _1093_ (.A1(net28),
    .A2(_0611_),
    .B1(_0612_),
    .B2(net24),
    .X(_0613_));
 sky130_fd_sc_hd__mux4_2 _1094_ (.A0(\RAM[60][1] ),
    .A1(\RAM[61][1] ),
    .A2(\RAM[62][1] ),
    .A3(\RAM[63][1] ),
    .S0(net131),
    .S1(net79),
    .X(_0614_));
 sky130_fd_sc_hd__mux4_2 _1095_ (.A0(\RAM[48][1] ),
    .A1(\RAM[49][1] ),
    .A2(\RAM[50][1] ),
    .A3(\RAM[51][1] ),
    .S0(net131),
    .S1(net79),
    .X(_0615_));
 sky130_fd_sc_hd__o221ai_4 _1096_ (.A1(net22),
    .A2(_0614_),
    .B1(_0615_),
    .B2(net25),
    .C1(_0613_),
    .Y(_0616_));
 sky130_fd_sc_hd__o21ai_1 _1097_ (.A1(net5),
    .A2(_0610_),
    .B1(net6),
    .Y(_0617_));
 sky130_fd_sc_hd__a21o_1 _1098_ (.A1(net5),
    .A2(_0616_),
    .B1(_0617_),
    .X(_0618_));
 sky130_fd_sc_hd__mux2_1 _1099_ (.A0(\RAM[6][1] ),
    .A1(\RAM[7][1] ),
    .S(net144),
    .X(_0619_));
 sky130_fd_sc_hd__nand2_1 _1100_ (.A(net93),
    .B(_0619_),
    .Y(_0620_));
 sky130_fd_sc_hd__mux2_1 _1101_ (.A0(\RAM[4][1] ),
    .A1(\RAM[5][1] ),
    .S(net145),
    .X(_0621_));
 sky130_fd_sc_hd__a21oi_1 _1102_ (.A1(net34),
    .A2(_0621_),
    .B1(net31),
    .Y(_0622_));
 sky130_fd_sc_hd__mux4_1 _1103_ (.A0(\RAM[0][1] ),
    .A1(\RAM[1][1] ),
    .A2(\RAM[2][1] ),
    .A3(\RAM[3][1] ),
    .S0(net146),
    .S1(net93),
    .X(_0623_));
 sky130_fd_sc_hd__a2bb2o_1 _1104_ (.A1_N(net74),
    .A2_N(_0623_),
    .B1(_0620_),
    .B2(_0622_),
    .X(_0624_));
 sky130_fd_sc_hd__mux4_1 _1105_ (.A0(\RAM[8][1] ),
    .A1(\RAM[9][1] ),
    .A2(\RAM[10][1] ),
    .A3(\RAM[11][1] ),
    .S0(net143),
    .S1(net90),
    .X(_0625_));
 sky130_fd_sc_hd__mux2_1 _1106_ (.A0(\RAM[12][1] ),
    .A1(\RAM[13][1] ),
    .S(net144),
    .X(_0626_));
 sky130_fd_sc_hd__mux2_1 _1107_ (.A0(\RAM[14][1] ),
    .A1(\RAM[15][1] ),
    .S(net147),
    .X(_0627_));
 sky130_fd_sc_hd__a21o_1 _1108_ (.A1(net34),
    .A2(_0626_),
    .B1(net31),
    .X(_0628_));
 sky130_fd_sc_hd__a21oi_1 _1109_ (.A1(net91),
    .A2(_0627_),
    .B1(_0628_),
    .Y(_0629_));
 sky130_fd_sc_hd__o21ai_1 _1110_ (.A1(net74),
    .A2(_0625_),
    .B1(net71),
    .Y(_0630_));
 sky130_fd_sc_hd__o22a_1 _1111_ (.A1(net71),
    .A2(_0624_),
    .B1(_0629_),
    .B2(_0630_),
    .X(_0631_));
 sky130_fd_sc_hd__mux4_2 _1112_ (.A0(\RAM[20][1] ),
    .A1(\RAM[21][1] ),
    .A2(\RAM[22][1] ),
    .A3(\RAM[23][1] ),
    .S0(net141),
    .S1(net88),
    .X(_0632_));
 sky130_fd_sc_hd__mux4_1 _1113_ (.A0(\RAM[24][1] ),
    .A1(\RAM[25][1] ),
    .A2(\RAM[26][1] ),
    .A3(\RAM[27][1] ),
    .S0(net141),
    .S1(net88),
    .X(_0633_));
 sky130_fd_sc_hd__a22o_1 _1114_ (.A1(net29),
    .A2(_0632_),
    .B1(_0633_),
    .B2(_0541_),
    .X(_0634_));
 sky130_fd_sc_hd__mux4_1 _1115_ (.A0(\RAM[28][1] ),
    .A1(\RAM[29][1] ),
    .A2(\RAM[30][1] ),
    .A3(\RAM[31][1] ),
    .S0(net140),
    .S1(net87),
    .X(_0635_));
 sky130_fd_sc_hd__mux4_2 _1116_ (.A0(\RAM[16][1] ),
    .A1(\RAM[17][1] ),
    .A2(\RAM[18][1] ),
    .A3(\RAM[19][1] ),
    .S0(net140),
    .S1(net87),
    .X(_0636_));
 sky130_fd_sc_hd__a22o_1 _1117_ (.A1(net23),
    .A2(_0635_),
    .B1(_0636_),
    .B2(net26),
    .X(_0637_));
 sky130_fd_sc_hd__nor2_1 _1118_ (.A(_0634_),
    .B(_0637_),
    .Y(_0638_));
 sky130_fd_sc_hd__o221a_2 _1119_ (.A1(_0516_),
    .A2(_0631_),
    .B1(_0638_),
    .B2(net21),
    .C1(_0512_),
    .X(_0639_));
 sky130_fd_sc_hd__mux2_1 _1120_ (.A0(\RAM[70][1] ),
    .A1(\RAM[71][1] ),
    .S(net142),
    .X(_0640_));
 sky130_fd_sc_hd__mux2_1 _1121_ (.A0(\RAM[68][1] ),
    .A1(\RAM[69][1] ),
    .S(net147),
    .X(_0641_));
 sky130_fd_sc_hd__a21o_1 _1122_ (.A1(net34),
    .A2(_0641_),
    .B1(net31),
    .X(_0642_));
 sky130_fd_sc_hd__a21oi_1 _1123_ (.A1(net91),
    .A2(_0640_),
    .B1(_0642_),
    .Y(_0643_));
 sky130_fd_sc_hd__mux4_1 _1124_ (.A0(\RAM[64][1] ),
    .A1(\RAM[65][1] ),
    .A2(\RAM[66][1] ),
    .A3(\RAM[67][1] ),
    .S0(net143),
    .S1(net91),
    .X(_0644_));
 sky130_fd_sc_hd__nor2_1 _1125_ (.A(net74),
    .B(_0644_),
    .Y(_0645_));
 sky130_fd_sc_hd__mux4_1 _1126_ (.A0(\RAM[72][1] ),
    .A1(\RAM[73][1] ),
    .A2(\RAM[74][1] ),
    .A3(\RAM[75][1] ),
    .S0(net135),
    .S1(net84),
    .X(_0646_));
 sky130_fd_sc_hd__mux2_1 _1127_ (.A0(\RAM[76][1] ),
    .A1(\RAM[77][1] ),
    .S(net135),
    .X(_0647_));
 sky130_fd_sc_hd__mux2_1 _1128_ (.A0(\RAM[78][1] ),
    .A1(\RAM[79][1] ),
    .S(net135),
    .X(_0648_));
 sky130_fd_sc_hd__a21o_1 _1129_ (.A1(net35),
    .A2(_0647_),
    .B1(net33),
    .X(_0649_));
 sky130_fd_sc_hd__a21oi_1 _1130_ (.A1(net84),
    .A2(_0648_),
    .B1(_0649_),
    .Y(_0650_));
 sky130_fd_sc_hd__o21ai_1 _1131_ (.A1(net73),
    .A2(_0646_),
    .B1(net70),
    .Y(_0651_));
 sky130_fd_sc_hd__o32a_1 _1132_ (.A1(net71),
    .A2(_0643_),
    .A3(_0645_),
    .B1(_0650_),
    .B2(_0651_),
    .X(_0652_));
 sky130_fd_sc_hd__mux4_1 _1133_ (.A0(\RAM[116][1] ),
    .A1(\RAM[117][1] ),
    .A2(\RAM[118][1] ),
    .A3(\RAM[119][1] ),
    .S0(net136),
    .S1(net83),
    .X(_0653_));
 sky130_fd_sc_hd__o21ba_1 _1134_ (.A1(net28),
    .A2(_0653_),
    .B1_N(_0531_),
    .X(_0654_));
 sky130_fd_sc_hd__mux4_1 _1135_ (.A0(\RAM[112][1] ),
    .A1(\RAM[113][1] ),
    .A2(\RAM[114][1] ),
    .A3(\RAM[115][1] ),
    .S0(net129),
    .S1(net81),
    .X(_0655_));
 sky130_fd_sc_hd__mux4_1 _1136_ (.A0(\RAM[120][1] ),
    .A1(\RAM[121][1] ),
    .A2(\RAM[122][1] ),
    .A3(\RAM[123][1] ),
    .S0(net136),
    .S1(net83),
    .X(_0656_));
 sky130_fd_sc_hd__mux4_2 _1137_ (.A0(\RAM[124][1] ),
    .A1(\RAM[125][1] ),
    .A2(\RAM[126][1] ),
    .A3(\RAM[127][1] ),
    .S0(net133),
    .S1(net81),
    .X(_0657_));
 sky130_fd_sc_hd__o22a_1 _1138_ (.A1(net24),
    .A2(_0656_),
    .B1(_0657_),
    .B2(net22),
    .X(_0658_));
 sky130_fd_sc_hd__o211a_1 _1139_ (.A1(net25),
    .A2(_0655_),
    .B1(_0658_),
    .C1(_0654_),
    .X(_0659_));
 sky130_fd_sc_hd__mux4_1 _1140_ (.A0(\RAM[100][1] ),
    .A1(\RAM[101][1] ),
    .A2(\RAM[102][1] ),
    .A3(\RAM[103][1] ),
    .S0(net133),
    .S1(net82),
    .X(_0660_));
 sky130_fd_sc_hd__mux4_1 _1141_ (.A0(\RAM[108][1] ),
    .A1(\RAM[109][1] ),
    .A2(\RAM[110][1] ),
    .A3(\RAM[111][1] ),
    .S0(net134),
    .S1(net82),
    .X(_0661_));
 sky130_fd_sc_hd__mux4_2 _1142_ (.A0(\RAM[96][1] ),
    .A1(\RAM[97][1] ),
    .A2(\RAM[98][1] ),
    .A3(\RAM[99][1] ),
    .S0(net133),
    .S1(net81),
    .X(_0662_));
 sky130_fd_sc_hd__a22o_1 _1143_ (.A1(net29),
    .A2(_0660_),
    .B1(_0662_),
    .B2(net26),
    .X(_0663_));
 sky130_fd_sc_hd__mux4_1 _1144_ (.A0(\RAM[104][1] ),
    .A1(\RAM[105][1] ),
    .A2(\RAM[106][1] ),
    .A3(\RAM[107][1] ),
    .S0(net134),
    .S1(net82),
    .X(_0664_));
 sky130_fd_sc_hd__or2_1 _1145_ (.A(net73),
    .B(_0664_),
    .X(_0665_));
 sky130_fd_sc_hd__or2_1 _1146_ (.A(net33),
    .B(_0661_),
    .X(_0666_));
 sky130_fd_sc_hd__a31o_1 _1147_ (.A1(net70),
    .A2(_0665_),
    .A3(_0666_),
    .B1(_0663_),
    .X(_0667_));
 sky130_fd_sc_hd__a21oi_2 _1148_ (.A1(_0558_),
    .A2(_0667_),
    .B1(_0659_),
    .Y(_0668_));
 sky130_fd_sc_hd__mux4_2 _1149_ (.A0(\RAM[84][1] ),
    .A1(\RAM[85][1] ),
    .A2(\RAM[86][1] ),
    .A3(\RAM[87][1] ),
    .S0(net146),
    .S1(net92),
    .X(_0669_));
 sky130_fd_sc_hd__mux4_1 _1150_ (.A0(\RAM[88][1] ),
    .A1(\RAM[89][1] ),
    .A2(\RAM[90][1] ),
    .A3(\RAM[91][1] ),
    .S0(net143),
    .S1(net90),
    .X(_0670_));
 sky130_fd_sc_hd__a22o_1 _1151_ (.A1(net30),
    .A2(_0669_),
    .B1(_0670_),
    .B2(_0541_),
    .X(_0671_));
 sky130_fd_sc_hd__mux4_1 _1152_ (.A0(\RAM[92][1] ),
    .A1(\RAM[93][1] ),
    .A2(\RAM[94][1] ),
    .A3(\RAM[95][1] ),
    .S0(net138),
    .S1(net86),
    .X(_0672_));
 sky130_fd_sc_hd__mux4_2 _1153_ (.A0(\RAM[80][1] ),
    .A1(\RAM[81][1] ),
    .A2(\RAM[82][1] ),
    .A3(\RAM[83][1] ),
    .S0(net138),
    .S1(net86),
    .X(_0673_));
 sky130_fd_sc_hd__a22o_1 _1154_ (.A1(net23),
    .A2(_0672_),
    .B1(_0673_),
    .B2(net27),
    .X(_0674_));
 sky130_fd_sc_hd__nor2_1 _1155_ (.A(_0671_),
    .B(_0674_),
    .Y(_0675_));
 sky130_fd_sc_hd__o221a_2 _1156_ (.A1(_0516_),
    .A2(_0652_),
    .B1(_0675_),
    .B2(net21),
    .C1(_0668_),
    .X(_0676_));
 sky130_fd_sc_hd__a22oi_4 _1157_ (.A1(_0618_),
    .A2(_0639_),
    .B1(_0676_),
    .B2(net7),
    .Y(net14));
 sky130_fd_sc_hd__mux4_1 _1158_ (.A0(\RAM[96][2] ),
    .A1(\RAM[97][2] ),
    .A2(\RAM[98][2] ),
    .A3(\RAM[99][2] ),
    .S0(net133),
    .S1(net81),
    .X(_0677_));
 sky130_fd_sc_hd__mux4_2 _1159_ (.A0(\RAM[108][2] ),
    .A1(\RAM[109][2] ),
    .A2(\RAM[110][2] ),
    .A3(\RAM[111][2] ),
    .S0(net134),
    .S1(net82),
    .X(_0678_));
 sky130_fd_sc_hd__mux4_1 _1160_ (.A0(\RAM[104][2] ),
    .A1(\RAM[105][2] ),
    .A2(\RAM[106][2] ),
    .A3(\RAM[107][2] ),
    .S0(net135),
    .S1(net84),
    .X(_0679_));
 sky130_fd_sc_hd__or2_1 _1161_ (.A(net73),
    .B(_0679_),
    .X(_0680_));
 sky130_fd_sc_hd__o211a_1 _1162_ (.A1(net33),
    .A2(_0678_),
    .B1(_0680_),
    .C1(net70),
    .X(_0681_));
 sky130_fd_sc_hd__mux4_1 _1163_ (.A0(\RAM[100][2] ),
    .A1(\RAM[101][2] ),
    .A2(\RAM[102][2] ),
    .A3(\RAM[103][2] ),
    .S0(net133),
    .S1(net81),
    .X(_0682_));
 sky130_fd_sc_hd__a22o_1 _1164_ (.A1(net26),
    .A2(_0677_),
    .B1(_0682_),
    .B2(net29),
    .X(_0683_));
 sky130_fd_sc_hd__mux4_1 _1165_ (.A0(\RAM[116][2] ),
    .A1(\RAM[117][2] ),
    .A2(\RAM[118][2] ),
    .A3(\RAM[119][2] ),
    .S0(net136),
    .S1(net83),
    .X(_0684_));
 sky130_fd_sc_hd__mux4_2 _1166_ (.A0(\RAM[120][2] ),
    .A1(\RAM[121][2] ),
    .A2(\RAM[122][2] ),
    .A3(\RAM[123][2] ),
    .S0(net136),
    .S1(net83),
    .X(_0685_));
 sky130_fd_sc_hd__o22a_1 _1167_ (.A1(net28),
    .A2(_0684_),
    .B1(_0685_),
    .B2(net24),
    .X(_0686_));
 sky130_fd_sc_hd__mux4_2 _1168_ (.A0(\RAM[124][2] ),
    .A1(\RAM[125][2] ),
    .A2(\RAM[126][2] ),
    .A3(\RAM[127][2] ),
    .S0(net129),
    .S1(net78),
    .X(_0687_));
 sky130_fd_sc_hd__mux4_1 _1169_ (.A0(\RAM[112][2] ),
    .A1(\RAM[113][2] ),
    .A2(\RAM[114][2] ),
    .A3(\RAM[115][2] ),
    .S0(net129),
    .S1(net78),
    .X(_0688_));
 sky130_fd_sc_hd__o22a_1 _1170_ (.A1(net22),
    .A2(_0687_),
    .B1(_0688_),
    .B2(net25),
    .X(_0689_));
 sky130_fd_sc_hd__a21bo_1 _1171_ (.A1(_0686_),
    .A2(_0689_),
    .B1_N(net69),
    .X(_0690_));
 sky130_fd_sc_hd__o311a_1 _1172_ (.A1(net69),
    .A2(_0681_),
    .A3(_0683_),
    .B1(_0690_),
    .C1(net6),
    .X(_0691_));
 sky130_fd_sc_hd__mux2_1 _1173_ (.A0(\RAM[70][2] ),
    .A1(\RAM[71][2] ),
    .S(net142),
    .X(_0692_));
 sky130_fd_sc_hd__and2_1 _1174_ (.A(net91),
    .B(_0692_),
    .X(_0693_));
 sky130_fd_sc_hd__mux2_1 _1175_ (.A0(\RAM[68][2] ),
    .A1(\RAM[69][2] ),
    .S(net142),
    .X(_0694_));
 sky130_fd_sc_hd__a211o_1 _1176_ (.A1(net34),
    .A2(_0694_),
    .B1(_0693_),
    .C1(net31),
    .X(_0695_));
 sky130_fd_sc_hd__mux4_1 _1177_ (.A0(\RAM[64][2] ),
    .A1(\RAM[65][2] ),
    .A2(\RAM[66][2] ),
    .A3(\RAM[67][2] ),
    .S0(net136),
    .S1(net83),
    .X(_0696_));
 sky130_fd_sc_hd__o21ba_1 _1178_ (.A1(net76),
    .A2(_0696_),
    .B1_N(net71),
    .X(_0697_));
 sky130_fd_sc_hd__mux4_1 _1179_ (.A0(\RAM[72][2] ),
    .A1(\RAM[73][2] ),
    .A2(\RAM[74][2] ),
    .A3(\RAM[75][2] ),
    .S0(net135),
    .S1(net84),
    .X(_0698_));
 sky130_fd_sc_hd__or2_1 _1180_ (.A(net76),
    .B(_0698_),
    .X(_0699_));
 sky130_fd_sc_hd__mux2_1 _1181_ (.A0(\RAM[76][2] ),
    .A1(\RAM[77][2] ),
    .S(net135),
    .X(_0700_));
 sky130_fd_sc_hd__mux2_1 _1182_ (.A0(\RAM[78][2] ),
    .A1(\RAM[79][2] ),
    .S(net137),
    .X(_0701_));
 sky130_fd_sc_hd__a21o_1 _1183_ (.A1(net35),
    .A2(_0700_),
    .B1(net33),
    .X(_0702_));
 sky130_fd_sc_hd__a21o_1 _1184_ (.A1(net84),
    .A2(_0701_),
    .B1(_0702_),
    .X(_0703_));
 sky130_fd_sc_hd__a32o_2 _1185_ (.A1(net71),
    .A2(_0699_),
    .A3(_0703_),
    .B1(_0695_),
    .B2(_0697_),
    .X(_0704_));
 sky130_fd_sc_hd__mux4_2 _1186_ (.A0(\RAM[84][2] ),
    .A1(\RAM[85][2] ),
    .A2(\RAM[86][2] ),
    .A3(\RAM[87][2] ),
    .S0(net146),
    .S1(net92),
    .X(_0705_));
 sky130_fd_sc_hd__mux4_1 _1187_ (.A0(\RAM[88][2] ),
    .A1(\RAM[89][2] ),
    .A2(\RAM[90][2] ),
    .A3(\RAM[91][2] ),
    .S0(net143),
    .S1(net90),
    .X(_0706_));
 sky130_fd_sc_hd__a22o_1 _1188_ (.A1(net30),
    .A2(_0705_),
    .B1(_0706_),
    .B2(_0541_),
    .X(_0707_));
 sky130_fd_sc_hd__mux4_1 _1189_ (.A0(\RAM[92][2] ),
    .A1(\RAM[93][2] ),
    .A2(\RAM[94][2] ),
    .A3(\RAM[95][2] ),
    .S0(net138),
    .S1(net86),
    .X(_0708_));
 sky130_fd_sc_hd__mux4_2 _1190_ (.A0(\RAM[80][2] ),
    .A1(\RAM[81][2] ),
    .A2(\RAM[82][2] ),
    .A3(\RAM[83][2] ),
    .S0(net138),
    .S1(net86),
    .X(_0709_));
 sky130_fd_sc_hd__a22o_1 _1191_ (.A1(net23),
    .A2(_0708_),
    .B1(_0709_),
    .B2(net27),
    .X(_0710_));
 sky130_fd_sc_hd__o21ba_1 _1192_ (.A1(_0707_),
    .A2(_0710_),
    .B1_N(net21),
    .X(_0711_));
 sky130_fd_sc_hd__a211o_1 _1193_ (.A1(_0515_),
    .A2(_0704_),
    .B1(_0711_),
    .C1(_0691_),
    .X(_0712_));
 sky130_fd_sc_hd__mux2_1 _1194_ (.A0(\RAM[6][2] ),
    .A1(\RAM[7][2] ),
    .S(net145),
    .X(_0713_));
 sky130_fd_sc_hd__mux2_1 _1195_ (.A0(\RAM[4][2] ),
    .A1(\RAM[5][2] ),
    .S(net145),
    .X(_0714_));
 sky130_fd_sc_hd__a21o_1 _1196_ (.A1(net34),
    .A2(_0714_),
    .B1(net32),
    .X(_0715_));
 sky130_fd_sc_hd__a21oi_1 _1197_ (.A1(net93),
    .A2(_0713_),
    .B1(_0715_),
    .Y(_0716_));
 sky130_fd_sc_hd__mux4_1 _1198_ (.A0(\RAM[0][2] ),
    .A1(\RAM[1][2] ),
    .A2(\RAM[2][2] ),
    .A3(\RAM[3][2] ),
    .S0(net145),
    .S1(net93),
    .X(_0717_));
 sky130_fd_sc_hd__nor2_1 _1199_ (.A(net74),
    .B(_0717_),
    .Y(_0718_));
 sky130_fd_sc_hd__mux4_1 _1200_ (.A0(\RAM[8][2] ),
    .A1(\RAM[9][2] ),
    .A2(\RAM[10][2] ),
    .A3(\RAM[11][2] ),
    .S0(net146),
    .S1(net93),
    .X(_0719_));
 sky130_fd_sc_hd__mux2_1 _1201_ (.A0(\RAM[12][2] ),
    .A1(\RAM[13][2] ),
    .S(net144),
    .X(_0720_));
 sky130_fd_sc_hd__mux2_1 _1202_ (.A0(\RAM[14][2] ),
    .A1(\RAM[15][2] ),
    .S(net144),
    .X(_0721_));
 sky130_fd_sc_hd__a21o_1 _1203_ (.A1(net34),
    .A2(_0720_),
    .B1(net32),
    .X(_0722_));
 sky130_fd_sc_hd__a21oi_1 _1204_ (.A1(net93),
    .A2(_0721_),
    .B1(_0722_),
    .Y(_0723_));
 sky130_fd_sc_hd__o21ai_1 _1205_ (.A1(net74),
    .A2(_0719_),
    .B1(net72),
    .Y(_0724_));
 sky130_fd_sc_hd__o32a_2 _1206_ (.A1(net72),
    .A2(_0716_),
    .A3(_0718_),
    .B1(_0723_),
    .B2(_0724_),
    .X(_0725_));
 sky130_fd_sc_hd__nor2_1 _1207_ (.A(_0516_),
    .B(_0725_),
    .Y(_0726_));
 sky130_fd_sc_hd__mux4_1 _1208_ (.A0(\RAM[52][2] ),
    .A1(\RAM[53][2] ),
    .A2(\RAM[54][2] ),
    .A3(\RAM[55][2] ),
    .S0(net139),
    .S1(net89),
    .X(_0727_));
 sky130_fd_sc_hd__o21ba_1 _1209_ (.A1(net28),
    .A2(_0727_),
    .B1_N(_0531_),
    .X(_0728_));
 sky130_fd_sc_hd__mux4_2 _1210_ (.A0(\RAM[48][2] ),
    .A1(\RAM[49][2] ),
    .A2(\RAM[50][2] ),
    .A3(\RAM[51][2] ),
    .S0(net138),
    .S1(net86),
    .X(_0729_));
 sky130_fd_sc_hd__mux4_1 _1211_ (.A0(\RAM[56][2] ),
    .A1(\RAM[57][2] ),
    .A2(\RAM[58][2] ),
    .A3(\RAM[59][2] ),
    .S0(net131),
    .S1(net80),
    .X(_0730_));
 sky130_fd_sc_hd__mux4_1 _1212_ (.A0(\RAM[60][2] ),
    .A1(\RAM[61][2] ),
    .A2(\RAM[62][2] ),
    .A3(\RAM[63][2] ),
    .S0(net131),
    .S1(net79),
    .X(_0731_));
 sky130_fd_sc_hd__o22a_1 _1213_ (.A1(net24),
    .A2(_0730_),
    .B1(_0731_),
    .B2(net22),
    .X(_0732_));
 sky130_fd_sc_hd__o211a_1 _1214_ (.A1(net25),
    .A2(_0729_),
    .B1(_0732_),
    .C1(_0728_),
    .X(_0733_));
 sky130_fd_sc_hd__mux4_1 _1215_ (.A0(\RAM[36][2] ),
    .A1(\RAM[37][2] ),
    .A2(\RAM[38][2] ),
    .A3(\RAM[39][2] ),
    .S0(net128),
    .S1(net77),
    .X(_0734_));
 sky130_fd_sc_hd__mux4_1 _1216_ (.A0(\RAM[32][2] ),
    .A1(\RAM[33][2] ),
    .A2(\RAM[34][2] ),
    .A3(\RAM[35][2] ),
    .S0(net128),
    .S1(net77),
    .X(_0735_));
 sky130_fd_sc_hd__a22o_1 _1217_ (.A1(net29),
    .A2(_0734_),
    .B1(_0735_),
    .B2(net26),
    .X(_0736_));
 sky130_fd_sc_hd__mux4_1 _1218_ (.A0(\RAM[44][2] ),
    .A1(\RAM[45][2] ),
    .A2(\RAM[46][2] ),
    .A3(\RAM[47][2] ),
    .S0(net128),
    .S1(net77),
    .X(_0737_));
 sky130_fd_sc_hd__mux4_1 _1219_ (.A0(\RAM[40][2] ),
    .A1(\RAM[41][2] ),
    .A2(\RAM[42][2] ),
    .A3(\RAM[43][2] ),
    .S0(net129),
    .S1(net78),
    .X(_0738_));
 sky130_fd_sc_hd__or2_1 _1220_ (.A(net73),
    .B(_0738_),
    .X(_0739_));
 sky130_fd_sc_hd__o211a_1 _1221_ (.A1(net33),
    .A2(_0737_),
    .B1(_0739_),
    .C1(net70),
    .X(_0740_));
 sky130_fd_sc_hd__o21a_1 _1222_ (.A1(_0736_),
    .A2(_0740_),
    .B1(_0558_),
    .X(_0741_));
 sky130_fd_sc_hd__mux4_1 _1223_ (.A0(\RAM[20][2] ),
    .A1(\RAM[21][2] ),
    .A2(\RAM[22][2] ),
    .A3(\RAM[23][2] ),
    .S0(net141),
    .S1(net88),
    .X(_0742_));
 sky130_fd_sc_hd__mux4_1 _1224_ (.A0(\RAM[24][2] ),
    .A1(\RAM[25][2] ),
    .A2(\RAM[26][2] ),
    .A3(\RAM[27][2] ),
    .S0(net140),
    .S1(net88),
    .X(_0743_));
 sky130_fd_sc_hd__a22o_1 _1225_ (.A1(net30),
    .A2(_0742_),
    .B1(_0743_),
    .B2(_0541_),
    .X(_0744_));
 sky130_fd_sc_hd__mux4_1 _1226_ (.A0(\RAM[28][2] ),
    .A1(\RAM[29][2] ),
    .A2(\RAM[30][2] ),
    .A3(\RAM[31][2] ),
    .S0(net140),
    .S1(net87),
    .X(_0745_));
 sky130_fd_sc_hd__mux4_1 _1227_ (.A0(\RAM[16][2] ),
    .A1(\RAM[17][2] ),
    .A2(\RAM[18][2] ),
    .A3(\RAM[19][2] ),
    .S0(net140),
    .S1(net87),
    .X(_0746_));
 sky130_fd_sc_hd__a22o_1 _1228_ (.A1(net23),
    .A2(_0745_),
    .B1(_0746_),
    .B2(net27),
    .X(_0747_));
 sky130_fd_sc_hd__o21ba_1 _1229_ (.A1(_0744_),
    .A2(_0747_),
    .B1_N(net21),
    .X(_0748_));
 sky130_fd_sc_hd__or4_1 _1230_ (.A(net7),
    .B(_0733_),
    .C(_0741_),
    .D(_0748_),
    .X(_0749_));
 sky130_fd_sc_hd__o22a_2 _1231_ (.A1(_0512_),
    .A2(_0712_),
    .B1(_0726_),
    .B2(_0749_),
    .X(net15));
 sky130_fd_sc_hd__mux2_1 _1232_ (.A0(\RAM[70][3] ),
    .A1(\RAM[71][3] ),
    .S(net142),
    .X(_0750_));
 sky130_fd_sc_hd__mux2_1 _1233_ (.A0(\RAM[68][3] ),
    .A1(\RAM[69][3] ),
    .S(net147),
    .X(_0751_));
 sky130_fd_sc_hd__a21o_1 _1234_ (.A1(net34),
    .A2(_0751_),
    .B1(net31),
    .X(_0752_));
 sky130_fd_sc_hd__a21oi_1 _1235_ (.A1(net91),
    .A2(_0750_),
    .B1(_0752_),
    .Y(_0753_));
 sky130_fd_sc_hd__mux4_1 _1236_ (.A0(\RAM[64][3] ),
    .A1(\RAM[65][3] ),
    .A2(\RAM[66][3] ),
    .A3(\RAM[67][3] ),
    .S0(net143),
    .S1(net91),
    .X(_0754_));
 sky130_fd_sc_hd__nor2_1 _1237_ (.A(net74),
    .B(_0754_),
    .Y(_0755_));
 sky130_fd_sc_hd__mux4_1 _1238_ (.A0(\RAM[72][3] ),
    .A1(\RAM[73][3] ),
    .A2(\RAM[74][3] ),
    .A3(\RAM[75][3] ),
    .S0(net135),
    .S1(net84),
    .X(_0756_));
 sky130_fd_sc_hd__mux2_1 _1239_ (.A0(\RAM[76][3] ),
    .A1(\RAM[77][3] ),
    .S(net142),
    .X(_0757_));
 sky130_fd_sc_hd__mux2_1 _1240_ (.A0(\RAM[78][3] ),
    .A1(\RAM[79][3] ),
    .S(net142),
    .X(_0758_));
 sky130_fd_sc_hd__a21o_1 _1241_ (.A1(net35),
    .A2(_0757_),
    .B1(net31),
    .X(_0759_));
 sky130_fd_sc_hd__a21oi_1 _1242_ (.A1(net91),
    .A2(_0758_),
    .B1(_0759_),
    .Y(_0760_));
 sky130_fd_sc_hd__o21ai_1 _1243_ (.A1(net76),
    .A2(_0756_),
    .B1(net70),
    .Y(_0761_));
 sky130_fd_sc_hd__o32a_1 _1244_ (.A1(net71),
    .A2(_0753_),
    .A3(_0755_),
    .B1(_0760_),
    .B2(_0761_),
    .X(_0762_));
 sky130_fd_sc_hd__mux4_1 _1245_ (.A0(\RAM[116][3] ),
    .A1(\RAM[117][3] ),
    .A2(\RAM[118][3] ),
    .A3(\RAM[119][3] ),
    .S0(net143),
    .S1(net90),
    .X(_0763_));
 sky130_fd_sc_hd__o21ba_1 _1246_ (.A1(_0533_),
    .A2(_0763_),
    .B1_N(_0531_),
    .X(_0764_));
 sky130_fd_sc_hd__mux4_1 _1247_ (.A0(\RAM[112][3] ),
    .A1(\RAM[113][3] ),
    .A2(\RAM[114][3] ),
    .A3(\RAM[115][3] ),
    .S0(net130),
    .S1(net80),
    .X(_0765_));
 sky130_fd_sc_hd__mux4_2 _1248_ (.A0(\RAM[120][3] ),
    .A1(\RAM[121][3] ),
    .A2(\RAM[122][3] ),
    .A3(\RAM[123][3] ),
    .S0(net136),
    .S1(net83),
    .X(_0766_));
 sky130_fd_sc_hd__mux4_2 _1249_ (.A0(\RAM[124][3] ),
    .A1(\RAM[125][3] ),
    .A2(\RAM[126][3] ),
    .A3(\RAM[127][3] ),
    .S0(net133),
    .S1(net81),
    .X(_0767_));
 sky130_fd_sc_hd__o22a_1 _1250_ (.A1(net24),
    .A2(_0766_),
    .B1(_0767_),
    .B2(net22),
    .X(_0768_));
 sky130_fd_sc_hd__o211a_1 _1251_ (.A1(net25),
    .A2(_0765_),
    .B1(_0768_),
    .C1(_0764_),
    .X(_0769_));
 sky130_fd_sc_hd__mux4_1 _1252_ (.A0(\RAM[100][3] ),
    .A1(\RAM[101][3] ),
    .A2(\RAM[102][3] ),
    .A3(\RAM[103][3] ),
    .S0(net133),
    .S1(net82),
    .X(_0770_));
 sky130_fd_sc_hd__mux4_1 _1253_ (.A0(\RAM[96][3] ),
    .A1(\RAM[97][3] ),
    .A2(\RAM[98][3] ),
    .A3(\RAM[99][3] ),
    .S0(net133),
    .S1(net81),
    .X(_0771_));
 sky130_fd_sc_hd__a22o_1 _1254_ (.A1(net29),
    .A2(_0770_),
    .B1(_0771_),
    .B2(net26),
    .X(_0772_));
 sky130_fd_sc_hd__mux4_1 _1255_ (.A0(\RAM[108][3] ),
    .A1(\RAM[109][3] ),
    .A2(\RAM[110][3] ),
    .A3(\RAM[111][3] ),
    .S0(net134),
    .S1(net82),
    .X(_0773_));
 sky130_fd_sc_hd__mux4_1 _1256_ (.A0(\RAM[104][3] ),
    .A1(\RAM[105][3] ),
    .A2(\RAM[106][3] ),
    .A3(\RAM[107][3] ),
    .S0(net134),
    .S1(net82),
    .X(_0774_));
 sky130_fd_sc_hd__o21a_1 _1257_ (.A1(net76),
    .A2(_0774_),
    .B1(net4),
    .X(_0775_));
 sky130_fd_sc_hd__or2_1 _1258_ (.A(net33),
    .B(_0773_),
    .X(_0776_));
 sky130_fd_sc_hd__a21o_1 _1259_ (.A1(_0775_),
    .A2(_0776_),
    .B1(_0772_),
    .X(_0777_));
 sky130_fd_sc_hd__a21oi_2 _1260_ (.A1(_0558_),
    .A2(_0777_),
    .B1(_0769_),
    .Y(_0778_));
 sky130_fd_sc_hd__mux4_2 _1261_ (.A0(\RAM[84][3] ),
    .A1(\RAM[85][3] ),
    .A2(\RAM[86][3] ),
    .A3(\RAM[87][3] ),
    .S0(net146),
    .S1(net92),
    .X(_0779_));
 sky130_fd_sc_hd__mux4_1 _1262_ (.A0(\RAM[88][3] ),
    .A1(\RAM[89][3] ),
    .A2(\RAM[90][3] ),
    .A3(\RAM[91][3] ),
    .S0(net141),
    .S1(net92),
    .X(_0780_));
 sky130_fd_sc_hd__a22o_1 _1263_ (.A1(net30),
    .A2(_0779_),
    .B1(_0780_),
    .B2(_0541_),
    .X(_0781_));
 sky130_fd_sc_hd__mux4_1 _1264_ (.A0(\RAM[92][3] ),
    .A1(\RAM[93][3] ),
    .A2(\RAM[94][3] ),
    .A3(\RAM[95][3] ),
    .S0(net139),
    .S1(net89),
    .X(_0782_));
 sky130_fd_sc_hd__mux4_2 _1265_ (.A0(\RAM[80][3] ),
    .A1(\RAM[81][3] ),
    .A2(\RAM[82][3] ),
    .A3(\RAM[83][3] ),
    .S0(net138),
    .S1(net86),
    .X(_0783_));
 sky130_fd_sc_hd__a22o_1 _1266_ (.A1(net23),
    .A2(_0782_),
    .B1(_0783_),
    .B2(net27),
    .X(_0784_));
 sky130_fd_sc_hd__nor2_1 _1267_ (.A(_0781_),
    .B(_0784_),
    .Y(_0785_));
 sky130_fd_sc_hd__o221a_1 _1268_ (.A1(_0516_),
    .A2(_0762_),
    .B1(_0785_),
    .B2(net21),
    .C1(_0778_),
    .X(_0786_));
 sky130_fd_sc_hd__mux2_1 _1269_ (.A0(\RAM[6][3] ),
    .A1(\RAM[7][3] ),
    .S(net145),
    .X(_0787_));
 sky130_fd_sc_hd__mux2_1 _1270_ (.A0(\RAM[4][3] ),
    .A1(\RAM[5][3] ),
    .S(net145),
    .X(_0788_));
 sky130_fd_sc_hd__a21o_1 _1271_ (.A1(_0513_),
    .A2(_0788_),
    .B1(net32),
    .X(_0789_));
 sky130_fd_sc_hd__a21oi_1 _1272_ (.A1(net93),
    .A2(_0787_),
    .B1(_0789_),
    .Y(_0790_));
 sky130_fd_sc_hd__mux4_1 _1273_ (.A0(\RAM[0][3] ),
    .A1(\RAM[1][3] ),
    .A2(\RAM[2][3] ),
    .A3(\RAM[3][3] ),
    .S0(net146),
    .S1(net92),
    .X(_0791_));
 sky130_fd_sc_hd__nor2_1 _1274_ (.A(net75),
    .B(_0791_),
    .Y(_0792_));
 sky130_fd_sc_hd__mux4_1 _1275_ (.A0(\RAM[8][3] ),
    .A1(\RAM[9][3] ),
    .A2(\RAM[10][3] ),
    .A3(\RAM[11][3] ),
    .S0(net146),
    .S1(net92),
    .X(_0793_));
 sky130_fd_sc_hd__mux2_1 _1276_ (.A0(\RAM[12][3] ),
    .A1(\RAM[13][3] ),
    .S(net144),
    .X(_0794_));
 sky130_fd_sc_hd__mux2_1 _1277_ (.A0(\RAM[14][3] ),
    .A1(\RAM[15][3] ),
    .S(net144),
    .X(_0795_));
 sky130_fd_sc_hd__a21o_1 _1278_ (.A1(_0513_),
    .A2(_0794_),
    .B1(net32),
    .X(_0796_));
 sky130_fd_sc_hd__a21oi_1 _1279_ (.A1(net93),
    .A2(_0795_),
    .B1(_0796_),
    .Y(_0797_));
 sky130_fd_sc_hd__o21ai_1 _1280_ (.A1(net75),
    .A2(_0793_),
    .B1(net72),
    .Y(_0798_));
 sky130_fd_sc_hd__o32a_1 _1281_ (.A1(net72),
    .A2(_0790_),
    .A3(_0792_),
    .B1(_0797_),
    .B2(_0798_),
    .X(_0799_));
 sky130_fd_sc_hd__nor2_1 _1282_ (.A(_0516_),
    .B(_0799_),
    .Y(_0800_));
 sky130_fd_sc_hd__mux4_1 _1283_ (.A0(\RAM[52][3] ),
    .A1(\RAM[53][3] ),
    .A2(\RAM[54][3] ),
    .A3(\RAM[55][3] ),
    .S0(net139),
    .S1(net89),
    .X(_0801_));
 sky130_fd_sc_hd__o21ba_1 _1284_ (.A1(net28),
    .A2(_0801_),
    .B1_N(_0531_),
    .X(_0802_));
 sky130_fd_sc_hd__mux4_1 _1285_ (.A0(\RAM[48][3] ),
    .A1(\RAM[49][3] ),
    .A2(\RAM[50][3] ),
    .A3(\RAM[51][3] ),
    .S0(net138),
    .S1(net86),
    .X(_0803_));
 sky130_fd_sc_hd__mux4_1 _1286_ (.A0(\RAM[56][3] ),
    .A1(\RAM[57][3] ),
    .A2(\RAM[58][3] ),
    .A3(\RAM[59][3] ),
    .S0(net131),
    .S1(net80),
    .X(_0804_));
 sky130_fd_sc_hd__mux4_1 _1287_ (.A0(\RAM[60][3] ),
    .A1(\RAM[61][3] ),
    .A2(\RAM[62][3] ),
    .A3(\RAM[63][3] ),
    .S0(net131),
    .S1(net79),
    .X(_0805_));
 sky130_fd_sc_hd__o22a_1 _1288_ (.A1(net24),
    .A2(_0804_),
    .B1(_0805_),
    .B2(net22),
    .X(_0806_));
 sky130_fd_sc_hd__o211a_1 _1289_ (.A1(net25),
    .A2(_0803_),
    .B1(_0806_),
    .C1(_0802_),
    .X(_0807_));
 sky130_fd_sc_hd__mux2_1 _1290_ (.A0(\RAM[40][3] ),
    .A1(\RAM[41][3] ),
    .S(net129),
    .X(_0808_));
 sky130_fd_sc_hd__or2_1 _1291_ (.A(net78),
    .B(_0808_),
    .X(_0809_));
 sky130_fd_sc_hd__mux2_1 _1292_ (.A0(\RAM[42][3] ),
    .A1(\RAM[43][3] ),
    .S(net129),
    .X(_0810_));
 sky130_fd_sc_hd__or2_1 _1293_ (.A(net35),
    .B(_0810_),
    .X(_0811_));
 sky130_fd_sc_hd__mux4_1 _1294_ (.A0(\RAM[32][3] ),
    .A1(\RAM[33][3] ),
    .A2(\RAM[34][3] ),
    .A3(\RAM[35][3] ),
    .S0(net128),
    .S1(net78),
    .X(_0812_));
 sky130_fd_sc_hd__a32o_1 _1295_ (.A1(_0541_),
    .A2(_0809_),
    .A3(_0811_),
    .B1(_0812_),
    .B2(net26),
    .X(_0813_));
 sky130_fd_sc_hd__mux4_2 _1296_ (.A0(\RAM[44][3] ),
    .A1(\RAM[45][3] ),
    .A2(\RAM[46][3] ),
    .A3(\RAM[47][3] ),
    .S0(net128),
    .S1(net77),
    .X(_0814_));
 sky130_fd_sc_hd__mux4_1 _1297_ (.A0(\RAM[36][3] ),
    .A1(\RAM[37][3] ),
    .A2(\RAM[38][3] ),
    .A3(\RAM[39][3] ),
    .S0(net128),
    .S1(net77),
    .X(_0815_));
 sky130_fd_sc_hd__a22o_1 _1298_ (.A1(net23),
    .A2(_0814_),
    .B1(_0815_),
    .B2(net29),
    .X(_0816_));
 sky130_fd_sc_hd__o21a_1 _1299_ (.A1(_0813_),
    .A2(_0816_),
    .B1(_0558_),
    .X(_0817_));
 sky130_fd_sc_hd__mux4_1 _1300_ (.A0(\RAM[20][3] ),
    .A1(\RAM[21][3] ),
    .A2(\RAM[22][3] ),
    .A3(\RAM[23][3] ),
    .S0(net141),
    .S1(net88),
    .X(_0818_));
 sky130_fd_sc_hd__mux4_1 _1301_ (.A0(\RAM[24][3] ),
    .A1(\RAM[25][3] ),
    .A2(\RAM[26][3] ),
    .A3(\RAM[27][3] ),
    .S0(net140),
    .S1(net88),
    .X(_0819_));
 sky130_fd_sc_hd__a22o_1 _1302_ (.A1(net30),
    .A2(_0818_),
    .B1(_0819_),
    .B2(_0541_),
    .X(_0820_));
 sky130_fd_sc_hd__mux4_1 _1303_ (.A0(\RAM[28][3] ),
    .A1(\RAM[29][3] ),
    .A2(\RAM[30][3] ),
    .A3(\RAM[31][3] ),
    .S0(net140),
    .S1(net87),
    .X(_0821_));
 sky130_fd_sc_hd__mux4_1 _1304_ (.A0(\RAM[16][3] ),
    .A1(\RAM[17][3] ),
    .A2(\RAM[18][3] ),
    .A3(\RAM[19][3] ),
    .S0(net141),
    .S1(net87),
    .X(_0822_));
 sky130_fd_sc_hd__a22o_1 _1305_ (.A1(_0544_),
    .A2(_0821_),
    .B1(_0822_),
    .B2(net27),
    .X(_0823_));
 sky130_fd_sc_hd__o21ba_1 _1306_ (.A1(_0820_),
    .A2(_0823_),
    .B1_N(net21),
    .X(_0824_));
 sky130_fd_sc_hd__or4_1 _1307_ (.A(net7),
    .B(_0807_),
    .C(_0817_),
    .D(_0824_),
    .X(_0825_));
 sky130_fd_sc_hd__o2bb2a_2 _1308_ (.A1_N(net7),
    .A2_N(_0786_),
    .B1(_0800_),
    .B2(_0825_),
    .X(net16));
 sky130_fd_sc_hd__nor2_8 _1309_ (.A(_0533_),
    .B(_0535_),
    .Y(_0826_));
 sky130_fd_sc_hd__or2_4 _1310_ (.A(_0533_),
    .B(_0535_),
    .X(_0827_));
 sky130_fd_sc_hd__nand2_8 _1311_ (.A(net7),
    .B(net12),
    .Y(_0828_));
 sky130_fd_sc_hd__nor2_8 _1312_ (.A(_0516_),
    .B(_0828_),
    .Y(_0829_));
 sky130_fd_sc_hd__or2_4 _1313_ (.A(_0516_),
    .B(_0828_),
    .X(_0830_));
 sky130_fd_sc_hd__nor2_2 _1314_ (.A(_0827_),
    .B(net20),
    .Y(_0831_));
 sky130_fd_sc_hd__mux2_1 _1315_ (.A0(\RAM[69][0] ),
    .A1(net66),
    .S(_0831_),
    .X(_0000_));
 sky130_fd_sc_hd__mux2_1 _1316_ (.A0(\RAM[69][1] ),
    .A1(net49),
    .S(_0831_),
    .X(_0001_));
 sky130_fd_sc_hd__mux2_1 _1317_ (.A0(\RAM[69][2] ),
    .A1(net125),
    .S(_0831_),
    .X(_0002_));
 sky130_fd_sc_hd__mux2_1 _1318_ (.A0(\RAM[69][3] ),
    .A1(net105),
    .S(_0831_),
    .X(_0003_));
 sky130_fd_sc_hd__nor2_8 _1319_ (.A(_0535_),
    .B(net24),
    .Y(_0832_));
 sky130_fd_sc_hd__or2_4 _1320_ (.A(_0535_),
    .B(_0542_),
    .X(_0833_));
 sky130_fd_sc_hd__nor2_8 _1321_ (.A(_0561_),
    .B(_0828_),
    .Y(_0834_));
 sky130_fd_sc_hd__or2_4 _1322_ (.A(_0561_),
    .B(_0828_),
    .X(_0835_));
 sky130_fd_sc_hd__nand2_2 _1323_ (.A(_0832_),
    .B(_0834_),
    .Y(_0836_));
 sky130_fd_sc_hd__mux2_1 _1324_ (.A0(net58),
    .A1(\RAM[89][0] ),
    .S(_0836_),
    .X(_0004_));
 sky130_fd_sc_hd__mux2_1 _1325_ (.A0(net49),
    .A1(\RAM[89][1] ),
    .S(_0836_),
    .X(_0005_));
 sky130_fd_sc_hd__mux2_1 _1326_ (.A0(net123),
    .A1(\RAM[89][2] ),
    .S(_0836_),
    .X(_0006_));
 sky130_fd_sc_hd__mux2_1 _1327_ (.A0(net104),
    .A1(\RAM[89][3] ),
    .S(_0836_),
    .X(_0007_));
 sky130_fd_sc_hd__nor2_8 _1328_ (.A(_0534_),
    .B(_0542_),
    .Y(_0837_));
 sky130_fd_sc_hd__nand2b_4 _1329_ (.A_N(net7),
    .B(net12),
    .Y(_0838_));
 sky130_fd_sc_hd__nor2_8 _1330_ (.A(_0531_),
    .B(_0838_),
    .Y(_0839_));
 sky130_fd_sc_hd__or2_4 _1331_ (.A(_0531_),
    .B(_0838_),
    .X(_0840_));
 sky130_fd_sc_hd__nand2_2 _1332_ (.A(_0837_),
    .B(_0839_),
    .Y(_0841_));
 sky130_fd_sc_hd__mux2_1 _1333_ (.A0(net55),
    .A1(\RAM[59][0] ),
    .S(_0841_),
    .X(_0008_));
 sky130_fd_sc_hd__mux2_1 _1334_ (.A0(net38),
    .A1(\RAM[59][1] ),
    .S(_0841_),
    .X(_0009_));
 sky130_fd_sc_hd__mux2_1 _1335_ (.A0(net112),
    .A1(\RAM[59][2] ),
    .S(_0841_),
    .X(_0010_));
 sky130_fd_sc_hd__mux2_1 _1336_ (.A0(net97),
    .A1(\RAM[59][3] ),
    .S(_0841_),
    .X(_0011_));
 sky130_fd_sc_hd__or2_4 _1337_ (.A(_0535_),
    .B(net25),
    .X(_0842_));
 sky130_fd_sc_hd__nor2_4 _1338_ (.A(_0840_),
    .B(_0842_),
    .Y(_0843_));
 sky130_fd_sc_hd__mux2_1 _1339_ (.A0(\RAM[49][0] ),
    .A1(net54),
    .S(_0843_),
    .X(_0012_));
 sky130_fd_sc_hd__mux2_1 _1340_ (.A0(\RAM[49][1] ),
    .A1(net38),
    .S(_0843_),
    .X(_0013_));
 sky130_fd_sc_hd__mux2_1 _1341_ (.A0(\RAM[49][2] ),
    .A1(net115),
    .S(_0843_),
    .X(_0014_));
 sky130_fd_sc_hd__mux2_1 _1342_ (.A0(\RAM[49][3] ),
    .A1(net101),
    .S(_0843_),
    .X(_0015_));
 sky130_fd_sc_hd__nor2_8 _1343_ (.A(net28),
    .B(_0534_),
    .Y(_0844_));
 sky130_fd_sc_hd__nor2_8 _1344_ (.A(_0559_),
    .B(_0838_),
    .Y(_0845_));
 sky130_fd_sc_hd__or2_4 _1345_ (.A(_0559_),
    .B(_0838_),
    .X(_0846_));
 sky130_fd_sc_hd__nand2_2 _1346_ (.A(_0844_),
    .B(_0845_),
    .Y(_0847_));
 sky130_fd_sc_hd__mux2_1 _1347_ (.A0(net53),
    .A1(\RAM[39][0] ),
    .S(_0847_),
    .X(_0016_));
 sky130_fd_sc_hd__mux2_1 _1348_ (.A0(net36),
    .A1(\RAM[39][1] ),
    .S(_0847_),
    .X(_0017_));
 sky130_fd_sc_hd__mux2_1 _1349_ (.A0(net111),
    .A1(\RAM[39][2] ),
    .S(_0847_),
    .X(_0018_));
 sky130_fd_sc_hd__mux2_1 _1350_ (.A0(net95),
    .A1(\RAM[39][3] ),
    .S(_0847_),
    .X(_0019_));
 sky130_fd_sc_hd__nor2_8 _1351_ (.A(_0534_),
    .B(_0539_),
    .Y(_0848_));
 sky130_fd_sc_hd__or2_4 _1352_ (.A(_0534_),
    .B(_0539_),
    .X(_0849_));
 sky130_fd_sc_hd__nor2_8 _1353_ (.A(net21),
    .B(_0838_),
    .Y(_0850_));
 sky130_fd_sc_hd__or2_4 _1354_ (.A(net21),
    .B(_0838_),
    .X(_0851_));
 sky130_fd_sc_hd__nor2_4 _1355_ (.A(_0849_),
    .B(net18),
    .Y(_0852_));
 sky130_fd_sc_hd__mux2_1 _1356_ (.A0(\RAM[19][0] ),
    .A1(net57),
    .S(_0852_),
    .X(_0020_));
 sky130_fd_sc_hd__mux2_1 _1357_ (.A0(\RAM[19][1] ),
    .A1(net46),
    .S(_0852_),
    .X(_0021_));
 sky130_fd_sc_hd__mux2_1 _1358_ (.A0(\RAM[19][2] ),
    .A1(net116),
    .S(_0852_),
    .X(_0022_));
 sky130_fd_sc_hd__mux2_1 _1359_ (.A0(\RAM[19][3] ),
    .A1(net103),
    .S(_0852_),
    .X(_0023_));
 sky130_fd_sc_hd__nor2_8 _1360_ (.A(_0534_),
    .B(_0545_),
    .Y(_0853_));
 sky130_fd_sc_hd__nand2_2 _1361_ (.A(_0829_),
    .B(_0853_),
    .Y(_0854_));
 sky130_fd_sc_hd__mux2_1 _1362_ (.A0(net63),
    .A1(\RAM[79][0] ),
    .S(_0854_),
    .X(_0024_));
 sky130_fd_sc_hd__mux2_1 _1363_ (.A0(net42),
    .A1(\RAM[79][1] ),
    .S(_0854_),
    .X(_0025_));
 sky130_fd_sc_hd__mux2_1 _1364_ (.A0(net125),
    .A1(\RAM[79][2] ),
    .S(_0854_),
    .X(_0026_));
 sky130_fd_sc_hd__mux2_1 _1365_ (.A0(net105),
    .A1(\RAM[79][3] ),
    .S(_0854_),
    .X(_0027_));
 sky130_fd_sc_hd__nor2_8 _1366_ (.A(_0535_),
    .B(net22),
    .Y(_0855_));
 sky130_fd_sc_hd__nand2_4 _1367_ (.A(_0850_),
    .B(_0855_),
    .Y(_0856_));
 sky130_fd_sc_hd__mux2_1 _1368_ (.A0(net57),
    .A1(\RAM[29][0] ),
    .S(_0856_),
    .X(_0028_));
 sky130_fd_sc_hd__mux2_1 _1369_ (.A0(net46),
    .A1(\RAM[29][1] ),
    .S(_0856_),
    .X(_0029_));
 sky130_fd_sc_hd__mux2_1 _1370_ (.A0(net116),
    .A1(\RAM[29][2] ),
    .S(_0856_),
    .X(_0030_));
 sky130_fd_sc_hd__mux2_1 _1371_ (.A0(net103),
    .A1(\RAM[29][3] ),
    .S(_0856_),
    .X(_0031_));
 sky130_fd_sc_hd__nor2_8 _1372_ (.A(_0559_),
    .B(_0828_),
    .Y(_0857_));
 sky130_fd_sc_hd__or2_4 _1373_ (.A(_0559_),
    .B(_0828_),
    .X(_0858_));
 sky130_fd_sc_hd__nand2_2 _1374_ (.A(_0848_),
    .B(_0857_),
    .Y(_0859_));
 sky130_fd_sc_hd__mux2_1 _1375_ (.A0(net60),
    .A1(\RAM[99][0] ),
    .S(_0859_),
    .X(_0032_));
 sky130_fd_sc_hd__mux2_1 _1376_ (.A0(net40),
    .A1(\RAM[99][1] ),
    .S(_0859_),
    .X(_0033_));
 sky130_fd_sc_hd__mux2_1 _1377_ (.A0(net119),
    .A1(\RAM[99][2] ),
    .S(_0859_),
    .X(_0034_));
 sky130_fd_sc_hd__mux2_1 _1378_ (.A0(net98),
    .A1(\RAM[99][3] ),
    .S(_0859_),
    .X(_0035_));
 sky130_fd_sc_hd__nand2_2 _1379_ (.A(_0855_),
    .B(_0857_),
    .Y(_0860_));
 sky130_fd_sc_hd__mux2_1 _1380_ (.A0(net62),
    .A1(\RAM[109][0] ),
    .S(_0860_),
    .X(_0036_));
 sky130_fd_sc_hd__mux2_1 _1381_ (.A0(net40),
    .A1(\RAM[109][1] ),
    .S(_0860_),
    .X(_0037_));
 sky130_fd_sc_hd__mux2_1 _1382_ (.A0(net121),
    .A1(\RAM[109][2] ),
    .S(_0860_),
    .X(_0038_));
 sky130_fd_sc_hd__mux2_1 _1383_ (.A0(net98),
    .A1(\RAM[109][3] ),
    .S(_0860_),
    .X(_0039_));
 sky130_fd_sc_hd__nor2_8 _1384_ (.A(_0531_),
    .B(_0828_),
    .Y(_0861_));
 sky130_fd_sc_hd__or2_4 _1385_ (.A(_0531_),
    .B(_0828_),
    .X(_0862_));
 sky130_fd_sc_hd__nand2_2 _1386_ (.A(_0844_),
    .B(_0861_),
    .Y(_0863_));
 sky130_fd_sc_hd__mux2_1 _1387_ (.A0(net60),
    .A1(\RAM[119][0] ),
    .S(_0863_),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_1 _1388_ (.A0(net42),
    .A1(\RAM[119][1] ),
    .S(_0863_),
    .X(_0041_));
 sky130_fd_sc_hd__mux2_1 _1389_ (.A0(net119),
    .A1(\RAM[119][2] ),
    .S(_0863_),
    .X(_0042_));
 sky130_fd_sc_hd__mux2_1 _1390_ (.A0(net105),
    .A1(\RAM[119][3] ),
    .S(_0863_),
    .X(_0043_));
 sky130_fd_sc_hd__nand2_2 _1391_ (.A(_0853_),
    .B(_0861_),
    .Y(_0864_));
 sky130_fd_sc_hd__mux2_1 _1392_ (.A0(net56),
    .A1(\RAM[127][0] ),
    .S(_0864_),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _1393_ (.A0(net37),
    .A1(\RAM[127][1] ),
    .S(_0864_),
    .X(_0045_));
 sky130_fd_sc_hd__mux2_1 _1394_ (.A0(net113),
    .A1(\RAM[127][2] ),
    .S(_0864_),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_1 _1395_ (.A0(net96),
    .A1(\RAM[127][3] ),
    .S(_0864_),
    .X(_0047_));
 sky130_fd_sc_hd__or3_4 _1396_ (.A(net130),
    .B(net80),
    .C(net22),
    .X(_0865_));
 sky130_fd_sc_hd__nor2_8 _1397_ (.A(_0516_),
    .B(_0838_),
    .Y(_0866_));
 sky130_fd_sc_hd__or2_4 _1398_ (.A(_0516_),
    .B(_0838_),
    .X(_0867_));
 sky130_fd_sc_hd__nor2_2 _1399_ (.A(_0865_),
    .B(net17),
    .Y(_0868_));
 sky130_fd_sc_hd__mux2_1 _1400_ (.A0(\RAM[12][0] ),
    .A1(net66),
    .S(_0868_),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _1401_ (.A0(\RAM[12][1] ),
    .A1(net51),
    .S(_0868_),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_1 _1402_ (.A0(\RAM[12][2] ),
    .A1(net124),
    .S(_0868_),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _1403_ (.A0(\RAM[12][3] ),
    .A1(net107),
    .S(_0868_),
    .X(_0051_));
 sky130_fd_sc_hd__nand2_4 _1404_ (.A(_0855_),
    .B(_0866_),
    .Y(_0869_));
 sky130_fd_sc_hd__mux2_1 _1405_ (.A0(net66),
    .A1(\RAM[13][0] ),
    .S(_0869_),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _1406_ (.A0(net49),
    .A1(\RAM[13][1] ),
    .S(_0869_),
    .X(_0053_));
 sky130_fd_sc_hd__mux2_1 _1407_ (.A0(net124),
    .A1(\RAM[13][2] ),
    .S(_0869_),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _1408_ (.A0(net107),
    .A1(\RAM[13][3] ),
    .S(_0869_),
    .X(_0055_));
 sky130_fd_sc_hd__and3b_4 _1409_ (.A_N(net143),
    .B(net90),
    .C(net23),
    .X(_0870_));
 sky130_fd_sc_hd__nand2_2 _1410_ (.A(_0866_),
    .B(_0870_),
    .Y(_0871_));
 sky130_fd_sc_hd__mux2_1 _1411_ (.A0(net66),
    .A1(\RAM[14][0] ),
    .S(_0871_),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _1412_ (.A0(net50),
    .A1(\RAM[14][1] ),
    .S(_0871_),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _1413_ (.A0(net124),
    .A1(\RAM[14][2] ),
    .S(_0871_),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_1 _1414_ (.A0(net107),
    .A1(\RAM[14][3] ),
    .S(_0871_),
    .X(_0059_));
 sky130_fd_sc_hd__and2_2 _1415_ (.A(_0853_),
    .B(_0866_),
    .X(_0872_));
 sky130_fd_sc_hd__mux2_1 _1416_ (.A0(\RAM[15][0] ),
    .A1(net66),
    .S(_0872_),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _1417_ (.A0(\RAM[15][1] ),
    .A1(net50),
    .S(_0872_),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _1418_ (.A0(\RAM[15][2] ),
    .A1(net124),
    .S(_0872_),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _1419_ (.A0(\RAM[15][3] ),
    .A1(net107),
    .S(_0872_),
    .X(_0063_));
 sky130_fd_sc_hd__or3_4 _1420_ (.A(net132),
    .B(net80),
    .C(net25),
    .X(_0873_));
 sky130_fd_sc_hd__nor2_4 _1421_ (.A(net18),
    .B(_0873_),
    .Y(_0874_));
 sky130_fd_sc_hd__mux2_1 _1422_ (.A0(\RAM[16][0] ),
    .A1(net57),
    .S(_0874_),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _1423_ (.A0(\RAM[16][1] ),
    .A1(net46),
    .S(_0874_),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _1424_ (.A0(\RAM[16][2] ),
    .A1(net116),
    .S(_0874_),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_1 _1425_ (.A0(\RAM[16][3] ),
    .A1(net103),
    .S(_0874_),
    .X(_0067_));
 sky130_fd_sc_hd__nor2_4 _1426_ (.A(_0842_),
    .B(net18),
    .Y(_0875_));
 sky130_fd_sc_hd__mux2_1 _1427_ (.A0(\RAM[17][0] ),
    .A1(net57),
    .S(_0875_),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _1428_ (.A0(\RAM[17][1] ),
    .A1(net46),
    .S(_0875_),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_1 _1429_ (.A0(\RAM[17][2] ),
    .A1(net116),
    .S(_0875_),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _1430_ (.A0(\RAM[17][3] ),
    .A1(net103),
    .S(_0875_),
    .X(_0071_));
 sky130_fd_sc_hd__or3_4 _1431_ (.A(net136),
    .B(net35),
    .C(_0539_),
    .X(_0876_));
 sky130_fd_sc_hd__nor2_4 _1432_ (.A(net18),
    .B(_0876_),
    .Y(_0877_));
 sky130_fd_sc_hd__mux2_1 _1433_ (.A0(\RAM[18][0] ),
    .A1(net57),
    .S(_0877_),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_1 _1434_ (.A0(\RAM[18][1] ),
    .A1(net46),
    .S(_0877_),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _1435_ (.A0(\RAM[18][2] ),
    .A1(net116),
    .S(_0877_),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _1436_ (.A0(\RAM[18][3] ),
    .A1(net103),
    .S(_0877_),
    .X(_0075_));
 sky130_fd_sc_hd__nor2_4 _1437_ (.A(_0842_),
    .B(net17),
    .Y(_0878_));
 sky130_fd_sc_hd__mux2_1 _1438_ (.A0(\RAM[1][0] ),
    .A1(net64),
    .S(_0878_),
    .X(_0076_));
 sky130_fd_sc_hd__mux2_1 _1439_ (.A0(\RAM[1][1] ),
    .A1(net51),
    .S(_0878_),
    .X(_0077_));
 sky130_fd_sc_hd__mux2_1 _1440_ (.A0(\RAM[1][2] ),
    .A1(net124),
    .S(_0878_),
    .X(_0078_));
 sky130_fd_sc_hd__mux2_1 _1441_ (.A0(\RAM[1][3] ),
    .A1(net106),
    .S(_0878_),
    .X(_0079_));
 sky130_fd_sc_hd__or3_4 _1442_ (.A(net130),
    .B(net80),
    .C(net28),
    .X(_0879_));
 sky130_fd_sc_hd__nor2_2 _1443_ (.A(net18),
    .B(_0879_),
    .Y(_0880_));
 sky130_fd_sc_hd__mux2_1 _1444_ (.A0(\RAM[20][0] ),
    .A1(net58),
    .S(_0880_),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _1445_ (.A0(\RAM[20][1] ),
    .A1(net46),
    .S(_0880_),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_1 _1446_ (.A0(\RAM[20][2] ),
    .A1(net117),
    .S(_0880_),
    .X(_0082_));
 sky130_fd_sc_hd__mux2_1 _1447_ (.A0(\RAM[20][3] ),
    .A1(net104),
    .S(_0880_),
    .X(_0083_));
 sky130_fd_sc_hd__nor2_2 _1448_ (.A(_0827_),
    .B(net18),
    .Y(_0881_));
 sky130_fd_sc_hd__mux2_1 _1449_ (.A0(\RAM[21][0] ),
    .A1(net58),
    .S(_0881_),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_1 _1450_ (.A0(\RAM[21][1] ),
    .A1(net47),
    .S(_0881_),
    .X(_0085_));
 sky130_fd_sc_hd__mux2_1 _1451_ (.A0(\RAM[21][2] ),
    .A1(net117),
    .S(_0881_),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_1 _1452_ (.A0(\RAM[21][3] ),
    .A1(net104),
    .S(_0881_),
    .X(_0087_));
 sky130_fd_sc_hd__or3_4 _1453_ (.A(net139),
    .B(net35),
    .C(net28),
    .X(_0882_));
 sky130_fd_sc_hd__nor2_2 _1454_ (.A(net18),
    .B(_0882_),
    .Y(_0883_));
 sky130_fd_sc_hd__mux2_1 _1455_ (.A0(\RAM[22][0] ),
    .A1(net58),
    .S(_0883_),
    .X(_0088_));
 sky130_fd_sc_hd__mux2_1 _1456_ (.A0(\RAM[22][1] ),
    .A1(net47),
    .S(_0883_),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _1457_ (.A0(\RAM[22][2] ),
    .A1(net117),
    .S(_0883_),
    .X(_0090_));
 sky130_fd_sc_hd__mux2_1 _1458_ (.A0(\RAM[22][3] ),
    .A1(net104),
    .S(_0883_),
    .X(_0091_));
 sky130_fd_sc_hd__nand2_2 _1459_ (.A(_0844_),
    .B(_0850_),
    .Y(_0884_));
 sky130_fd_sc_hd__mux2_1 _1460_ (.A0(net59),
    .A1(\RAM[23][0] ),
    .S(_0884_),
    .X(_0092_));
 sky130_fd_sc_hd__mux2_1 _1461_ (.A0(net47),
    .A1(\RAM[23][1] ),
    .S(_0884_),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _1462_ (.A0(net117),
    .A1(\RAM[23][2] ),
    .S(_0884_),
    .X(_0094_));
 sky130_fd_sc_hd__mux2_1 _1463_ (.A0(net104),
    .A1(\RAM[23][3] ),
    .S(_0884_),
    .X(_0095_));
 sky130_fd_sc_hd__or3_4 _1464_ (.A(net130),
    .B(net83),
    .C(net24),
    .X(_0885_));
 sky130_fd_sc_hd__nor2_2 _1465_ (.A(net18),
    .B(_0885_),
    .Y(_0886_));
 sky130_fd_sc_hd__mux2_1 _1466_ (.A0(\RAM[24][0] ),
    .A1(net59),
    .S(_0886_),
    .X(_0096_));
 sky130_fd_sc_hd__mux2_1 _1467_ (.A0(\RAM[24][1] ),
    .A1(net47),
    .S(_0886_),
    .X(_0097_));
 sky130_fd_sc_hd__mux2_1 _1468_ (.A0(\RAM[24][2] ),
    .A1(net117),
    .S(_0886_),
    .X(_0098_));
 sky130_fd_sc_hd__mux2_1 _1469_ (.A0(\RAM[24][3] ),
    .A1(net104),
    .S(_0886_),
    .X(_0099_));
 sky130_fd_sc_hd__nor2_4 _1470_ (.A(_0833_),
    .B(_0851_),
    .Y(_0887_));
 sky130_fd_sc_hd__mux2_1 _1471_ (.A0(\RAM[25][0] ),
    .A1(net59),
    .S(_0887_),
    .X(_0100_));
 sky130_fd_sc_hd__mux2_1 _1472_ (.A0(\RAM[25][1] ),
    .A1(net47),
    .S(_0887_),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _1473_ (.A0(\RAM[25][2] ),
    .A1(net118),
    .S(_0887_),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_1 _1474_ (.A0(\RAM[25][3] ),
    .A1(net104),
    .S(_0887_),
    .X(_0103_));
 sky130_fd_sc_hd__or3_4 _1475_ (.A(net136),
    .B(net35),
    .C(_0542_),
    .X(_0888_));
 sky130_fd_sc_hd__nor2_2 _1476_ (.A(net18),
    .B(_0888_),
    .Y(_0889_));
 sky130_fd_sc_hd__mux2_1 _1477_ (.A0(\RAM[26][0] ),
    .A1(net57),
    .S(_0889_),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _1478_ (.A0(\RAM[26][1] ),
    .A1(net46),
    .S(_0889_),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _1479_ (.A0(\RAM[26][2] ),
    .A1(net116),
    .S(_0889_),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _1480_ (.A0(\RAM[26][3] ),
    .A1(net103),
    .S(_0889_),
    .X(_0107_));
 sky130_fd_sc_hd__nand2_4 _1481_ (.A(_0837_),
    .B(_0850_),
    .Y(_0890_));
 sky130_fd_sc_hd__mux2_1 _1482_ (.A0(net59),
    .A1(\RAM[27][0] ),
    .S(_0890_),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _1483_ (.A0(net47),
    .A1(\RAM[27][1] ),
    .S(_0890_),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _1484_ (.A0(net116),
    .A1(\RAM[27][2] ),
    .S(_0890_),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_1 _1485_ (.A0(net103),
    .A1(\RAM[27][3] ),
    .S(_0890_),
    .X(_0111_));
 sky130_fd_sc_hd__nor2_2 _1486_ (.A(net18),
    .B(_0865_),
    .Y(_0891_));
 sky130_fd_sc_hd__mux2_1 _1487_ (.A0(\RAM[28][0] ),
    .A1(net59),
    .S(_0891_),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _1488_ (.A0(\RAM[28][1] ),
    .A1(net46),
    .S(_0891_),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _1489_ (.A0(\RAM[28][2] ),
    .A1(net118),
    .S(_0891_),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_1 _1490_ (.A0(\RAM[28][3] ),
    .A1(net103),
    .S(_0891_),
    .X(_0115_));
 sky130_fd_sc_hd__nor2_4 _1491_ (.A(net17),
    .B(_0876_),
    .Y(_0892_));
 sky130_fd_sc_hd__mux2_1 _1492_ (.A0(\RAM[2][0] ),
    .A1(net64),
    .S(_0892_),
    .X(_0116_));
 sky130_fd_sc_hd__mux2_1 _1493_ (.A0(\RAM[2][1] ),
    .A1(net51),
    .S(_0892_),
    .X(_0117_));
 sky130_fd_sc_hd__mux2_1 _1494_ (.A0(\RAM[2][2] ),
    .A1(net123),
    .S(_0892_),
    .X(_0118_));
 sky130_fd_sc_hd__mux2_1 _1495_ (.A0(\RAM[2][3] ),
    .A1(net106),
    .S(_0892_),
    .X(_0119_));
 sky130_fd_sc_hd__nand2_4 _1496_ (.A(_0850_),
    .B(_0870_),
    .Y(_0893_));
 sky130_fd_sc_hd__mux2_1 _1497_ (.A0(net59),
    .A1(\RAM[30][0] ),
    .S(_0893_),
    .X(_0120_));
 sky130_fd_sc_hd__mux2_1 _1498_ (.A0(net46),
    .A1(\RAM[30][1] ),
    .S(_0893_),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _1499_ (.A0(net118),
    .A1(\RAM[30][2] ),
    .S(_0893_),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _1500_ (.A0(net103),
    .A1(\RAM[30][3] ),
    .S(_0893_),
    .X(_0123_));
 sky130_fd_sc_hd__nand2_4 _1501_ (.A(_0850_),
    .B(_0853_),
    .Y(_0894_));
 sky130_fd_sc_hd__mux2_1 _1502_ (.A0(net59),
    .A1(\RAM[31][0] ),
    .S(_0894_),
    .X(_0124_));
 sky130_fd_sc_hd__mux2_1 _1503_ (.A0(net46),
    .A1(\RAM[31][1] ),
    .S(_0894_),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_1 _1504_ (.A0(net118),
    .A1(\RAM[31][2] ),
    .S(_0894_),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_1 _1505_ (.A0(net103),
    .A1(\RAM[31][3] ),
    .S(_0894_),
    .X(_0127_));
 sky130_fd_sc_hd__nor2_2 _1506_ (.A(net19),
    .B(_0873_),
    .Y(_0895_));
 sky130_fd_sc_hd__mux2_1 _1507_ (.A0(\RAM[32][0] ),
    .A1(net56),
    .S(_0895_),
    .X(_0128_));
 sky130_fd_sc_hd__mux2_1 _1508_ (.A0(\RAM[32][1] ),
    .A1(net37),
    .S(_0895_),
    .X(_0129_));
 sky130_fd_sc_hd__mux2_1 _1509_ (.A0(\RAM[32][2] ),
    .A1(net113),
    .S(_0895_),
    .X(_0130_));
 sky130_fd_sc_hd__mux2_1 _1510_ (.A0(\RAM[32][3] ),
    .A1(net96),
    .S(_0895_),
    .X(_0131_));
 sky130_fd_sc_hd__nor2_2 _1511_ (.A(_0842_),
    .B(net19),
    .Y(_0896_));
 sky130_fd_sc_hd__mux2_1 _1512_ (.A0(\RAM[33][0] ),
    .A1(net53),
    .S(_0896_),
    .X(_0132_));
 sky130_fd_sc_hd__mux2_1 _1513_ (.A0(\RAM[33][1] ),
    .A1(net36),
    .S(_0896_),
    .X(_0133_));
 sky130_fd_sc_hd__mux2_1 _1514_ (.A0(\RAM[33][2] ),
    .A1(net111),
    .S(_0896_),
    .X(_0134_));
 sky130_fd_sc_hd__mux2_1 _1515_ (.A0(\RAM[33][3] ),
    .A1(net95),
    .S(_0896_),
    .X(_0135_));
 sky130_fd_sc_hd__nor2_2 _1516_ (.A(net19),
    .B(_0876_),
    .Y(_0897_));
 sky130_fd_sc_hd__mux2_1 _1517_ (.A0(\RAM[34][0] ),
    .A1(net53),
    .S(_0897_),
    .X(_0136_));
 sky130_fd_sc_hd__mux2_1 _1518_ (.A0(\RAM[34][1] ),
    .A1(net36),
    .S(_0897_),
    .X(_0137_));
 sky130_fd_sc_hd__mux2_1 _1519_ (.A0(\RAM[34][2] ),
    .A1(net111),
    .S(_0897_),
    .X(_0138_));
 sky130_fd_sc_hd__mux2_1 _1520_ (.A0(\RAM[34][3] ),
    .A1(net95),
    .S(_0897_),
    .X(_0139_));
 sky130_fd_sc_hd__nor2_2 _1521_ (.A(net19),
    .B(_0849_),
    .Y(_0898_));
 sky130_fd_sc_hd__mux2_1 _1522_ (.A0(\RAM[35][0] ),
    .A1(net54),
    .S(_0898_),
    .X(_0140_));
 sky130_fd_sc_hd__mux2_1 _1523_ (.A0(\RAM[35][1] ),
    .A1(net36),
    .S(_0898_),
    .X(_0141_));
 sky130_fd_sc_hd__mux2_1 _1524_ (.A0(\RAM[35][2] ),
    .A1(net111),
    .S(_0898_),
    .X(_0142_));
 sky130_fd_sc_hd__mux2_1 _1525_ (.A0(\RAM[35][3] ),
    .A1(net95),
    .S(_0898_),
    .X(_0143_));
 sky130_fd_sc_hd__nor2_4 _1526_ (.A(net19),
    .B(_0879_),
    .Y(_0899_));
 sky130_fd_sc_hd__mux2_1 _1527_ (.A0(\RAM[36][0] ),
    .A1(net53),
    .S(_0899_),
    .X(_0144_));
 sky130_fd_sc_hd__mux2_1 _1528_ (.A0(\RAM[36][1] ),
    .A1(net36),
    .S(_0899_),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _1529_ (.A0(\RAM[36][2] ),
    .A1(net111),
    .S(_0899_),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_1 _1530_ (.A0(\RAM[36][3] ),
    .A1(net95),
    .S(_0899_),
    .X(_0147_));
 sky130_fd_sc_hd__nor2_4 _1531_ (.A(_0827_),
    .B(_0846_),
    .Y(_0900_));
 sky130_fd_sc_hd__mux2_1 _1532_ (.A0(\RAM[37][0] ),
    .A1(net53),
    .S(_0900_),
    .X(_0148_));
 sky130_fd_sc_hd__mux2_1 _1533_ (.A0(\RAM[37][1] ),
    .A1(net36),
    .S(_0900_),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_1 _1534_ (.A0(\RAM[37][2] ),
    .A1(net111),
    .S(_0900_),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_1 _1535_ (.A0(\RAM[37][3] ),
    .A1(net97),
    .S(_0900_),
    .X(_0151_));
 sky130_fd_sc_hd__nor2_4 _1536_ (.A(net19),
    .B(_0882_),
    .Y(_0901_));
 sky130_fd_sc_hd__mux2_1 _1537_ (.A0(\RAM[38][0] ),
    .A1(net53),
    .S(_0901_),
    .X(_0152_));
 sky130_fd_sc_hd__mux2_1 _1538_ (.A0(\RAM[38][1] ),
    .A1(net37),
    .S(_0901_),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _1539_ (.A0(\RAM[38][2] ),
    .A1(net111),
    .S(_0901_),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_1 _1540_ (.A0(\RAM[38][3] ),
    .A1(net95),
    .S(_0901_),
    .X(_0155_));
 sky130_fd_sc_hd__nor2_2 _1541_ (.A(_0849_),
    .B(net17),
    .Y(_0902_));
 sky130_fd_sc_hd__mux2_1 _1542_ (.A0(\RAM[3][0] ),
    .A1(net65),
    .S(_0902_),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _1543_ (.A0(\RAM[3][1] ),
    .A1(net51),
    .S(_0902_),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_1 _1544_ (.A0(\RAM[3][2] ),
    .A1(net123),
    .S(_0902_),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_1 _1545_ (.A0(\RAM[3][3] ),
    .A1(net106),
    .S(_0902_),
    .X(_0159_));
 sky130_fd_sc_hd__nor2_4 _1546_ (.A(net19),
    .B(_0885_),
    .Y(_0903_));
 sky130_fd_sc_hd__mux2_1 _1547_ (.A0(\RAM[40][0] ),
    .A1(net56),
    .S(_0903_),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _1548_ (.A0(\RAM[40][1] ),
    .A1(net37),
    .S(_0903_),
    .X(_0161_));
 sky130_fd_sc_hd__mux2_1 _1549_ (.A0(\RAM[40][2] ),
    .A1(net113),
    .S(_0903_),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _1550_ (.A0(\RAM[40][3] ),
    .A1(net96),
    .S(_0903_),
    .X(_0163_));
 sky130_fd_sc_hd__nor2_4 _1551_ (.A(_0833_),
    .B(net19),
    .Y(_0904_));
 sky130_fd_sc_hd__mux2_1 _1552_ (.A0(\RAM[41][0] ),
    .A1(net56),
    .S(_0904_),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_1 _1553_ (.A0(\RAM[41][1] ),
    .A1(net37),
    .S(_0904_),
    .X(_0165_));
 sky130_fd_sc_hd__mux2_1 _1554_ (.A0(\RAM[41][2] ),
    .A1(net113),
    .S(_0904_),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_1 _1555_ (.A0(\RAM[41][3] ),
    .A1(net96),
    .S(_0904_),
    .X(_0167_));
 sky130_fd_sc_hd__nor2_4 _1556_ (.A(net19),
    .B(_0888_),
    .Y(_0905_));
 sky130_fd_sc_hd__mux2_1 _1557_ (.A0(\RAM[42][0] ),
    .A1(net56),
    .S(_0905_),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _1558_ (.A0(\RAM[42][1] ),
    .A1(net37),
    .S(_0905_),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_1 _1559_ (.A0(\RAM[42][2] ),
    .A1(net113),
    .S(_0905_),
    .X(_0170_));
 sky130_fd_sc_hd__mux2_1 _1560_ (.A0(\RAM[42][3] ),
    .A1(net96),
    .S(_0905_),
    .X(_0171_));
 sky130_fd_sc_hd__nand2_4 _1561_ (.A(_0837_),
    .B(_0845_),
    .Y(_0906_));
 sky130_fd_sc_hd__mux2_1 _1562_ (.A0(net56),
    .A1(\RAM[43][0] ),
    .S(_0906_),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_1 _1563_ (.A0(net37),
    .A1(\RAM[43][1] ),
    .S(_0906_),
    .X(_0173_));
 sky130_fd_sc_hd__mux2_1 _1564_ (.A0(net113),
    .A1(\RAM[43][2] ),
    .S(_0906_),
    .X(_0174_));
 sky130_fd_sc_hd__mux2_1 _1565_ (.A0(net96),
    .A1(\RAM[43][3] ),
    .S(_0906_),
    .X(_0175_));
 sky130_fd_sc_hd__nor2_4 _1566_ (.A(net19),
    .B(_0865_),
    .Y(_0907_));
 sky130_fd_sc_hd__mux2_1 _1567_ (.A0(\RAM[44][0] ),
    .A1(net53),
    .S(_0907_),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _1568_ (.A0(\RAM[44][1] ),
    .A1(net36),
    .S(_0907_),
    .X(_0177_));
 sky130_fd_sc_hd__mux2_1 _1569_ (.A0(\RAM[44][2] ),
    .A1(net111),
    .S(_0907_),
    .X(_0178_));
 sky130_fd_sc_hd__mux2_1 _1570_ (.A0(\RAM[44][3] ),
    .A1(net95),
    .S(_0907_),
    .X(_0179_));
 sky130_fd_sc_hd__nand2_4 _1571_ (.A(_0845_),
    .B(_0855_),
    .Y(_0908_));
 sky130_fd_sc_hd__mux2_1 _1572_ (.A0(net53),
    .A1(\RAM[45][0] ),
    .S(_0908_),
    .X(_0180_));
 sky130_fd_sc_hd__mux2_1 _1573_ (.A0(net36),
    .A1(\RAM[45][1] ),
    .S(_0908_),
    .X(_0181_));
 sky130_fd_sc_hd__mux2_1 _1574_ (.A0(net111),
    .A1(\RAM[45][2] ),
    .S(_0908_),
    .X(_0182_));
 sky130_fd_sc_hd__mux2_1 _1575_ (.A0(net95),
    .A1(\RAM[45][3] ),
    .S(_0908_),
    .X(_0183_));
 sky130_fd_sc_hd__nand2_4 _1576_ (.A(_0845_),
    .B(_0870_),
    .Y(_0909_));
 sky130_fd_sc_hd__mux2_1 _1577_ (.A0(net53),
    .A1(\RAM[46][0] ),
    .S(_0909_),
    .X(_0184_));
 sky130_fd_sc_hd__mux2_1 _1578_ (.A0(net36),
    .A1(\RAM[46][1] ),
    .S(_0909_),
    .X(_0185_));
 sky130_fd_sc_hd__mux2_1 _1579_ (.A0(net111),
    .A1(\RAM[46][2] ),
    .S(_0909_),
    .X(_0186_));
 sky130_fd_sc_hd__mux2_1 _1580_ (.A0(net95),
    .A1(\RAM[46][3] ),
    .S(_0909_),
    .X(_0187_));
 sky130_fd_sc_hd__nand2_4 _1581_ (.A(_0845_),
    .B(_0853_),
    .Y(_0910_));
 sky130_fd_sc_hd__mux2_1 _1582_ (.A0(net53),
    .A1(\RAM[47][0] ),
    .S(_0910_),
    .X(_0188_));
 sky130_fd_sc_hd__mux2_1 _1583_ (.A0(net36),
    .A1(\RAM[47][1] ),
    .S(_0910_),
    .X(_0189_));
 sky130_fd_sc_hd__mux2_1 _1584_ (.A0(net112),
    .A1(\RAM[47][2] ),
    .S(_0910_),
    .X(_0190_));
 sky130_fd_sc_hd__mux2_1 _1585_ (.A0(net95),
    .A1(\RAM[47][3] ),
    .S(_0910_),
    .X(_0191_));
 sky130_fd_sc_hd__nor2_2 _1586_ (.A(_0840_),
    .B(_0873_),
    .Y(_0911_));
 sky130_fd_sc_hd__mux2_1 _1587_ (.A0(\RAM[48][0] ),
    .A1(net54),
    .S(_0911_),
    .X(_0192_));
 sky130_fd_sc_hd__mux2_1 _1588_ (.A0(\RAM[48][1] ),
    .A1(net38),
    .S(_0911_),
    .X(_0193_));
 sky130_fd_sc_hd__mux2_1 _1589_ (.A0(\RAM[48][2] ),
    .A1(net115),
    .S(_0911_),
    .X(_0194_));
 sky130_fd_sc_hd__mux2_1 _1590_ (.A0(\RAM[48][3] ),
    .A1(net101),
    .S(_0911_),
    .X(_0195_));
 sky130_fd_sc_hd__nor2_2 _1591_ (.A(net17),
    .B(_0879_),
    .Y(_0912_));
 sky130_fd_sc_hd__mux2_1 _1592_ (.A0(\RAM[4][0] ),
    .A1(net67),
    .S(_0912_),
    .X(_0196_));
 sky130_fd_sc_hd__mux2_1 _1593_ (.A0(\RAM[4][1] ),
    .A1(net51),
    .S(_0912_),
    .X(_0197_));
 sky130_fd_sc_hd__mux2_1 _1594_ (.A0(\RAM[4][2] ),
    .A1(net125),
    .S(_0912_),
    .X(_0198_));
 sky130_fd_sc_hd__mux2_1 _1595_ (.A0(\RAM[4][3] ),
    .A1(net107),
    .S(_0912_),
    .X(_0199_));
 sky130_fd_sc_hd__nor2_4 _1596_ (.A(_0840_),
    .B(_0876_),
    .Y(_0913_));
 sky130_fd_sc_hd__mux2_1 _1597_ (.A0(\RAM[50][0] ),
    .A1(net54),
    .S(_0913_),
    .X(_0200_));
 sky130_fd_sc_hd__mux2_1 _1598_ (.A0(\RAM[50][1] ),
    .A1(net38),
    .S(_0913_),
    .X(_0201_));
 sky130_fd_sc_hd__mux2_1 _1599_ (.A0(\RAM[50][2] ),
    .A1(net115),
    .S(_0913_),
    .X(_0202_));
 sky130_fd_sc_hd__mux2_1 _1600_ (.A0(\RAM[50][3] ),
    .A1(net101),
    .S(_0913_),
    .X(_0203_));
 sky130_fd_sc_hd__nand2_2 _1601_ (.A(_0839_),
    .B(_0848_),
    .Y(_0914_));
 sky130_fd_sc_hd__mux2_1 _1602_ (.A0(net54),
    .A1(\RAM[51][0] ),
    .S(_0914_),
    .X(_0204_));
 sky130_fd_sc_hd__mux2_1 _1603_ (.A0(net38),
    .A1(\RAM[51][1] ),
    .S(_0914_),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _1604_ (.A0(net115),
    .A1(\RAM[51][2] ),
    .S(_0914_),
    .X(_0206_));
 sky130_fd_sc_hd__mux2_1 _1605_ (.A0(net101),
    .A1(\RAM[51][3] ),
    .S(_0914_),
    .X(_0207_));
 sky130_fd_sc_hd__nor2_2 _1606_ (.A(_0840_),
    .B(_0879_),
    .Y(_0915_));
 sky130_fd_sc_hd__mux2_1 _1607_ (.A0(\RAM[52][0] ),
    .A1(net55),
    .S(_0915_),
    .X(_0208_));
 sky130_fd_sc_hd__mux2_1 _1608_ (.A0(\RAM[52][1] ),
    .A1(net45),
    .S(_0915_),
    .X(_0209_));
 sky130_fd_sc_hd__mux2_1 _1609_ (.A0(\RAM[52][2] ),
    .A1(net117),
    .S(_0915_),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_1 _1610_ (.A0(\RAM[52][3] ),
    .A1(net101),
    .S(_0915_),
    .X(_0211_));
 sky130_fd_sc_hd__nand2_2 _1611_ (.A(_0826_),
    .B(_0839_),
    .Y(_0916_));
 sky130_fd_sc_hd__mux2_1 _1612_ (.A0(net55),
    .A1(\RAM[53][0] ),
    .S(_0916_),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_1 _1613_ (.A0(net45),
    .A1(\RAM[53][1] ),
    .S(_0916_),
    .X(_0213_));
 sky130_fd_sc_hd__mux2_1 _1614_ (.A0(net117),
    .A1(\RAM[53][2] ),
    .S(_0916_),
    .X(_0214_));
 sky130_fd_sc_hd__mux2_1 _1615_ (.A0(net102),
    .A1(\RAM[53][3] ),
    .S(_0916_),
    .X(_0215_));
 sky130_fd_sc_hd__or2_4 _1616_ (.A(_0840_),
    .B(_0882_),
    .X(_0917_));
 sky130_fd_sc_hd__mux2_1 _1617_ (.A0(net55),
    .A1(\RAM[54][0] ),
    .S(_0917_),
    .X(_0216_));
 sky130_fd_sc_hd__mux2_1 _1618_ (.A0(net45),
    .A1(\RAM[54][1] ),
    .S(_0917_),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _1619_ (.A0(net115),
    .A1(\RAM[54][2] ),
    .S(_0917_),
    .X(_0218_));
 sky130_fd_sc_hd__mux2_1 _1620_ (.A0(net101),
    .A1(\RAM[54][3] ),
    .S(_0917_),
    .X(_0219_));
 sky130_fd_sc_hd__nand2_2 _1621_ (.A(_0839_),
    .B(_0844_),
    .Y(_0918_));
 sky130_fd_sc_hd__mux2_1 _1622_ (.A0(net55),
    .A1(\RAM[55][0] ),
    .S(_0918_),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _1623_ (.A0(net48),
    .A1(\RAM[55][1] ),
    .S(_0918_),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _1624_ (.A0(net117),
    .A1(\RAM[55][2] ),
    .S(_0918_),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _1625_ (.A0(net102),
    .A1(\RAM[55][3] ),
    .S(_0918_),
    .X(_0223_));
 sky130_fd_sc_hd__nor2_4 _1626_ (.A(_0840_),
    .B(_0885_),
    .Y(_0919_));
 sky130_fd_sc_hd__mux2_1 _1627_ (.A0(\RAM[56][0] ),
    .A1(net55),
    .S(_0919_),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_1 _1628_ (.A0(\RAM[56][1] ),
    .A1(net38),
    .S(_0919_),
    .X(_0225_));
 sky130_fd_sc_hd__mux2_1 _1629_ (.A0(\RAM[56][2] ),
    .A1(net114),
    .S(_0919_),
    .X(_0226_));
 sky130_fd_sc_hd__mux2_1 _1630_ (.A0(\RAM[56][3] ),
    .A1(net97),
    .S(_0919_),
    .X(_0227_));
 sky130_fd_sc_hd__nand2_2 _1631_ (.A(_0832_),
    .B(_0839_),
    .Y(_0920_));
 sky130_fd_sc_hd__mux2_1 _1632_ (.A0(net55),
    .A1(\RAM[57][0] ),
    .S(_0920_),
    .X(_0228_));
 sky130_fd_sc_hd__mux2_1 _1633_ (.A0(net39),
    .A1(\RAM[57][1] ),
    .S(_0920_),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_1 _1634_ (.A0(net114),
    .A1(\RAM[57][2] ),
    .S(_0920_),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_1 _1635_ (.A0(net97),
    .A1(\RAM[57][3] ),
    .S(_0920_),
    .X(_0231_));
 sky130_fd_sc_hd__or2_4 _1636_ (.A(_0840_),
    .B(_0888_),
    .X(_0921_));
 sky130_fd_sc_hd__mux2_1 _1637_ (.A0(net55),
    .A1(\RAM[58][0] ),
    .S(_0921_),
    .X(_0232_));
 sky130_fd_sc_hd__mux2_1 _1638_ (.A0(net39),
    .A1(\RAM[58][1] ),
    .S(_0921_),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_1 _1639_ (.A0(net112),
    .A1(\RAM[58][2] ),
    .S(_0921_),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _1640_ (.A0(net97),
    .A1(\RAM[58][3] ),
    .S(_0921_),
    .X(_0235_));
 sky130_fd_sc_hd__nor2_2 _1641_ (.A(_0827_),
    .B(net17),
    .Y(_0922_));
 sky130_fd_sc_hd__mux2_1 _1642_ (.A0(\RAM[5][0] ),
    .A1(net67),
    .S(_0922_),
    .X(_0236_));
 sky130_fd_sc_hd__mux2_1 _1643_ (.A0(\RAM[5][1] ),
    .A1(net51),
    .S(_0922_),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _1644_ (.A0(\RAM[5][2] ),
    .A1(net125),
    .S(_0922_),
    .X(_0238_));
 sky130_fd_sc_hd__mux2_1 _1645_ (.A0(\RAM[5][3] ),
    .A1(net107),
    .S(_0922_),
    .X(_0239_));
 sky130_fd_sc_hd__or2_4 _1646_ (.A(_0840_),
    .B(_0865_),
    .X(_0923_));
 sky130_fd_sc_hd__mux2_1 _1647_ (.A0(net54),
    .A1(\RAM[60][0] ),
    .S(_0923_),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _1648_ (.A0(net38),
    .A1(\RAM[60][1] ),
    .S(_0923_),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_1 _1649_ (.A0(net112),
    .A1(\RAM[60][2] ),
    .S(_0923_),
    .X(_0242_));
 sky130_fd_sc_hd__mux2_1 _1650_ (.A0(net97),
    .A1(\RAM[60][3] ),
    .S(_0923_),
    .X(_0243_));
 sky130_fd_sc_hd__nand2_2 _1651_ (.A(_0839_),
    .B(_0855_),
    .Y(_0924_));
 sky130_fd_sc_hd__mux2_1 _1652_ (.A0(net54),
    .A1(\RAM[61][0] ),
    .S(_0924_),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _1653_ (.A0(net38),
    .A1(\RAM[61][1] ),
    .S(_0924_),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _1654_ (.A0(net112),
    .A1(\RAM[61][2] ),
    .S(_0924_),
    .X(_0246_));
 sky130_fd_sc_hd__mux2_1 _1655_ (.A0(net97),
    .A1(\RAM[61][3] ),
    .S(_0924_),
    .X(_0247_));
 sky130_fd_sc_hd__nand2_2 _1656_ (.A(_0839_),
    .B(_0870_),
    .Y(_0925_));
 sky130_fd_sc_hd__mux2_1 _1657_ (.A0(net54),
    .A1(\RAM[62][0] ),
    .S(_0925_),
    .X(_0248_));
 sky130_fd_sc_hd__mux2_1 _1658_ (.A0(net38),
    .A1(\RAM[62][1] ),
    .S(_0925_),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _1659_ (.A0(net112),
    .A1(\RAM[62][2] ),
    .S(_0925_),
    .X(_0250_));
 sky130_fd_sc_hd__mux2_1 _1660_ (.A0(net97),
    .A1(\RAM[62][3] ),
    .S(_0925_),
    .X(_0251_));
 sky130_fd_sc_hd__nand2_4 _1661_ (.A(_0839_),
    .B(_0853_),
    .Y(_0926_));
 sky130_fd_sc_hd__mux2_1 _1662_ (.A0(net54),
    .A1(\RAM[63][0] ),
    .S(_0926_),
    .X(_0252_));
 sky130_fd_sc_hd__mux2_1 _1663_ (.A0(net38),
    .A1(\RAM[63][1] ),
    .S(_0926_),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _1664_ (.A0(net112),
    .A1(\RAM[63][2] ),
    .S(_0926_),
    .X(_0254_));
 sky130_fd_sc_hd__mux2_1 _1665_ (.A0(net110),
    .A1(\RAM[63][3] ),
    .S(_0926_),
    .X(_0255_));
 sky130_fd_sc_hd__nor2_4 _1666_ (.A(_0830_),
    .B(_0873_),
    .Y(_0927_));
 sky130_fd_sc_hd__mux2_1 _1667_ (.A0(\RAM[64][0] ),
    .A1(net64),
    .S(_0927_),
    .X(_0256_));
 sky130_fd_sc_hd__mux2_1 _1668_ (.A0(\RAM[64][1] ),
    .A1(net50),
    .S(_0927_),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _1669_ (.A0(\RAM[64][2] ),
    .A1(net123),
    .S(_0927_),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_1 _1670_ (.A0(\RAM[64][3] ),
    .A1(net105),
    .S(_0927_),
    .X(_0259_));
 sky130_fd_sc_hd__nor2_4 _1671_ (.A(net20),
    .B(_0842_),
    .Y(_0928_));
 sky130_fd_sc_hd__mux2_1 _1672_ (.A0(\RAM[65][0] ),
    .A1(net64),
    .S(_0928_),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_1 _1673_ (.A0(\RAM[65][1] ),
    .A1(net50),
    .S(_0928_),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _1674_ (.A0(\RAM[65][2] ),
    .A1(net123),
    .S(_0928_),
    .X(_0262_));
 sky130_fd_sc_hd__mux2_1 _1675_ (.A0(\RAM[65][3] ),
    .A1(net105),
    .S(_0928_),
    .X(_0263_));
 sky130_fd_sc_hd__nor2_4 _1676_ (.A(net20),
    .B(_0876_),
    .Y(_0929_));
 sky130_fd_sc_hd__mux2_1 _1677_ (.A0(\RAM[66][0] ),
    .A1(net64),
    .S(_0929_),
    .X(_0264_));
 sky130_fd_sc_hd__mux2_1 _1678_ (.A0(\RAM[66][1] ),
    .A1(net49),
    .S(_0929_),
    .X(_0265_));
 sky130_fd_sc_hd__mux2_1 _1679_ (.A0(\RAM[66][2] ),
    .A1(net123),
    .S(_0929_),
    .X(_0266_));
 sky130_fd_sc_hd__mux2_1 _1680_ (.A0(\RAM[66][3] ),
    .A1(net105),
    .S(_0929_),
    .X(_0267_));
 sky130_fd_sc_hd__nor2_4 _1681_ (.A(net20),
    .B(_0849_),
    .Y(_0930_));
 sky130_fd_sc_hd__mux2_1 _1682_ (.A0(\RAM[67][0] ),
    .A1(net64),
    .S(_0930_),
    .X(_0268_));
 sky130_fd_sc_hd__mux2_1 _1683_ (.A0(\RAM[67][1] ),
    .A1(net49),
    .S(_0930_),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _1684_ (.A0(\RAM[67][2] ),
    .A1(net123),
    .S(_0930_),
    .X(_0270_));
 sky130_fd_sc_hd__mux2_1 _1685_ (.A0(\RAM[67][3] ),
    .A1(net105),
    .S(_0930_),
    .X(_0271_));
 sky130_fd_sc_hd__nor2_2 _1686_ (.A(net20),
    .B(_0879_),
    .Y(_0931_));
 sky130_fd_sc_hd__mux2_1 _1687_ (.A0(\RAM[68][0] ),
    .A1(net66),
    .S(_0931_),
    .X(_0272_));
 sky130_fd_sc_hd__mux2_1 _1688_ (.A0(\RAM[68][1] ),
    .A1(net50),
    .S(_0931_),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _1689_ (.A0(\RAM[68][2] ),
    .A1(net125),
    .S(_0931_),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_1 _1690_ (.A0(\RAM[68][3] ),
    .A1(net105),
    .S(_0931_),
    .X(_0275_));
 sky130_fd_sc_hd__nor2_2 _1691_ (.A(_0867_),
    .B(_0882_),
    .Y(_0932_));
 sky130_fd_sc_hd__mux2_1 _1692_ (.A0(\RAM[6][0] ),
    .A1(net67),
    .S(_0932_),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_1 _1693_ (.A0(\RAM[6][1] ),
    .A1(net51),
    .S(_0932_),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_1 _1694_ (.A0(\RAM[6][2] ),
    .A1(net124),
    .S(_0932_),
    .X(_0278_));
 sky130_fd_sc_hd__mux2_1 _1695_ (.A0(\RAM[6][3] ),
    .A1(net107),
    .S(_0932_),
    .X(_0279_));
 sky130_fd_sc_hd__nor2_4 _1696_ (.A(net20),
    .B(_0882_),
    .Y(_0933_));
 sky130_fd_sc_hd__mux2_1 _1697_ (.A0(\RAM[70][0] ),
    .A1(net66),
    .S(_0933_),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_1 _1698_ (.A0(\RAM[70][1] ),
    .A1(net50),
    .S(_0933_),
    .X(_0281_));
 sky130_fd_sc_hd__mux2_1 _1699_ (.A0(\RAM[70][2] ),
    .A1(net125),
    .S(_0933_),
    .X(_0282_));
 sky130_fd_sc_hd__mux2_1 _1700_ (.A0(\RAM[70][3] ),
    .A1(net108),
    .S(_0933_),
    .X(_0283_));
 sky130_fd_sc_hd__nand2_4 _1701_ (.A(_0829_),
    .B(_0844_),
    .Y(_0934_));
 sky130_fd_sc_hd__mux2_1 _1702_ (.A0(net66),
    .A1(\RAM[71][0] ),
    .S(_0934_),
    .X(_0284_));
 sky130_fd_sc_hd__mux2_1 _1703_ (.A0(net50),
    .A1(\RAM[71][1] ),
    .S(_0934_),
    .X(_0285_));
 sky130_fd_sc_hd__mux2_1 _1704_ (.A0(net125),
    .A1(\RAM[71][2] ),
    .S(_0934_),
    .X(_0286_));
 sky130_fd_sc_hd__mux2_1 _1705_ (.A0(net108),
    .A1(\RAM[71][3] ),
    .S(_0934_),
    .X(_0287_));
 sky130_fd_sc_hd__nor2_2 _1706_ (.A(net20),
    .B(_0885_),
    .Y(_0935_));
 sky130_fd_sc_hd__mux2_1 _1707_ (.A0(\RAM[72][0] ),
    .A1(net63),
    .S(_0935_),
    .X(_0288_));
 sky130_fd_sc_hd__mux2_1 _1708_ (.A0(\RAM[72][1] ),
    .A1(net42),
    .S(_0935_),
    .X(_0289_));
 sky130_fd_sc_hd__mux2_1 _1709_ (.A0(\RAM[72][2] ),
    .A1(net121),
    .S(_0935_),
    .X(_0290_));
 sky130_fd_sc_hd__mux2_1 _1710_ (.A0(\RAM[72][3] ),
    .A1(net100),
    .S(_0935_),
    .X(_0291_));
 sky130_fd_sc_hd__nor2_4 _1711_ (.A(net20),
    .B(_0833_),
    .Y(_0936_));
 sky130_fd_sc_hd__mux2_1 _1712_ (.A0(\RAM[73][0] ),
    .A1(net63),
    .S(_0936_),
    .X(_0292_));
 sky130_fd_sc_hd__mux2_1 _1713_ (.A0(\RAM[73][1] ),
    .A1(net42),
    .S(_0936_),
    .X(_0293_));
 sky130_fd_sc_hd__mux2_1 _1714_ (.A0(\RAM[73][2] ),
    .A1(net121),
    .S(_0936_),
    .X(_0294_));
 sky130_fd_sc_hd__mux2_1 _1715_ (.A0(\RAM[73][3] ),
    .A1(net100),
    .S(_0936_),
    .X(_0295_));
 sky130_fd_sc_hd__nor2_2 _1716_ (.A(net20),
    .B(_0888_),
    .Y(_0937_));
 sky130_fd_sc_hd__mux2_1 _1717_ (.A0(\RAM[74][0] ),
    .A1(net63),
    .S(_0937_),
    .X(_0296_));
 sky130_fd_sc_hd__mux2_1 _1718_ (.A0(\RAM[74][1] ),
    .A1(net43),
    .S(_0937_),
    .X(_0297_));
 sky130_fd_sc_hd__mux2_1 _1719_ (.A0(\RAM[74][2] ),
    .A1(net121),
    .S(_0937_),
    .X(_0298_));
 sky130_fd_sc_hd__mux2_1 _1720_ (.A0(\RAM[74][3] ),
    .A1(net100),
    .S(_0937_),
    .X(_0299_));
 sky130_fd_sc_hd__nand2_4 _1721_ (.A(_0829_),
    .B(_0837_),
    .Y(_0938_));
 sky130_fd_sc_hd__mux2_1 _1722_ (.A0(net63),
    .A1(\RAM[75][0] ),
    .S(_0938_),
    .X(_0300_));
 sky130_fd_sc_hd__mux2_1 _1723_ (.A0(net43),
    .A1(\RAM[75][1] ),
    .S(_0938_),
    .X(_0301_));
 sky130_fd_sc_hd__mux2_1 _1724_ (.A0(net121),
    .A1(\RAM[75][2] ),
    .S(_0938_),
    .X(_0302_));
 sky130_fd_sc_hd__mux2_1 _1725_ (.A0(net100),
    .A1(\RAM[75][3] ),
    .S(_0938_),
    .X(_0303_));
 sky130_fd_sc_hd__nor2_2 _1726_ (.A(net20),
    .B(_0865_),
    .Y(_0939_));
 sky130_fd_sc_hd__mux2_1 _1727_ (.A0(\RAM[76][0] ),
    .A1(net63),
    .S(_0939_),
    .X(_0304_));
 sky130_fd_sc_hd__mux2_1 _1728_ (.A0(\RAM[76][1] ),
    .A1(net43),
    .S(_0939_),
    .X(_0305_));
 sky130_fd_sc_hd__mux2_1 _1729_ (.A0(\RAM[76][2] ),
    .A1(net125),
    .S(_0939_),
    .X(_0306_));
 sky130_fd_sc_hd__mux2_1 _1730_ (.A0(\RAM[76][3] ),
    .A1(net108),
    .S(_0939_),
    .X(_0307_));
 sky130_fd_sc_hd__nand2_2 _1731_ (.A(_0829_),
    .B(_0855_),
    .Y(_0940_));
 sky130_fd_sc_hd__mux2_1 _1732_ (.A0(net63),
    .A1(\RAM[77][0] ),
    .S(_0940_),
    .X(_0308_));
 sky130_fd_sc_hd__mux2_1 _1733_ (.A0(net43),
    .A1(\RAM[77][1] ),
    .S(_0940_),
    .X(_0309_));
 sky130_fd_sc_hd__mux2_1 _1734_ (.A0(net121),
    .A1(\RAM[77][2] ),
    .S(_0940_),
    .X(_0310_));
 sky130_fd_sc_hd__mux2_1 _1735_ (.A0(net100),
    .A1(\RAM[77][3] ),
    .S(_0940_),
    .X(_0311_));
 sky130_fd_sc_hd__nand2_2 _1736_ (.A(_0829_),
    .B(_0870_),
    .Y(_0941_));
 sky130_fd_sc_hd__mux2_1 _1737_ (.A0(net66),
    .A1(\RAM[78][0] ),
    .S(_0941_),
    .X(_0312_));
 sky130_fd_sc_hd__mux2_1 _1738_ (.A0(net43),
    .A1(\RAM[78][1] ),
    .S(_0941_),
    .X(_0313_));
 sky130_fd_sc_hd__mux2_1 _1739_ (.A0(net125),
    .A1(\RAM[78][2] ),
    .S(_0941_),
    .X(_0314_));
 sky130_fd_sc_hd__mux2_1 _1740_ (.A0(net108),
    .A1(\RAM[78][3] ),
    .S(_0941_),
    .X(_0315_));
 sky130_fd_sc_hd__nand2_4 _1741_ (.A(_0844_),
    .B(_0866_),
    .Y(_0942_));
 sky130_fd_sc_hd__mux2_1 _1742_ (.A0(net67),
    .A1(\RAM[7][0] ),
    .S(_0942_),
    .X(_0316_));
 sky130_fd_sc_hd__mux2_1 _1743_ (.A0(net52),
    .A1(\RAM[7][1] ),
    .S(_0942_),
    .X(_0317_));
 sky130_fd_sc_hd__mux2_1 _1744_ (.A0(net124),
    .A1(\RAM[7][2] ),
    .S(_0942_),
    .X(_0318_));
 sky130_fd_sc_hd__mux2_1 _1745_ (.A0(net107),
    .A1(\RAM[7][3] ),
    .S(_0942_),
    .X(_0319_));
 sky130_fd_sc_hd__nor2_2 _1746_ (.A(_0835_),
    .B(_0873_),
    .Y(_0943_));
 sky130_fd_sc_hd__mux2_1 _1747_ (.A0(\RAM[80][0] ),
    .A1(net57),
    .S(_0943_),
    .X(_0320_));
 sky130_fd_sc_hd__mux2_1 _1748_ (.A0(\RAM[80][1] ),
    .A1(net45),
    .S(_0943_),
    .X(_0321_));
 sky130_fd_sc_hd__mux2_1 _1749_ (.A0(\RAM[80][2] ),
    .A1(net115),
    .S(_0943_),
    .X(_0322_));
 sky130_fd_sc_hd__mux2_1 _1750_ (.A0(\RAM[80][3] ),
    .A1(net101),
    .S(_0943_),
    .X(_0323_));
 sky130_fd_sc_hd__nor2_4 _1751_ (.A(_0835_),
    .B(_0842_),
    .Y(_0944_));
 sky130_fd_sc_hd__mux2_1 _1752_ (.A0(\RAM[81][0] ),
    .A1(net57),
    .S(_0944_),
    .X(_0324_));
 sky130_fd_sc_hd__mux2_1 _1753_ (.A0(\RAM[81][1] ),
    .A1(net45),
    .S(_0944_),
    .X(_0325_));
 sky130_fd_sc_hd__mux2_1 _1754_ (.A0(\RAM[81][2] ),
    .A1(net115),
    .S(_0944_),
    .X(_0326_));
 sky130_fd_sc_hd__mux2_1 _1755_ (.A0(\RAM[81][3] ),
    .A1(net101),
    .S(_0944_),
    .X(_0327_));
 sky130_fd_sc_hd__nor2_4 _1756_ (.A(_0835_),
    .B(_0876_),
    .Y(_0945_));
 sky130_fd_sc_hd__mux2_1 _1757_ (.A0(\RAM[82][0] ),
    .A1(net57),
    .S(_0945_),
    .X(_0328_));
 sky130_fd_sc_hd__mux2_1 _1758_ (.A0(\RAM[82][1] ),
    .A1(net45),
    .S(_0945_),
    .X(_0329_));
 sky130_fd_sc_hd__mux2_1 _1759_ (.A0(\RAM[82][2] ),
    .A1(net115),
    .S(_0945_),
    .X(_0330_));
 sky130_fd_sc_hd__mux2_1 _1760_ (.A0(\RAM[82][3] ),
    .A1(net101),
    .S(_0945_),
    .X(_0331_));
 sky130_fd_sc_hd__nand2_4 _1761_ (.A(_0834_),
    .B(_0848_),
    .Y(_0946_));
 sky130_fd_sc_hd__mux2_1 _1762_ (.A0(net57),
    .A1(\RAM[83][0] ),
    .S(_0946_),
    .X(_0332_));
 sky130_fd_sc_hd__mux2_1 _1763_ (.A0(net45),
    .A1(\RAM[83][1] ),
    .S(_0946_),
    .X(_0333_));
 sky130_fd_sc_hd__mux2_1 _1764_ (.A0(net115),
    .A1(\RAM[83][2] ),
    .S(_0946_),
    .X(_0334_));
 sky130_fd_sc_hd__mux2_1 _1765_ (.A0(net101),
    .A1(\RAM[83][3] ),
    .S(_0946_),
    .X(_0335_));
 sky130_fd_sc_hd__nor2_2 _1766_ (.A(_0835_),
    .B(_0879_),
    .Y(_0947_));
 sky130_fd_sc_hd__mux2_1 _1767_ (.A0(\RAM[84][0] ),
    .A1(net65),
    .S(_0947_),
    .X(_0336_));
 sky130_fd_sc_hd__mux2_1 _1768_ (.A0(\RAM[84][1] ),
    .A1(net51),
    .S(_0947_),
    .X(_0337_));
 sky130_fd_sc_hd__mux2_1 _1769_ (.A0(\RAM[84][2] ),
    .A1(net123),
    .S(_0947_),
    .X(_0338_));
 sky130_fd_sc_hd__mux2_1 _1770_ (.A0(\RAM[84][3] ),
    .A1(net106),
    .S(_0947_),
    .X(_0339_));
 sky130_fd_sc_hd__nand2_4 _1771_ (.A(_0826_),
    .B(_0834_),
    .Y(_0948_));
 sky130_fd_sc_hd__mux2_1 _1772_ (.A0(net65),
    .A1(\RAM[85][0] ),
    .S(_0948_),
    .X(_0340_));
 sky130_fd_sc_hd__mux2_1 _1773_ (.A0(net51),
    .A1(\RAM[85][1] ),
    .S(_0948_),
    .X(_0341_));
 sky130_fd_sc_hd__mux2_1 _1774_ (.A0(net126),
    .A1(\RAM[85][2] ),
    .S(_0948_),
    .X(_0342_));
 sky130_fd_sc_hd__mux2_1 _1775_ (.A0(net106),
    .A1(\RAM[85][3] ),
    .S(_0948_),
    .X(_0343_));
 sky130_fd_sc_hd__or2_4 _1776_ (.A(_0835_),
    .B(_0882_),
    .X(_0949_));
 sky130_fd_sc_hd__mux2_1 _1777_ (.A0(net59),
    .A1(\RAM[86][0] ),
    .S(_0949_),
    .X(_0344_));
 sky130_fd_sc_hd__mux2_1 _1778_ (.A0(net47),
    .A1(\RAM[86][1] ),
    .S(_0949_),
    .X(_0345_));
 sky130_fd_sc_hd__mux2_1 _1779_ (.A0(net118),
    .A1(\RAM[86][2] ),
    .S(_0949_),
    .X(_0346_));
 sky130_fd_sc_hd__mux2_1 _1780_ (.A0(net104),
    .A1(\RAM[86][3] ),
    .S(_0949_),
    .X(_0347_));
 sky130_fd_sc_hd__nand2_2 _1781_ (.A(_0834_),
    .B(_0844_),
    .Y(_0950_));
 sky130_fd_sc_hd__mux2_1 _1782_ (.A0(net65),
    .A1(\RAM[87][0] ),
    .S(_0950_),
    .X(_0348_));
 sky130_fd_sc_hd__mux2_1 _1783_ (.A0(net51),
    .A1(\RAM[87][1] ),
    .S(_0950_),
    .X(_0349_));
 sky130_fd_sc_hd__mux2_1 _1784_ (.A0(net118),
    .A1(\RAM[87][2] ),
    .S(_0950_),
    .X(_0350_));
 sky130_fd_sc_hd__mux2_1 _1785_ (.A0(net104),
    .A1(\RAM[87][3] ),
    .S(_0950_),
    .X(_0351_));
 sky130_fd_sc_hd__nor2_2 _1786_ (.A(_0835_),
    .B(_0885_),
    .Y(_0951_));
 sky130_fd_sc_hd__mux2_1 _1787_ (.A0(\RAM[88][0] ),
    .A1(net64),
    .S(_0951_),
    .X(_0352_));
 sky130_fd_sc_hd__mux2_1 _1788_ (.A0(\RAM[88][1] ),
    .A1(net49),
    .S(_0951_),
    .X(_0353_));
 sky130_fd_sc_hd__mux2_1 _1789_ (.A0(\RAM[88][2] ),
    .A1(net123),
    .S(_0951_),
    .X(_0354_));
 sky130_fd_sc_hd__mux2_1 _1790_ (.A0(\RAM[88][3] ),
    .A1(net106),
    .S(_0951_),
    .X(_0355_));
 sky130_fd_sc_hd__nor2_2 _1791_ (.A(net17),
    .B(_0885_),
    .Y(_0952_));
 sky130_fd_sc_hd__mux2_1 _1792_ (.A0(\RAM[8][0] ),
    .A1(net66),
    .S(_0952_),
    .X(_0356_));
 sky130_fd_sc_hd__mux2_1 _1793_ (.A0(\RAM[8][1] ),
    .A1(net50),
    .S(_0952_),
    .X(_0357_));
 sky130_fd_sc_hd__mux2_1 _1794_ (.A0(\RAM[8][2] ),
    .A1(net124),
    .S(_0952_),
    .X(_0358_));
 sky130_fd_sc_hd__mux2_1 _1795_ (.A0(\RAM[8][3] ),
    .A1(net106),
    .S(_0952_),
    .X(_0359_));
 sky130_fd_sc_hd__or2_2 _1796_ (.A(_0835_),
    .B(_0888_),
    .X(_0953_));
 sky130_fd_sc_hd__mux2_1 _1797_ (.A0(net58),
    .A1(\RAM[90][0] ),
    .S(_0953_),
    .X(_0360_));
 sky130_fd_sc_hd__mux2_1 _1798_ (.A0(net48),
    .A1(\RAM[90][1] ),
    .S(_0953_),
    .X(_0361_));
 sky130_fd_sc_hd__mux2_1 _1799_ (.A0(net117),
    .A1(\RAM[90][2] ),
    .S(_0953_),
    .X(_0362_));
 sky130_fd_sc_hd__mux2_1 _1800_ (.A0(net104),
    .A1(\RAM[90][3] ),
    .S(_0953_),
    .X(_0363_));
 sky130_fd_sc_hd__nand2_2 _1801_ (.A(_0834_),
    .B(_0837_),
    .Y(_0954_));
 sky130_fd_sc_hd__mux2_1 _1802_ (.A0(net58),
    .A1(\RAM[91][0] ),
    .S(_0954_),
    .X(_0364_));
 sky130_fd_sc_hd__mux2_1 _1803_ (.A0(net49),
    .A1(\RAM[91][1] ),
    .S(_0954_),
    .X(_0365_));
 sky130_fd_sc_hd__mux2_1 _1804_ (.A0(net123),
    .A1(\RAM[91][2] ),
    .S(_0954_),
    .X(_0366_));
 sky130_fd_sc_hd__mux2_1 _1805_ (.A0(net102),
    .A1(\RAM[91][3] ),
    .S(_0954_),
    .X(_0367_));
 sky130_fd_sc_hd__or2_4 _1806_ (.A(_0835_),
    .B(_0865_),
    .X(_0955_));
 sky130_fd_sc_hd__mux2_1 _1807_ (.A0(net58),
    .A1(\RAM[92][0] ),
    .S(_0955_),
    .X(_0368_));
 sky130_fd_sc_hd__mux2_1 _1808_ (.A0(net48),
    .A1(\RAM[92][1] ),
    .S(_0955_),
    .X(_0369_));
 sky130_fd_sc_hd__mux2_1 _1809_ (.A0(net117),
    .A1(\RAM[92][2] ),
    .S(_0955_),
    .X(_0370_));
 sky130_fd_sc_hd__mux2_1 _1810_ (.A0(net102),
    .A1(\RAM[92][3] ),
    .S(_0955_),
    .X(_0371_));
 sky130_fd_sc_hd__nand2_2 _1811_ (.A(_0834_),
    .B(_0855_),
    .Y(_0956_));
 sky130_fd_sc_hd__mux2_1 _1812_ (.A0(net58),
    .A1(\RAM[93][0] ),
    .S(_0956_),
    .X(_0372_));
 sky130_fd_sc_hd__mux2_1 _1813_ (.A0(net45),
    .A1(\RAM[93][1] ),
    .S(_0956_),
    .X(_0373_));
 sky130_fd_sc_hd__mux2_1 _1814_ (.A0(net115),
    .A1(\RAM[93][2] ),
    .S(_0956_),
    .X(_0374_));
 sky130_fd_sc_hd__mux2_1 _1815_ (.A0(net102),
    .A1(\RAM[93][3] ),
    .S(_0956_),
    .X(_0375_));
 sky130_fd_sc_hd__nand2_2 _1816_ (.A(_0834_),
    .B(_0870_),
    .Y(_0957_));
 sky130_fd_sc_hd__mux2_1 _1817_ (.A0(net58),
    .A1(\RAM[94][0] ),
    .S(_0957_),
    .X(_0376_));
 sky130_fd_sc_hd__mux2_1 _1818_ (.A0(net45),
    .A1(\RAM[94][1] ),
    .S(_0957_),
    .X(_0377_));
 sky130_fd_sc_hd__mux2_1 _1819_ (.A0(net116),
    .A1(\RAM[94][2] ),
    .S(_0957_),
    .X(_0378_));
 sky130_fd_sc_hd__mux2_1 _1820_ (.A0(net102),
    .A1(\RAM[94][3] ),
    .S(_0957_),
    .X(_0379_));
 sky130_fd_sc_hd__nand2_2 _1821_ (.A(_0834_),
    .B(_0853_),
    .Y(_0958_));
 sky130_fd_sc_hd__mux2_1 _1822_ (.A0(net58),
    .A1(\RAM[95][0] ),
    .S(_0958_),
    .X(_0380_));
 sky130_fd_sc_hd__mux2_1 _1823_ (.A0(net45),
    .A1(\RAM[95][1] ),
    .S(_0958_),
    .X(_0381_));
 sky130_fd_sc_hd__mux2_1 _1824_ (.A0(net116),
    .A1(\RAM[95][2] ),
    .S(_0958_),
    .X(_0382_));
 sky130_fd_sc_hd__mux2_1 _1825_ (.A0(net102),
    .A1(\RAM[95][3] ),
    .S(_0958_),
    .X(_0383_));
 sky130_fd_sc_hd__nor2_2 _1826_ (.A(_0858_),
    .B(_0873_),
    .Y(_0959_));
 sky130_fd_sc_hd__mux2_1 _1827_ (.A0(\RAM[96][0] ),
    .A1(net60),
    .S(_0959_),
    .X(_0384_));
 sky130_fd_sc_hd__mux2_1 _1828_ (.A0(\RAM[96][1] ),
    .A1(net40),
    .S(_0959_),
    .X(_0385_));
 sky130_fd_sc_hd__mux2_1 _1829_ (.A0(\RAM[96][2] ),
    .A1(net119),
    .S(_0959_),
    .X(_0386_));
 sky130_fd_sc_hd__mux2_1 _1830_ (.A0(\RAM[96][3] ),
    .A1(net98),
    .S(_0959_),
    .X(_0387_));
 sky130_fd_sc_hd__nor2_4 _1831_ (.A(_0842_),
    .B(_0858_),
    .Y(_0960_));
 sky130_fd_sc_hd__mux2_1 _1832_ (.A0(\RAM[97][0] ),
    .A1(net60),
    .S(_0960_),
    .X(_0388_));
 sky130_fd_sc_hd__mux2_1 _1833_ (.A0(\RAM[97][1] ),
    .A1(net40),
    .S(_0960_),
    .X(_0389_));
 sky130_fd_sc_hd__mux2_1 _1834_ (.A0(\RAM[97][2] ),
    .A1(net119),
    .S(_0960_),
    .X(_0390_));
 sky130_fd_sc_hd__mux2_1 _1835_ (.A0(\RAM[97][3] ),
    .A1(net98),
    .S(_0960_),
    .X(_0391_));
 sky130_fd_sc_hd__nor2_2 _1836_ (.A(_0858_),
    .B(_0876_),
    .Y(_0961_));
 sky130_fd_sc_hd__mux2_1 _1837_ (.A0(\RAM[98][0] ),
    .A1(net60),
    .S(_0961_),
    .X(_0392_));
 sky130_fd_sc_hd__mux2_1 _1838_ (.A0(\RAM[98][1] ),
    .A1(net40),
    .S(_0961_),
    .X(_0393_));
 sky130_fd_sc_hd__mux2_1 _1839_ (.A0(\RAM[98][2] ),
    .A1(net119),
    .S(_0961_),
    .X(_0394_));
 sky130_fd_sc_hd__mux2_1 _1840_ (.A0(\RAM[98][3] ),
    .A1(net98),
    .S(_0961_),
    .X(_0395_));
 sky130_fd_sc_hd__nor2_4 _1841_ (.A(net17),
    .B(_0873_),
    .Y(_0962_));
 sky130_fd_sc_hd__mux2_1 _1842_ (.A0(\RAM[0][0] ),
    .A1(net65),
    .S(_0962_),
    .X(_0396_));
 sky130_fd_sc_hd__mux2_1 _1843_ (.A0(\RAM[0][1] ),
    .A1(net52),
    .S(_0962_),
    .X(_0397_));
 sky130_fd_sc_hd__mux2_1 _1844_ (.A0(\RAM[0][2] ),
    .A1(net124),
    .S(_0962_),
    .X(_0398_));
 sky130_fd_sc_hd__mux2_1 _1845_ (.A0(\RAM[0][3] ),
    .A1(net107),
    .S(_0962_),
    .X(_0399_));
 sky130_fd_sc_hd__nor2_2 _1846_ (.A(_0858_),
    .B(_0879_),
    .Y(_0963_));
 sky130_fd_sc_hd__mux2_1 _1847_ (.A0(\RAM[100][0] ),
    .A1(net62),
    .S(_0963_),
    .X(_0400_));
 sky130_fd_sc_hd__mux2_1 _1848_ (.A0(\RAM[100][1] ),
    .A1(net41),
    .S(_0963_),
    .X(_0401_));
 sky130_fd_sc_hd__mux2_1 _1849_ (.A0(\RAM[100][2] ),
    .A1(net121),
    .S(_0963_),
    .X(_0402_));
 sky130_fd_sc_hd__mux2_1 _1850_ (.A0(\RAM[100][3] ),
    .A1(net99),
    .S(_0963_),
    .X(_0403_));
 sky130_fd_sc_hd__nand2_4 _1851_ (.A(_0826_),
    .B(_0857_),
    .Y(_0964_));
 sky130_fd_sc_hd__mux2_1 _1852_ (.A0(net62),
    .A1(\RAM[101][0] ),
    .S(_0964_),
    .X(_0404_));
 sky130_fd_sc_hd__mux2_1 _1853_ (.A0(net41),
    .A1(\RAM[101][1] ),
    .S(_0964_),
    .X(_0405_));
 sky130_fd_sc_hd__mux2_1 _1854_ (.A0(net119),
    .A1(\RAM[101][2] ),
    .S(_0964_),
    .X(_0406_));
 sky130_fd_sc_hd__mux2_1 _1855_ (.A0(net99),
    .A1(\RAM[101][3] ),
    .S(_0964_),
    .X(_0407_));
 sky130_fd_sc_hd__or2_4 _1856_ (.A(_0858_),
    .B(_0882_),
    .X(_0965_));
 sky130_fd_sc_hd__mux2_1 _1857_ (.A0(net60),
    .A1(\RAM[102][0] ),
    .S(_0965_),
    .X(_0408_));
 sky130_fd_sc_hd__mux2_1 _1858_ (.A0(net40),
    .A1(\RAM[102][1] ),
    .S(_0965_),
    .X(_0409_));
 sky130_fd_sc_hd__mux2_1 _1859_ (.A0(net119),
    .A1(\RAM[102][2] ),
    .S(_0965_),
    .X(_0410_));
 sky130_fd_sc_hd__mux2_1 _1860_ (.A0(net98),
    .A1(\RAM[102][3] ),
    .S(_0965_),
    .X(_0411_));
 sky130_fd_sc_hd__nand2_2 _1861_ (.A(_0844_),
    .B(_0857_),
    .Y(_0966_));
 sky130_fd_sc_hd__mux2_1 _1862_ (.A0(net60),
    .A1(\RAM[103][0] ),
    .S(_0966_),
    .X(_0412_));
 sky130_fd_sc_hd__mux2_1 _1863_ (.A0(net40),
    .A1(\RAM[103][1] ),
    .S(_0966_),
    .X(_0413_));
 sky130_fd_sc_hd__mux2_1 _1864_ (.A0(net119),
    .A1(\RAM[103][2] ),
    .S(_0966_),
    .X(_0414_));
 sky130_fd_sc_hd__mux2_1 _1865_ (.A0(net98),
    .A1(\RAM[103][3] ),
    .S(_0966_),
    .X(_0415_));
 sky130_fd_sc_hd__nor2_4 _1866_ (.A(_0858_),
    .B(_0885_),
    .Y(_0967_));
 sky130_fd_sc_hd__mux2_1 _1867_ (.A0(\RAM[104][0] ),
    .A1(net62),
    .S(_0967_),
    .X(_0416_));
 sky130_fd_sc_hd__mux2_1 _1868_ (.A0(\RAM[104][1] ),
    .A1(net41),
    .S(_0967_),
    .X(_0417_));
 sky130_fd_sc_hd__mux2_1 _1869_ (.A0(\RAM[104][2] ),
    .A1(net122),
    .S(_0967_),
    .X(_0418_));
 sky130_fd_sc_hd__mux2_1 _1870_ (.A0(\RAM[104][3] ),
    .A1(net99),
    .S(_0967_),
    .X(_0419_));
 sky130_fd_sc_hd__nand2_4 _1871_ (.A(_0832_),
    .B(_0857_),
    .Y(_0968_));
 sky130_fd_sc_hd__mux2_1 _1872_ (.A0(net62),
    .A1(\RAM[105][0] ),
    .S(_0968_),
    .X(_0420_));
 sky130_fd_sc_hd__mux2_1 _1873_ (.A0(net41),
    .A1(\RAM[105][1] ),
    .S(_0968_),
    .X(_0421_));
 sky130_fd_sc_hd__mux2_1 _1874_ (.A0(net122),
    .A1(\RAM[105][2] ),
    .S(_0968_),
    .X(_0422_));
 sky130_fd_sc_hd__mux2_1 _1875_ (.A0(net99),
    .A1(\RAM[105][3] ),
    .S(_0968_),
    .X(_0423_));
 sky130_fd_sc_hd__or2_4 _1876_ (.A(_0858_),
    .B(_0888_),
    .X(_0969_));
 sky130_fd_sc_hd__mux2_1 _1877_ (.A0(net62),
    .A1(\RAM[106][0] ),
    .S(_0969_),
    .X(_0424_));
 sky130_fd_sc_hd__mux2_1 _1878_ (.A0(net41),
    .A1(\RAM[106][1] ),
    .S(_0969_),
    .X(_0425_));
 sky130_fd_sc_hd__mux2_1 _1879_ (.A0(net122),
    .A1(\RAM[106][2] ),
    .S(_0969_),
    .X(_0426_));
 sky130_fd_sc_hd__mux2_1 _1880_ (.A0(net99),
    .A1(\RAM[106][3] ),
    .S(_0969_),
    .X(_0427_));
 sky130_fd_sc_hd__nand2_2 _1881_ (.A(_0837_),
    .B(_0857_),
    .Y(_0970_));
 sky130_fd_sc_hd__mux2_1 _1882_ (.A0(net62),
    .A1(\RAM[107][0] ),
    .S(_0970_),
    .X(_0428_));
 sky130_fd_sc_hd__mux2_1 _1883_ (.A0(net41),
    .A1(\RAM[107][1] ),
    .S(_0970_),
    .X(_0429_));
 sky130_fd_sc_hd__mux2_1 _1884_ (.A0(net122),
    .A1(\RAM[107][2] ),
    .S(_0970_),
    .X(_0430_));
 sky130_fd_sc_hd__mux2_1 _1885_ (.A0(net99),
    .A1(\RAM[107][3] ),
    .S(_0970_),
    .X(_0431_));
 sky130_fd_sc_hd__or2_4 _1886_ (.A(_0858_),
    .B(_0865_),
    .X(_0971_));
 sky130_fd_sc_hd__mux2_1 _1887_ (.A0(net62),
    .A1(\RAM[108][0] ),
    .S(_0971_),
    .X(_0432_));
 sky130_fd_sc_hd__mux2_1 _1888_ (.A0(net41),
    .A1(\RAM[108][1] ),
    .S(_0971_),
    .X(_0433_));
 sky130_fd_sc_hd__mux2_1 _1889_ (.A0(net121),
    .A1(\RAM[108][2] ),
    .S(_0971_),
    .X(_0434_));
 sky130_fd_sc_hd__mux2_1 _1890_ (.A0(net99),
    .A1(\RAM[108][3] ),
    .S(_0971_),
    .X(_0435_));
 sky130_fd_sc_hd__nor2_2 _1891_ (.A(net17),
    .B(_0888_),
    .Y(_0972_));
 sky130_fd_sc_hd__mux2_1 _1892_ (.A0(\RAM[10][0] ),
    .A1(net64),
    .S(_0972_),
    .X(_0436_));
 sky130_fd_sc_hd__mux2_1 _1893_ (.A0(\RAM[10][1] ),
    .A1(net49),
    .S(_0972_),
    .X(_0437_));
 sky130_fd_sc_hd__mux2_1 _1894_ (.A0(\RAM[10][2] ),
    .A1(net126),
    .S(_0972_),
    .X(_0438_));
 sky130_fd_sc_hd__mux2_1 _1895_ (.A0(\RAM[10][3] ),
    .A1(net106),
    .S(_0972_),
    .X(_0439_));
 sky130_fd_sc_hd__nand2_2 _1896_ (.A(_0857_),
    .B(_0870_),
    .Y(_0973_));
 sky130_fd_sc_hd__mux2_1 _1897_ (.A0(net62),
    .A1(\RAM[110][0] ),
    .S(_0973_),
    .X(_0440_));
 sky130_fd_sc_hd__mux2_1 _1898_ (.A0(net41),
    .A1(\RAM[110][1] ),
    .S(_0973_),
    .X(_0441_));
 sky130_fd_sc_hd__mux2_1 _1899_ (.A0(net121),
    .A1(\RAM[110][2] ),
    .S(_0973_),
    .X(_0442_));
 sky130_fd_sc_hd__mux2_1 _1900_ (.A0(net99),
    .A1(\RAM[110][3] ),
    .S(_0973_),
    .X(_0443_));
 sky130_fd_sc_hd__nand2_2 _1901_ (.A(_0853_),
    .B(_0857_),
    .Y(_0974_));
 sky130_fd_sc_hd__mux2_1 _1902_ (.A0(net62),
    .A1(\RAM[111][0] ),
    .S(_0974_),
    .X(_0444_));
 sky130_fd_sc_hd__mux2_1 _1903_ (.A0(net41),
    .A1(\RAM[111][1] ),
    .S(_0974_),
    .X(_0445_));
 sky130_fd_sc_hd__mux2_1 _1904_ (.A0(net121),
    .A1(\RAM[111][2] ),
    .S(_0974_),
    .X(_0446_));
 sky130_fd_sc_hd__mux2_1 _1905_ (.A0(net99),
    .A1(\RAM[111][3] ),
    .S(_0974_),
    .X(_0447_));
 sky130_fd_sc_hd__nor2_2 _1906_ (.A(_0862_),
    .B(_0873_),
    .Y(_0975_));
 sky130_fd_sc_hd__mux2_1 _1907_ (.A0(\RAM[112][0] ),
    .A1(net60),
    .S(_0975_),
    .X(_0448_));
 sky130_fd_sc_hd__mux2_1 _1908_ (.A0(\RAM[112][1] ),
    .A1(net40),
    .S(_0975_),
    .X(_0449_));
 sky130_fd_sc_hd__mux2_1 _1909_ (.A0(\RAM[112][2] ),
    .A1(net119),
    .S(_0975_),
    .X(_0450_));
 sky130_fd_sc_hd__mux2_1 _1910_ (.A0(\RAM[112][3] ),
    .A1(net98),
    .S(_0975_),
    .X(_0451_));
 sky130_fd_sc_hd__nor2_2 _1911_ (.A(_0842_),
    .B(_0862_),
    .Y(_0976_));
 sky130_fd_sc_hd__mux2_1 _1912_ (.A0(\RAM[113][0] ),
    .A1(net55),
    .S(_0976_),
    .X(_0452_));
 sky130_fd_sc_hd__mux2_1 _1913_ (.A0(\RAM[113][1] ),
    .A1(net37),
    .S(_0976_),
    .X(_0453_));
 sky130_fd_sc_hd__mux2_1 _1914_ (.A0(\RAM[113][2] ),
    .A1(net113),
    .S(_0976_),
    .X(_0454_));
 sky130_fd_sc_hd__mux2_1 _1915_ (.A0(\RAM[113][3] ),
    .A1(net96),
    .S(_0976_),
    .X(_0455_));
 sky130_fd_sc_hd__nor2_2 _1916_ (.A(_0862_),
    .B(_0876_),
    .Y(_0977_));
 sky130_fd_sc_hd__mux2_1 _1917_ (.A0(\RAM[114][0] ),
    .A1(net55),
    .S(_0977_),
    .X(_0456_));
 sky130_fd_sc_hd__mux2_1 _1918_ (.A0(\RAM[114][1] ),
    .A1(net37),
    .S(_0977_),
    .X(_0457_));
 sky130_fd_sc_hd__mux2_1 _1919_ (.A0(\RAM[114][2] ),
    .A1(net113),
    .S(_0977_),
    .X(_0458_));
 sky130_fd_sc_hd__mux2_1 _1920_ (.A0(\RAM[114][3] ),
    .A1(net96),
    .S(_0977_),
    .X(_0459_));
 sky130_fd_sc_hd__nand2_2 _1921_ (.A(_0848_),
    .B(_0861_),
    .Y(_0978_));
 sky130_fd_sc_hd__mux2_1 _1922_ (.A0(net56),
    .A1(\RAM[115][0] ),
    .S(_0978_),
    .X(_0460_));
 sky130_fd_sc_hd__mux2_1 _1923_ (.A0(net39),
    .A1(\RAM[115][1] ),
    .S(_0978_),
    .X(_0461_));
 sky130_fd_sc_hd__mux2_1 _1924_ (.A0(net113),
    .A1(\RAM[115][2] ),
    .S(_0978_),
    .X(_0462_));
 sky130_fd_sc_hd__mux2_1 _1925_ (.A0(net96),
    .A1(\RAM[115][3] ),
    .S(_0978_),
    .X(_0463_));
 sky130_fd_sc_hd__nor2_2 _1926_ (.A(_0862_),
    .B(_0879_),
    .Y(_0979_));
 sky130_fd_sc_hd__mux2_1 _1927_ (.A0(\RAM[116][0] ),
    .A1(net61),
    .S(_0979_),
    .X(_0464_));
 sky130_fd_sc_hd__mux2_1 _1928_ (.A0(\RAM[116][1] ),
    .A1(net42),
    .S(_0979_),
    .X(_0465_));
 sky130_fd_sc_hd__mux2_1 _1929_ (.A0(\RAM[116][2] ),
    .A1(net120),
    .S(_0979_),
    .X(_0466_));
 sky130_fd_sc_hd__mux2_1 _1930_ (.A0(\RAM[116][3] ),
    .A1(net105),
    .S(_0979_),
    .X(_0467_));
 sky130_fd_sc_hd__nand2_2 _1931_ (.A(_0826_),
    .B(_0861_),
    .Y(_0980_));
 sky130_fd_sc_hd__mux2_1 _1932_ (.A0(net61),
    .A1(\RAM[117][0] ),
    .S(_0980_),
    .X(_0468_));
 sky130_fd_sc_hd__mux2_1 _1933_ (.A0(net42),
    .A1(\RAM[117][1] ),
    .S(_0980_),
    .X(_0469_));
 sky130_fd_sc_hd__mux2_1 _1934_ (.A0(net120),
    .A1(\RAM[117][2] ),
    .S(_0980_),
    .X(_0470_));
 sky130_fd_sc_hd__mux2_1 _1935_ (.A0(net105),
    .A1(\RAM[117][3] ),
    .S(_0980_),
    .X(_0471_));
 sky130_fd_sc_hd__or2_4 _1936_ (.A(_0862_),
    .B(_0882_),
    .X(_0981_));
 sky130_fd_sc_hd__mux2_1 _1937_ (.A0(net56),
    .A1(\RAM[118][0] ),
    .S(_0981_),
    .X(_0472_));
 sky130_fd_sc_hd__mux2_1 _1938_ (.A0(net39),
    .A1(\RAM[118][1] ),
    .S(_0981_),
    .X(_0473_));
 sky130_fd_sc_hd__mux2_1 _1939_ (.A0(net114),
    .A1(\RAM[118][2] ),
    .S(_0981_),
    .X(_0474_));
 sky130_fd_sc_hd__mux2_1 _1940_ (.A0(net102),
    .A1(\RAM[118][3] ),
    .S(_0981_),
    .X(_0475_));
 sky130_fd_sc_hd__nand2_2 _1941_ (.A(_0837_),
    .B(_0866_),
    .Y(_0982_));
 sky130_fd_sc_hd__mux2_1 _1942_ (.A0(net64),
    .A1(\RAM[11][0] ),
    .S(_0982_),
    .X(_0476_));
 sky130_fd_sc_hd__mux2_1 _1943_ (.A0(net49),
    .A1(\RAM[11][1] ),
    .S(_0982_),
    .X(_0477_));
 sky130_fd_sc_hd__mux2_1 _1944_ (.A0(net126),
    .A1(\RAM[11][2] ),
    .S(_0982_),
    .X(_0478_));
 sky130_fd_sc_hd__mux2_1 _1945_ (.A0(net106),
    .A1(\RAM[11][3] ),
    .S(_0982_),
    .X(_0479_));
 sky130_fd_sc_hd__nor2_2 _1946_ (.A(_0862_),
    .B(_0885_),
    .Y(_0983_));
 sky130_fd_sc_hd__mux2_1 _1947_ (.A0(\RAM[120][0] ),
    .A1(net61),
    .S(_0983_),
    .X(_0480_));
 sky130_fd_sc_hd__mux2_1 _1948_ (.A0(\RAM[120][1] ),
    .A1(net42),
    .S(_0983_),
    .X(_0481_));
 sky130_fd_sc_hd__mux2_1 _1949_ (.A0(\RAM[120][2] ),
    .A1(net120),
    .S(_0983_),
    .X(_0482_));
 sky130_fd_sc_hd__mux2_1 _1950_ (.A0(\RAM[120][3] ),
    .A1(net100),
    .S(_0983_),
    .X(_0483_));
 sky130_fd_sc_hd__nand2_4 _1951_ (.A(_0832_),
    .B(_0861_),
    .Y(_0984_));
 sky130_fd_sc_hd__mux2_1 _1952_ (.A0(net61),
    .A1(\RAM[121][0] ),
    .S(_0984_),
    .X(_0484_));
 sky130_fd_sc_hd__mux2_1 _1953_ (.A0(net42),
    .A1(\RAM[121][1] ),
    .S(_0984_),
    .X(_0485_));
 sky130_fd_sc_hd__mux2_1 _1954_ (.A0(net120),
    .A1(\RAM[121][2] ),
    .S(_0984_),
    .X(_0486_));
 sky130_fd_sc_hd__mux2_1 _1955_ (.A0(net100),
    .A1(\RAM[121][3] ),
    .S(_0984_),
    .X(_0487_));
 sky130_fd_sc_hd__or2_4 _1956_ (.A(_0862_),
    .B(_0888_),
    .X(_0985_));
 sky130_fd_sc_hd__mux2_1 _1957_ (.A0(net61),
    .A1(\RAM[122][0] ),
    .S(_0985_),
    .X(_0488_));
 sky130_fd_sc_hd__mux2_1 _1958_ (.A0(net42),
    .A1(\RAM[122][1] ),
    .S(_0985_),
    .X(_0489_));
 sky130_fd_sc_hd__mux2_1 _1959_ (.A0(net120),
    .A1(\RAM[122][2] ),
    .S(_0985_),
    .X(_0490_));
 sky130_fd_sc_hd__mux2_1 _1960_ (.A0(net100),
    .A1(\RAM[122][3] ),
    .S(_0985_),
    .X(_0491_));
 sky130_fd_sc_hd__nand2_2 _1961_ (.A(_0837_),
    .B(_0861_),
    .Y(_0986_));
 sky130_fd_sc_hd__mux2_1 _1962_ (.A0(net61),
    .A1(\RAM[123][0] ),
    .S(_0986_),
    .X(_0492_));
 sky130_fd_sc_hd__mux2_1 _1963_ (.A0(net42),
    .A1(\RAM[123][1] ),
    .S(_0986_),
    .X(_0493_));
 sky130_fd_sc_hd__mux2_1 _1964_ (.A0(net120),
    .A1(\RAM[123][2] ),
    .S(_0986_),
    .X(_0494_));
 sky130_fd_sc_hd__mux2_1 _1965_ (.A0(net110),
    .A1(\RAM[123][3] ),
    .S(_0986_),
    .X(_0495_));
 sky130_fd_sc_hd__or2_4 _1966_ (.A(_0862_),
    .B(_0865_),
    .X(_0987_));
 sky130_fd_sc_hd__mux2_1 _1967_ (.A0(net60),
    .A1(\RAM[124][0] ),
    .S(_0987_),
    .X(_0496_));
 sky130_fd_sc_hd__mux2_1 _1968_ (.A0(net40),
    .A1(\RAM[124][1] ),
    .S(_0987_),
    .X(_0497_));
 sky130_fd_sc_hd__mux2_1 _1969_ (.A0(net119),
    .A1(\RAM[124][2] ),
    .S(_0987_),
    .X(_0498_));
 sky130_fd_sc_hd__mux2_1 _1970_ (.A0(net98),
    .A1(\RAM[124][3] ),
    .S(_0987_),
    .X(_0499_));
 sky130_fd_sc_hd__nand2_2 _1971_ (.A(_0855_),
    .B(_0861_),
    .Y(_0988_));
 sky130_fd_sc_hd__mux2_1 _1972_ (.A0(net60),
    .A1(\RAM[125][0] ),
    .S(_0988_),
    .X(_0500_));
 sky130_fd_sc_hd__mux2_1 _1973_ (.A0(net40),
    .A1(\RAM[125][1] ),
    .S(_0988_),
    .X(_0501_));
 sky130_fd_sc_hd__mux2_1 _1974_ (.A0(net113),
    .A1(\RAM[125][2] ),
    .S(_0988_),
    .X(_0502_));
 sky130_fd_sc_hd__mux2_1 _1975_ (.A0(net98),
    .A1(\RAM[125][3] ),
    .S(_0988_),
    .X(_0503_));
 sky130_fd_sc_hd__nand2_2 _1976_ (.A(_0861_),
    .B(_0870_),
    .Y(_0989_));
 sky130_fd_sc_hd__mux2_1 _1977_ (.A0(net56),
    .A1(\RAM[126][0] ),
    .S(_0989_),
    .X(_0504_));
 sky130_fd_sc_hd__mux2_1 _1978_ (.A0(net39),
    .A1(\RAM[126][1] ),
    .S(_0989_),
    .X(_0505_));
 sky130_fd_sc_hd__mux2_1 _1979_ (.A0(net114),
    .A1(\RAM[126][2] ),
    .S(_0989_),
    .X(_0506_));
 sky130_fd_sc_hd__mux2_1 _1980_ (.A0(net96),
    .A1(\RAM[126][3] ),
    .S(_0989_),
    .X(_0507_));
 sky130_fd_sc_hd__nor2_2 _1981_ (.A(_0833_),
    .B(net17),
    .Y(_0990_));
 sky130_fd_sc_hd__mux2_1 _1982_ (.A0(\RAM[9][0] ),
    .A1(net64),
    .S(_0990_),
    .X(_0508_));
 sky130_fd_sc_hd__mux2_1 _1983_ (.A0(\RAM[9][1] ),
    .A1(net49),
    .S(_0990_),
    .X(_0509_));
 sky130_fd_sc_hd__mux2_1 _1984_ (.A0(\RAM[9][2] ),
    .A1(net124),
    .S(_0990_),
    .X(_0510_));
 sky130_fd_sc_hd__mux2_1 _1985_ (.A0(\RAM[9][3] ),
    .A1(net106),
    .S(_0990_),
    .X(_0511_));
 sky130_fd_sc_hd__dfxtp_1 _1986_ (.CLK(clknet_leaf_24_clk),
    .D(_0000_),
    .Q(\RAM[69][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1987_ (.CLK(clknet_leaf_25_clk),
    .D(_0001_),
    .Q(\RAM[69][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1988_ (.CLK(clknet_leaf_26_clk),
    .D(_0002_),
    .Q(\RAM[69][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1989_ (.CLK(clknet_leaf_25_clk),
    .D(_0003_),
    .Q(\RAM[69][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1990_ (.CLK(clknet_leaf_16_clk),
    .D(_0004_),
    .Q(\RAM[89][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1991_ (.CLK(clknet_leaf_19_clk),
    .D(_0005_),
    .Q(\RAM[89][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1992_ (.CLK(clknet_leaf_16_clk),
    .D(_0006_),
    .Q(\RAM[89][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1993_ (.CLK(clknet_leaf_13_clk),
    .D(_0007_),
    .Q(\RAM[89][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1994_ (.CLK(clknet_leaf_3_clk),
    .D(_0008_),
    .Q(\RAM[59][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1995_ (.CLK(clknet_leaf_3_clk),
    .D(_0009_),
    .Q(\RAM[59][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1996_ (.CLK(clknet_leaf_3_clk),
    .D(_0010_),
    .Q(\RAM[59][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1997_ (.CLK(clknet_leaf_3_clk),
    .D(_0011_),
    .Q(\RAM[59][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1998_ (.CLK(clknet_leaf_2_clk),
    .D(_0012_),
    .Q(\RAM[49][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1999_ (.CLK(clknet_leaf_2_clk),
    .D(_0013_),
    .Q(\RAM[49][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2000_ (.CLK(clknet_leaf_6_clk),
    .D(_0014_),
    .Q(\RAM[49][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2001_ (.CLK(clknet_leaf_6_clk),
    .D(_0015_),
    .Q(\RAM[49][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2002_ (.CLK(clknet_leaf_0_clk),
    .D(_0016_),
    .Q(\RAM[39][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2003_ (.CLK(clknet_leaf_44_clk),
    .D(_0017_),
    .Q(\RAM[39][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2004_ (.CLK(clknet_leaf_0_clk),
    .D(_0018_),
    .Q(\RAM[39][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2005_ (.CLK(clknet_leaf_1_clk),
    .D(_0019_),
    .Q(\RAM[39][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2006_ (.CLK(clknet_leaf_10_clk),
    .D(_0020_),
    .Q(\RAM[19][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2007_ (.CLK(clknet_leaf_10_clk),
    .D(_0021_),
    .Q(\RAM[19][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2008_ (.CLK(clknet_leaf_9_clk),
    .D(_0022_),
    .Q(\RAM[19][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2009_ (.CLK(clknet_leaf_9_clk),
    .D(_0023_),
    .Q(\RAM[19][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2010_ (.CLK(clknet_leaf_26_clk),
    .D(_0024_),
    .Q(\RAM[79][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2011_ (.CLK(clknet_leaf_30_clk),
    .D(_0025_),
    .Q(\RAM[79][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2012_ (.CLK(clknet_leaf_29_clk),
    .D(_0026_),
    .Q(\RAM[79][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2013_ (.CLK(clknet_leaf_26_clk),
    .D(_0027_),
    .Q(\RAM[79][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2014_ (.CLK(clknet_leaf_11_clk),
    .D(_0028_),
    .Q(\RAM[29][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2015_ (.CLK(clknet_leaf_9_clk),
    .D(_0029_),
    .Q(\RAM[29][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2016_ (.CLK(clknet_leaf_7_clk),
    .D(_0030_),
    .Q(\RAM[29][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2017_ (.CLK(clknet_leaf_8_clk),
    .D(_0031_),
    .Q(\RAM[29][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2018_ (.CLK(clknet_leaf_37_clk),
    .D(_0032_),
    .Q(\RAM[99][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2019_ (.CLK(clknet_leaf_35_clk),
    .D(_0033_),
    .Q(\RAM[99][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2020_ (.CLK(clknet_leaf_35_clk),
    .D(_0034_),
    .Q(\RAM[99][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2021_ (.CLK(clknet_leaf_36_clk),
    .D(_0035_),
    .Q(\RAM[99][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2022_ (.CLK(clknet_leaf_32_clk),
    .D(_0036_),
    .Q(\RAM[109][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2023_ (.CLK(clknet_leaf_33_clk),
    .D(_0037_),
    .Q(\RAM[109][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2024_ (.CLK(clknet_leaf_33_clk),
    .D(_0038_),
    .Q(\RAM[109][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2025_ (.CLK(clknet_leaf_34_clk),
    .D(_0039_),
    .Q(\RAM[109][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2026_ (.CLK(clknet_leaf_16_clk),
    .D(_0040_),
    .Q(\RAM[119][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2027_ (.CLK(clknet_leaf_4_clk),
    .D(_0041_),
    .Q(\RAM[119][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2028_ (.CLK(clknet_leaf_38_clk),
    .D(_0042_),
    .Q(\RAM[119][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2029_ (.CLK(clknet_leaf_16_clk),
    .D(_0043_),
    .Q(\RAM[119][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2030_ (.CLK(clknet_leaf_41_clk),
    .D(_0044_),
    .Q(\RAM[127][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2031_ (.CLK(clknet_leaf_41_clk),
    .D(_0045_),
    .Q(\RAM[127][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2032_ (.CLK(clknet_leaf_41_clk),
    .D(_0046_),
    .Q(\RAM[127][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2033_ (.CLK(clknet_leaf_41_clk),
    .D(_0047_),
    .Q(\RAM[127][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2034_ (.CLK(clknet_leaf_23_clk),
    .D(_0048_),
    .Q(\RAM[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2035_ (.CLK(clknet_leaf_23_clk),
    .D(_0049_),
    .Q(\RAM[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2036_ (.CLK(clknet_leaf_23_clk),
    .D(_0050_),
    .Q(\RAM[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2037_ (.CLK(clknet_leaf_23_clk),
    .D(_0051_),
    .Q(\RAM[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2038_ (.CLK(clknet_leaf_23_clk),
    .D(_0052_),
    .Q(\RAM[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2039_ (.CLK(clknet_leaf_24_clk),
    .D(_0053_),
    .Q(\RAM[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2040_ (.CLK(clknet_leaf_23_clk),
    .D(_0054_),
    .Q(\RAM[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2041_ (.CLK(clknet_leaf_23_clk),
    .D(_0055_),
    .Q(\RAM[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2042_ (.CLK(clknet_leaf_24_clk),
    .D(_0056_),
    .Q(\RAM[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2043_ (.CLK(clknet_leaf_24_clk),
    .D(_0057_),
    .Q(\RAM[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2044_ (.CLK(clknet_leaf_21_clk),
    .D(_0058_),
    .Q(\RAM[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2045_ (.CLK(clknet_leaf_21_clk),
    .D(_0059_),
    .Q(\RAM[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2046_ (.CLK(clknet_leaf_24_clk),
    .D(_0060_),
    .Q(\RAM[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2047_ (.CLK(clknet_leaf_24_clk),
    .D(_0061_),
    .Q(\RAM[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2048_ (.CLK(clknet_leaf_23_clk),
    .D(_0062_),
    .Q(\RAM[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2049_ (.CLK(clknet_leaf_23_clk),
    .D(_0063_),
    .Q(\RAM[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2050_ (.CLK(clknet_leaf_10_clk),
    .D(_0064_),
    .Q(\RAM[16][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2051_ (.CLK(clknet_leaf_10_clk),
    .D(_0065_),
    .Q(\RAM[16][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2052_ (.CLK(clknet_leaf_10_clk),
    .D(_0066_),
    .Q(\RAM[16][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2053_ (.CLK(clknet_leaf_10_clk),
    .D(_0067_),
    .Q(\RAM[16][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2054_ (.CLK(clknet_leaf_10_clk),
    .D(_0068_),
    .Q(\RAM[17][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2055_ (.CLK(clknet_leaf_10_clk),
    .D(_0069_),
    .Q(\RAM[17][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2056_ (.CLK(clknet_leaf_9_clk),
    .D(_0070_),
    .Q(\RAM[17][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2057_ (.CLK(clknet_leaf_10_clk),
    .D(_0071_),
    .Q(\RAM[17][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2058_ (.CLK(clknet_leaf_10_clk),
    .D(_0072_),
    .Q(\RAM[18][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2059_ (.CLK(clknet_leaf_9_clk),
    .D(_0073_),
    .Q(\RAM[18][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2060_ (.CLK(clknet_leaf_9_clk),
    .D(_0074_),
    .Q(\RAM[18][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2061_ (.CLK(clknet_leaf_9_clk),
    .D(_0075_),
    .Q(\RAM[18][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2062_ (.CLK(clknet_leaf_20_clk),
    .D(_0076_),
    .Q(\RAM[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2063_ (.CLK(clknet_leaf_20_clk),
    .D(_0077_),
    .Q(\RAM[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2064_ (.CLK(clknet_leaf_21_clk),
    .D(_0078_),
    .Q(\RAM[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2065_ (.CLK(clknet_leaf_20_clk),
    .D(_0079_),
    .Q(\RAM[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2066_ (.CLK(clknet_leaf_12_clk),
    .D(_0080_),
    .Q(\RAM[20][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2067_ (.CLK(clknet_leaf_12_clk),
    .D(_0081_),
    .Q(\RAM[20][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2068_ (.CLK(clknet_leaf_13_clk),
    .D(_0082_),
    .Q(\RAM[20][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2069_ (.CLK(clknet_leaf_13_clk),
    .D(_0083_),
    .Q(\RAM[20][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2070_ (.CLK(clknet_leaf_13_clk),
    .D(_0084_),
    .Q(\RAM[21][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2071_ (.CLK(clknet_leaf_12_clk),
    .D(_0085_),
    .Q(\RAM[21][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2072_ (.CLK(clknet_leaf_14_clk),
    .D(_0086_),
    .Q(\RAM[21][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2073_ (.CLK(clknet_leaf_12_clk),
    .D(_0087_),
    .Q(\RAM[21][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2074_ (.CLK(clknet_leaf_12_clk),
    .D(_0088_),
    .Q(\RAM[22][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2075_ (.CLK(clknet_leaf_12_clk),
    .D(_0089_),
    .Q(\RAM[22][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2076_ (.CLK(clknet_leaf_14_clk),
    .D(_0090_),
    .Q(\RAM[22][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2077_ (.CLK(clknet_leaf_11_clk),
    .D(_0091_),
    .Q(\RAM[22][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2078_ (.CLK(clknet_leaf_12_clk),
    .D(_0092_),
    .Q(\RAM[23][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2079_ (.CLK(clknet_leaf_12_clk),
    .D(_0093_),
    .Q(\RAM[23][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2080_ (.CLK(clknet_leaf_14_clk),
    .D(_0094_),
    .Q(\RAM[23][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2081_ (.CLK(clknet_leaf_11_clk),
    .D(_0095_),
    .Q(\RAM[23][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2082_ (.CLK(clknet_leaf_11_clk),
    .D(_0096_),
    .Q(\RAM[24][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2083_ (.CLK(clknet_leaf_11_clk),
    .D(_0097_),
    .Q(\RAM[24][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2084_ (.CLK(clknet_leaf_14_clk),
    .D(_0098_),
    .Q(\RAM[24][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2085_ (.CLK(clknet_leaf_11_clk),
    .D(_0099_),
    .Q(\RAM[24][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2086_ (.CLK(clknet_leaf_10_clk),
    .D(_0100_),
    .Q(\RAM[25][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2087_ (.CLK(clknet_leaf_12_clk),
    .D(_0101_),
    .Q(\RAM[25][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2088_ (.CLK(clknet_leaf_11_clk),
    .D(_0102_),
    .Q(\RAM[25][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2089_ (.CLK(clknet_leaf_11_clk),
    .D(_0103_),
    .Q(\RAM[25][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2090_ (.CLK(clknet_leaf_11_clk),
    .D(_0104_),
    .Q(\RAM[26][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2091_ (.CLK(clknet_leaf_11_clk),
    .D(_0105_),
    .Q(\RAM[26][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2092_ (.CLK(clknet_leaf_8_clk),
    .D(_0106_),
    .Q(\RAM[26][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2093_ (.CLK(clknet_leaf_11_clk),
    .D(_0107_),
    .Q(\RAM[26][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2094_ (.CLK(clknet_leaf_10_clk),
    .D(_0108_),
    .Q(\RAM[27][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2095_ (.CLK(clknet_leaf_11_clk),
    .D(_0109_),
    .Q(\RAM[27][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2096_ (.CLK(clknet_leaf_11_clk),
    .D(_0110_),
    .Q(\RAM[27][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2097_ (.CLK(clknet_leaf_11_clk),
    .D(_0111_),
    .Q(\RAM[27][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2098_ (.CLK(clknet_leaf_8_clk),
    .D(_0112_),
    .Q(\RAM[28][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2099_ (.CLK(clknet_leaf_8_clk),
    .D(_0113_),
    .Q(\RAM[28][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2100_ (.CLK(clknet_leaf_7_clk),
    .D(_0114_),
    .Q(\RAM[28][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2101_ (.CLK(clknet_leaf_8_clk),
    .D(_0115_),
    .Q(\RAM[28][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2102_ (.CLK(clknet_leaf_19_clk),
    .D(_0116_),
    .Q(\RAM[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2103_ (.CLK(clknet_leaf_20_clk),
    .D(_0117_),
    .Q(\RAM[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2104_ (.CLK(clknet_leaf_21_clk),
    .D(_0118_),
    .Q(\RAM[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2105_ (.CLK(clknet_leaf_20_clk),
    .D(_0119_),
    .Q(\RAM[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2106_ (.CLK(clknet_leaf_8_clk),
    .D(_0120_),
    .Q(\RAM[30][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2107_ (.CLK(clknet_leaf_9_clk),
    .D(_0121_),
    .Q(\RAM[30][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2108_ (.CLK(clknet_leaf_9_clk),
    .D(_0122_),
    .Q(\RAM[30][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2109_ (.CLK(clknet_leaf_9_clk),
    .D(_0123_),
    .Q(\RAM[30][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2110_ (.CLK(clknet_leaf_8_clk),
    .D(_0124_),
    .Q(\RAM[31][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2111_ (.CLK(clknet_leaf_9_clk),
    .D(_0125_),
    .Q(\RAM[31][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2112_ (.CLK(clknet_leaf_7_clk),
    .D(_0126_),
    .Q(\RAM[31][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2113_ (.CLK(clknet_leaf_9_clk),
    .D(_0127_),
    .Q(\RAM[31][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2114_ (.CLK(clknet_leaf_3_clk),
    .D(_0128_),
    .Q(\RAM[32][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2115_ (.CLK(clknet_leaf_43_clk),
    .D(_0129_),
    .Q(\RAM[32][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2116_ (.CLK(clknet_leaf_42_clk),
    .D(_0130_),
    .Q(\RAM[32][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2117_ (.CLK(clknet_leaf_40_clk),
    .D(_0131_),
    .Q(\RAM[32][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2118_ (.CLK(clknet_leaf_0_clk),
    .D(_0132_),
    .Q(\RAM[33][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2119_ (.CLK(clknet_leaf_42_clk),
    .D(_0133_),
    .Q(\RAM[33][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2120_ (.CLK(clknet_leaf_43_clk),
    .D(_0134_),
    .Q(\RAM[33][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2121_ (.CLK(clknet_leaf_39_clk),
    .D(_0135_),
    .Q(\RAM[33][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2122_ (.CLK(clknet_leaf_0_clk),
    .D(_0136_),
    .Q(\RAM[34][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2123_ (.CLK(clknet_leaf_43_clk),
    .D(_0137_),
    .Q(\RAM[34][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2124_ (.CLK(clknet_leaf_0_clk),
    .D(_0138_),
    .Q(\RAM[34][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2125_ (.CLK(clknet_leaf_0_clk),
    .D(_0139_),
    .Q(\RAM[34][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2126_ (.CLK(clknet_leaf_0_clk),
    .D(_0140_),
    .Q(\RAM[35][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2127_ (.CLK(clknet_leaf_43_clk),
    .D(_0141_),
    .Q(\RAM[35][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2128_ (.CLK(clknet_leaf_0_clk),
    .D(_0142_),
    .Q(\RAM[35][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2129_ (.CLK(clknet_leaf_0_clk),
    .D(_0143_),
    .Q(\RAM[35][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2130_ (.CLK(clknet_leaf_0_clk),
    .D(_0144_),
    .Q(\RAM[36][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2131_ (.CLK(clknet_leaf_44_clk),
    .D(_0145_),
    .Q(\RAM[36][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2132_ (.CLK(clknet_leaf_0_clk),
    .D(_0146_),
    .Q(\RAM[36][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2133_ (.CLK(clknet_leaf_0_clk),
    .D(_0147_),
    .Q(\RAM[36][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2134_ (.CLK(clknet_leaf_0_clk),
    .D(_0148_),
    .Q(\RAM[37][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2135_ (.CLK(clknet_leaf_44_clk),
    .D(_0149_),
    .Q(\RAM[37][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2136_ (.CLK(clknet_leaf_0_clk),
    .D(_0150_),
    .Q(\RAM[37][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2137_ (.CLK(clknet_leaf_1_clk),
    .D(_0151_),
    .Q(\RAM[37][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2138_ (.CLK(clknet_leaf_0_clk),
    .D(_0152_),
    .Q(\RAM[38][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2139_ (.CLK(clknet_leaf_44_clk),
    .D(_0153_),
    .Q(\RAM[38][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2140_ (.CLK(clknet_leaf_0_clk),
    .D(_0154_),
    .Q(\RAM[38][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2141_ (.CLK(clknet_leaf_44_clk),
    .D(_0155_),
    .Q(\RAM[38][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2142_ (.CLK(clknet_leaf_19_clk),
    .D(_0156_),
    .Q(\RAM[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2143_ (.CLK(clknet_leaf_20_clk),
    .D(_0157_),
    .Q(\RAM[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2144_ (.CLK(clknet_leaf_21_clk),
    .D(_0158_),
    .Q(\RAM[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2145_ (.CLK(clknet_leaf_20_clk),
    .D(_0159_),
    .Q(\RAM[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2146_ (.CLK(clknet_leaf_41_clk),
    .D(_0160_),
    .Q(\RAM[40][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2147_ (.CLK(clknet_leaf_41_clk),
    .D(_0161_),
    .Q(\RAM[40][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2148_ (.CLK(clknet_leaf_42_clk),
    .D(_0162_),
    .Q(\RAM[40][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2149_ (.CLK(clknet_leaf_42_clk),
    .D(_0163_),
    .Q(\RAM[40][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2150_ (.CLK(clknet_leaf_40_clk),
    .D(_0164_),
    .Q(\RAM[41][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2151_ (.CLK(clknet_leaf_41_clk),
    .D(_0165_),
    .Q(\RAM[41][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2152_ (.CLK(clknet_leaf_42_clk),
    .D(_0166_),
    .Q(\RAM[41][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2153_ (.CLK(clknet_leaf_42_clk),
    .D(_0167_),
    .Q(\RAM[41][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2154_ (.CLK(clknet_leaf_42_clk),
    .D(_0168_),
    .Q(\RAM[42][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2155_ (.CLK(clknet_leaf_42_clk),
    .D(_0169_),
    .Q(\RAM[42][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2156_ (.CLK(clknet_leaf_43_clk),
    .D(_0170_),
    .Q(\RAM[42][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2157_ (.CLK(clknet_leaf_39_clk),
    .D(_0171_),
    .Q(\RAM[42][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2158_ (.CLK(clknet_leaf_42_clk),
    .D(_0172_),
    .Q(\RAM[43][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2159_ (.CLK(clknet_leaf_42_clk),
    .D(_0173_),
    .Q(\RAM[43][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2160_ (.CLK(clknet_leaf_43_clk),
    .D(_0174_),
    .Q(\RAM[43][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2161_ (.CLK(clknet_leaf_40_clk),
    .D(_0175_),
    .Q(\RAM[43][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2162_ (.CLK(clknet_leaf_44_clk),
    .D(_0176_),
    .Q(\RAM[44][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2163_ (.CLK(clknet_leaf_43_clk),
    .D(_0177_),
    .Q(\RAM[44][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2164_ (.CLK(clknet_leaf_43_clk),
    .D(_0178_),
    .Q(\RAM[44][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2165_ (.CLK(clknet_leaf_43_clk),
    .D(_0179_),
    .Q(\RAM[44][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2166_ (.CLK(clknet_leaf_44_clk),
    .D(_0180_),
    .Q(\RAM[45][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2167_ (.CLK(clknet_leaf_43_clk),
    .D(_0181_),
    .Q(\RAM[45][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2168_ (.CLK(clknet_leaf_43_clk),
    .D(_0182_),
    .Q(\RAM[45][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2169_ (.CLK(clknet_leaf_43_clk),
    .D(_0183_),
    .Q(\RAM[45][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2170_ (.CLK(clknet_leaf_44_clk),
    .D(_0184_),
    .Q(\RAM[46][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2171_ (.CLK(clknet_leaf_44_clk),
    .D(_0185_),
    .Q(\RAM[46][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2172_ (.CLK(clknet_leaf_43_clk),
    .D(_0186_),
    .Q(\RAM[46][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2173_ (.CLK(clknet_leaf_44_clk),
    .D(_0187_),
    .Q(\RAM[46][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2174_ (.CLK(clknet_leaf_44_clk),
    .D(_0188_),
    .Q(\RAM[47][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2175_ (.CLK(clknet_leaf_44_clk),
    .D(_0189_),
    .Q(\RAM[47][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2176_ (.CLK(clknet_leaf_43_clk),
    .D(_0190_),
    .Q(\RAM[47][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2177_ (.CLK(clknet_leaf_44_clk),
    .D(_0191_),
    .Q(\RAM[47][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2178_ (.CLK(clknet_leaf_2_clk),
    .D(_0192_),
    .Q(\RAM[48][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2179_ (.CLK(clknet_leaf_2_clk),
    .D(_0193_),
    .Q(\RAM[48][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2180_ (.CLK(clknet_leaf_6_clk),
    .D(_0194_),
    .Q(\RAM[48][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2181_ (.CLK(clknet_leaf_5_clk),
    .D(_0195_),
    .Q(\RAM[48][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2182_ (.CLK(clknet_leaf_22_clk),
    .D(_0196_),
    .Q(\RAM[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2183_ (.CLK(clknet_leaf_22_clk),
    .D(_0197_),
    .Q(\RAM[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2184_ (.CLK(clknet_leaf_22_clk),
    .D(_0198_),
    .Q(\RAM[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2185_ (.CLK(clknet_leaf_22_clk),
    .D(_0199_),
    .Q(\RAM[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2186_ (.CLK(clknet_leaf_2_clk),
    .D(_0200_),
    .Q(\RAM[50][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2187_ (.CLK(clknet_leaf_2_clk),
    .D(_0201_),
    .Q(\RAM[50][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2188_ (.CLK(clknet_leaf_6_clk),
    .D(_0202_),
    .Q(\RAM[50][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2189_ (.CLK(clknet_leaf_6_clk),
    .D(_0203_),
    .Q(\RAM[50][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2190_ (.CLK(clknet_leaf_1_clk),
    .D(_0204_),
    .Q(\RAM[51][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2191_ (.CLK(clknet_leaf_2_clk),
    .D(_0205_),
    .Q(\RAM[51][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2192_ (.CLK(clknet_leaf_6_clk),
    .D(_0206_),
    .Q(\RAM[51][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2193_ (.CLK(clknet_leaf_6_clk),
    .D(_0207_),
    .Q(\RAM[51][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2194_ (.CLK(clknet_leaf_4_clk),
    .D(_0208_),
    .Q(\RAM[52][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2195_ (.CLK(clknet_leaf_4_clk),
    .D(_0209_),
    .Q(\RAM[52][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2196_ (.CLK(clknet_leaf_4_clk),
    .D(_0210_),
    .Q(\RAM[52][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2197_ (.CLK(clknet_leaf_5_clk),
    .D(_0211_),
    .Q(\RAM[52][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2198_ (.CLK(clknet_leaf_4_clk),
    .D(_0212_),
    .Q(\RAM[53][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2199_ (.CLK(clknet_leaf_4_clk),
    .D(_0213_),
    .Q(\RAM[53][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2200_ (.CLK(clknet_leaf_4_clk),
    .D(_0214_),
    .Q(\RAM[53][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2201_ (.CLK(clknet_leaf_16_clk),
    .D(_0215_),
    .Q(\RAM[53][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2202_ (.CLK(clknet_leaf_3_clk),
    .D(_0216_),
    .Q(\RAM[54][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2203_ (.CLK(clknet_leaf_5_clk),
    .D(_0217_),
    .Q(\RAM[54][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2204_ (.CLK(clknet_leaf_5_clk),
    .D(_0218_),
    .Q(\RAM[54][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2205_ (.CLK(clknet_leaf_5_clk),
    .D(_0219_),
    .Q(\RAM[54][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2206_ (.CLK(clknet_leaf_3_clk),
    .D(_0220_),
    .Q(\RAM[55][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2207_ (.CLK(clknet_leaf_4_clk),
    .D(_0221_),
    .Q(\RAM[55][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2208_ (.CLK(clknet_leaf_5_clk),
    .D(_0222_),
    .Q(\RAM[55][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2209_ (.CLK(clknet_leaf_5_clk),
    .D(_0223_),
    .Q(\RAM[55][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2210_ (.CLK(clknet_leaf_39_clk),
    .D(_0224_),
    .Q(\RAM[56][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2211_ (.CLK(clknet_leaf_38_clk),
    .D(_0225_),
    .Q(\RAM[56][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2212_ (.CLK(clknet_leaf_3_clk),
    .D(_0226_),
    .Q(\RAM[56][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2213_ (.CLK(clknet_leaf_3_clk),
    .D(_0227_),
    .Q(\RAM[56][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2214_ (.CLK(clknet_leaf_38_clk),
    .D(_0228_),
    .Q(\RAM[57][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2215_ (.CLK(clknet_leaf_38_clk),
    .D(_0229_),
    .Q(\RAM[57][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2216_ (.CLK(clknet_leaf_3_clk),
    .D(_0230_),
    .Q(\RAM[57][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2217_ (.CLK(clknet_leaf_3_clk),
    .D(_0231_),
    .Q(\RAM[57][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2218_ (.CLK(clknet_leaf_3_clk),
    .D(_0232_),
    .Q(\RAM[58][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2219_ (.CLK(clknet_leaf_3_clk),
    .D(_0233_),
    .Q(\RAM[58][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2220_ (.CLK(clknet_leaf_3_clk),
    .D(_0234_),
    .Q(\RAM[58][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2221_ (.CLK(clknet_leaf_3_clk),
    .D(_0235_),
    .Q(\RAM[58][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2222_ (.CLK(clknet_leaf_22_clk),
    .D(_0236_),
    .Q(\RAM[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2223_ (.CLK(clknet_leaf_22_clk),
    .D(_0237_),
    .Q(\RAM[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2224_ (.CLK(clknet_leaf_22_clk),
    .D(_0238_),
    .Q(\RAM[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2225_ (.CLK(clknet_leaf_22_clk),
    .D(_0239_),
    .Q(\RAM[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2226_ (.CLK(clknet_leaf_1_clk),
    .D(_0240_),
    .Q(\RAM[60][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2227_ (.CLK(clknet_leaf_1_clk),
    .D(_0241_),
    .Q(\RAM[60][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2228_ (.CLK(clknet_leaf_3_clk),
    .D(_0242_),
    .Q(\RAM[60][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2229_ (.CLK(clknet_leaf_3_clk),
    .D(_0243_),
    .Q(\RAM[60][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2230_ (.CLK(clknet_leaf_1_clk),
    .D(_0244_),
    .Q(\RAM[61][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2231_ (.CLK(clknet_leaf_1_clk),
    .D(_0245_),
    .Q(\RAM[61][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2232_ (.CLK(clknet_leaf_0_clk),
    .D(_0246_),
    .Q(\RAM[61][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2233_ (.CLK(clknet_leaf_2_clk),
    .D(_0247_),
    .Q(\RAM[61][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2234_ (.CLK(clknet_leaf_1_clk),
    .D(_0248_),
    .Q(\RAM[62][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2235_ (.CLK(clknet_leaf_1_clk),
    .D(_0249_),
    .Q(\RAM[62][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2236_ (.CLK(clknet_leaf_1_clk),
    .D(_0250_),
    .Q(\RAM[62][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2237_ (.CLK(clknet_leaf_2_clk),
    .D(_0251_),
    .Q(\RAM[62][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2238_ (.CLK(clknet_leaf_1_clk),
    .D(_0252_),
    .Q(\RAM[63][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2239_ (.CLK(clknet_leaf_1_clk),
    .D(_0253_),
    .Q(\RAM[63][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2240_ (.CLK(clknet_leaf_1_clk),
    .D(_0254_),
    .Q(\RAM[63][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2241_ (.CLK(clknet_leaf_2_clk),
    .D(_0255_),
    .Q(\RAM[63][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2242_ (.CLK(clknet_leaf_27_clk),
    .D(_0256_),
    .Q(\RAM[64][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2243_ (.CLK(clknet_leaf_26_clk),
    .D(_0257_),
    .Q(\RAM[64][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2244_ (.CLK(clknet_leaf_29_clk),
    .D(_0258_),
    .Q(\RAM[64][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2245_ (.CLK(clknet_leaf_26_clk),
    .D(_0259_),
    .Q(\RAM[64][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2246_ (.CLK(clknet_leaf_17_clk),
    .D(_0260_),
    .Q(\RAM[65][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2247_ (.CLK(clknet_leaf_27_clk),
    .D(_0261_),
    .Q(\RAM[65][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2248_ (.CLK(clknet_leaf_28_clk),
    .D(_0262_),
    .Q(\RAM[65][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2249_ (.CLK(clknet_leaf_27_clk),
    .D(_0263_),
    .Q(\RAM[65][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2250_ (.CLK(clknet_leaf_16_clk),
    .D(_0264_),
    .Q(\RAM[66][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2251_ (.CLK(clknet_leaf_28_clk),
    .D(_0265_),
    .Q(\RAM[66][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2252_ (.CLK(clknet_leaf_28_clk),
    .D(_0266_),
    .Q(\RAM[66][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2253_ (.CLK(clknet_leaf_27_clk),
    .D(_0267_),
    .Q(\RAM[66][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2254_ (.CLK(clknet_leaf_16_clk),
    .D(_0268_),
    .Q(\RAM[67][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2255_ (.CLK(clknet_leaf_28_clk),
    .D(_0269_),
    .Q(\RAM[67][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2256_ (.CLK(clknet_leaf_28_clk),
    .D(_0270_),
    .Q(\RAM[67][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2257_ (.CLK(clknet_leaf_27_clk),
    .D(_0271_),
    .Q(\RAM[67][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2258_ (.CLK(clknet_leaf_24_clk),
    .D(_0272_),
    .Q(\RAM[68][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2259_ (.CLK(clknet_leaf_24_clk),
    .D(_0273_),
    .Q(\RAM[68][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2260_ (.CLK(clknet_leaf_26_clk),
    .D(_0274_),
    .Q(\RAM[68][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2261_ (.CLK(clknet_leaf_24_clk),
    .D(_0275_),
    .Q(\RAM[68][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2262_ (.CLK(clknet_leaf_22_clk),
    .D(_0276_),
    .Q(\RAM[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2263_ (.CLK(clknet_leaf_22_clk),
    .D(_0277_),
    .Q(\RAM[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2264_ (.CLK(clknet_leaf_21_clk),
    .D(_0278_),
    .Q(\RAM[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2265_ (.CLK(clknet_leaf_21_clk),
    .D(_0279_),
    .Q(\RAM[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2266_ (.CLK(clknet_leaf_27_clk),
    .D(_0280_),
    .Q(\RAM[70][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2267_ (.CLK(clknet_leaf_26_clk),
    .D(_0281_),
    .Q(\RAM[70][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2268_ (.CLK(clknet_leaf_26_clk),
    .D(_0282_),
    .Q(\RAM[70][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2269_ (.CLK(clknet_leaf_25_clk),
    .D(_0283_),
    .Q(\RAM[70][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2270_ (.CLK(clknet_leaf_27_clk),
    .D(_0284_),
    .Q(\RAM[71][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2271_ (.CLK(clknet_leaf_25_clk),
    .D(_0285_),
    .Q(\RAM[71][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2272_ (.CLK(clknet_leaf_26_clk),
    .D(_0286_),
    .Q(\RAM[71][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2273_ (.CLK(clknet_leaf_25_clk),
    .D(_0287_),
    .Q(\RAM[71][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2274_ (.CLK(clknet_leaf_30_clk),
    .D(_0288_),
    .Q(\RAM[72][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2275_ (.CLK(clknet_leaf_31_clk),
    .D(_0289_),
    .Q(\RAM[72][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2276_ (.CLK(clknet_leaf_29_clk),
    .D(_0290_),
    .Q(\RAM[72][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2277_ (.CLK(clknet_leaf_31_clk),
    .D(_0291_),
    .Q(\RAM[72][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2278_ (.CLK(clknet_leaf_30_clk),
    .D(_0292_),
    .Q(\RAM[73][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2279_ (.CLK(clknet_leaf_29_clk),
    .D(_0293_),
    .Q(\RAM[73][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2280_ (.CLK(clknet_leaf_29_clk),
    .D(_0294_),
    .Q(\RAM[73][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2281_ (.CLK(clknet_leaf_30_clk),
    .D(_0295_),
    .Q(\RAM[73][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2282_ (.CLK(clknet_leaf_29_clk),
    .D(_0296_),
    .Q(\RAM[74][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2283_ (.CLK(clknet_leaf_29_clk),
    .D(_0297_),
    .Q(\RAM[74][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2284_ (.CLK(clknet_leaf_29_clk),
    .D(_0298_),
    .Q(\RAM[74][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2285_ (.CLK(clknet_leaf_31_clk),
    .D(_0299_),
    .Q(\RAM[74][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2286_ (.CLK(clknet_leaf_30_clk),
    .D(_0300_),
    .Q(\RAM[75][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2287_ (.CLK(clknet_leaf_29_clk),
    .D(_0301_),
    .Q(\RAM[75][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2288_ (.CLK(clknet_leaf_29_clk),
    .D(_0302_),
    .Q(\RAM[75][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2289_ (.CLK(clknet_leaf_31_clk),
    .D(_0303_),
    .Q(\RAM[75][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2290_ (.CLK(clknet_leaf_26_clk),
    .D(_0304_),
    .Q(\RAM[76][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2291_ (.CLK(clknet_leaf_30_clk),
    .D(_0305_),
    .Q(\RAM[76][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2292_ (.CLK(clknet_leaf_30_clk),
    .D(_0306_),
    .Q(\RAM[76][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2293_ (.CLK(clknet_leaf_25_clk),
    .D(_0307_),
    .Q(\RAM[76][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2294_ (.CLK(clknet_leaf_25_clk),
    .D(_0308_),
    .Q(\RAM[77][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2295_ (.CLK(clknet_leaf_30_clk),
    .D(_0309_),
    .Q(\RAM[77][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2296_ (.CLK(clknet_leaf_30_clk),
    .D(_0310_),
    .Q(\RAM[77][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2297_ (.CLK(clknet_leaf_25_clk),
    .D(_0311_),
    .Q(\RAM[77][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2298_ (.CLK(clknet_leaf_26_clk),
    .D(_0312_),
    .Q(\RAM[78][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2299_ (.CLK(clknet_leaf_26_clk),
    .D(_0313_),
    .Q(\RAM[78][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2300_ (.CLK(clknet_leaf_28_clk),
    .D(_0314_),
    .Q(\RAM[78][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2301_ (.CLK(clknet_leaf_26_clk),
    .D(_0315_),
    .Q(\RAM[78][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2302_ (.CLK(clknet_leaf_22_clk),
    .D(_0316_),
    .Q(\RAM[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2303_ (.CLK(clknet_leaf_20_clk),
    .D(_0317_),
    .Q(\RAM[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2304_ (.CLK(clknet_leaf_21_clk),
    .D(_0318_),
    .Q(\RAM[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2305_ (.CLK(clknet_leaf_21_clk),
    .D(_0319_),
    .Q(\RAM[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2306_ (.CLK(clknet_leaf_5_clk),
    .D(_0320_),
    .Q(\RAM[80][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2307_ (.CLK(clknet_leaf_6_clk),
    .D(_0321_),
    .Q(\RAM[80][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2308_ (.CLK(clknet_leaf_6_clk),
    .D(_0322_),
    .Q(\RAM[80][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2309_ (.CLK(clknet_leaf_7_clk),
    .D(_0323_),
    .Q(\RAM[80][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2310_ (.CLK(clknet_leaf_6_clk),
    .D(_0324_),
    .Q(\RAM[81][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2311_ (.CLK(clknet_leaf_7_clk),
    .D(_0325_),
    .Q(\RAM[81][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2312_ (.CLK(clknet_leaf_6_clk),
    .D(_0326_),
    .Q(\RAM[81][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2313_ (.CLK(clknet_leaf_7_clk),
    .D(_0327_),
    .Q(\RAM[81][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2314_ (.CLK(clknet_leaf_6_clk),
    .D(_0328_),
    .Q(\RAM[82][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2315_ (.CLK(clknet_leaf_7_clk),
    .D(_0329_),
    .Q(\RAM[82][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2316_ (.CLK(clknet_leaf_6_clk),
    .D(_0330_),
    .Q(\RAM[82][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2317_ (.CLK(clknet_leaf_7_clk),
    .D(_0331_),
    .Q(\RAM[82][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2318_ (.CLK(clknet_leaf_6_clk),
    .D(_0332_),
    .Q(\RAM[83][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2319_ (.CLK(clknet_leaf_7_clk),
    .D(_0333_),
    .Q(\RAM[83][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2320_ (.CLK(clknet_leaf_6_clk),
    .D(_0334_),
    .Q(\RAM[83][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2321_ (.CLK(clknet_leaf_7_clk),
    .D(_0335_),
    .Q(\RAM[83][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2322_ (.CLK(clknet_leaf_19_clk),
    .D(_0336_),
    .Q(\RAM[84][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2323_ (.CLK(clknet_leaf_20_clk),
    .D(_0337_),
    .Q(\RAM[84][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2324_ (.CLK(clknet_leaf_19_clk),
    .D(_0338_),
    .Q(\RAM[84][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2325_ (.CLK(clknet_leaf_20_clk),
    .D(_0339_),
    .Q(\RAM[84][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2326_ (.CLK(clknet_leaf_13_clk),
    .D(_0340_),
    .Q(\RAM[85][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2327_ (.CLK(clknet_leaf_13_clk),
    .D(_0341_),
    .Q(\RAM[85][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2328_ (.CLK(clknet_leaf_19_clk),
    .D(_0342_),
    .Q(\RAM[85][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2329_ (.CLK(clknet_leaf_19_clk),
    .D(_0343_),
    .Q(\RAM[85][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2330_ (.CLK(clknet_leaf_13_clk),
    .D(_0344_),
    .Q(\RAM[86][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2331_ (.CLK(clknet_leaf_12_clk),
    .D(_0345_),
    .Q(\RAM[86][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2332_ (.CLK(clknet_leaf_13_clk),
    .D(_0346_),
    .Q(\RAM[86][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2333_ (.CLK(clknet_leaf_13_clk),
    .D(_0347_),
    .Q(\RAM[86][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2334_ (.CLK(clknet_leaf_13_clk),
    .D(_0348_),
    .Q(\RAM[87][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2335_ (.CLK(clknet_leaf_12_clk),
    .D(_0349_),
    .Q(\RAM[87][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2336_ (.CLK(clknet_leaf_13_clk),
    .D(_0350_),
    .Q(\RAM[87][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2337_ (.CLK(clknet_leaf_13_clk),
    .D(_0351_),
    .Q(\RAM[87][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2338_ (.CLK(clknet_leaf_17_clk),
    .D(_0352_),
    .Q(\RAM[88][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2339_ (.CLK(clknet_leaf_17_clk),
    .D(_0353_),
    .Q(\RAM[88][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2340_ (.CLK(clknet_leaf_17_clk),
    .D(_0354_),
    .Q(\RAM[88][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2341_ (.CLK(clknet_leaf_18_clk),
    .D(_0355_),
    .Q(\RAM[88][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2342_ (.CLK(clknet_leaf_18_clk),
    .D(_0356_),
    .Q(\RAM[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2343_ (.CLK(clknet_leaf_27_clk),
    .D(_0357_),
    .Q(\RAM[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2344_ (.CLK(clknet_leaf_21_clk),
    .D(_0358_),
    .Q(\RAM[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2345_ (.CLK(clknet_leaf_18_clk),
    .D(_0359_),
    .Q(\RAM[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2346_ (.CLK(clknet_leaf_15_clk),
    .D(_0360_),
    .Q(\RAM[90][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2347_ (.CLK(clknet_leaf_15_clk),
    .D(_0361_),
    .Q(\RAM[90][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2348_ (.CLK(clknet_leaf_15_clk),
    .D(_0362_),
    .Q(\RAM[90][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2349_ (.CLK(clknet_leaf_14_clk),
    .D(_0363_),
    .Q(\RAM[90][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2350_ (.CLK(clknet_leaf_15_clk),
    .D(_0364_),
    .Q(\RAM[91][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2351_ (.CLK(clknet_leaf_15_clk),
    .D(_0365_),
    .Q(\RAM[91][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2352_ (.CLK(clknet_leaf_16_clk),
    .D(_0366_),
    .Q(\RAM[91][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2353_ (.CLK(clknet_leaf_15_clk),
    .D(_0367_),
    .Q(\RAM[91][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2354_ (.CLK(clknet_leaf_15_clk),
    .D(_0368_),
    .Q(\RAM[92][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2355_ (.CLK(clknet_leaf_15_clk),
    .D(_0369_),
    .Q(\RAM[92][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2356_ (.CLK(clknet_leaf_5_clk),
    .D(_0370_),
    .Q(\RAM[92][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2357_ (.CLK(clknet_leaf_15_clk),
    .D(_0371_),
    .Q(\RAM[92][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2358_ (.CLK(clknet_leaf_5_clk),
    .D(_0372_),
    .Q(\RAM[93][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2359_ (.CLK(clknet_leaf_8_clk),
    .D(_0373_),
    .Q(\RAM[93][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2360_ (.CLK(clknet_leaf_5_clk),
    .D(_0374_),
    .Q(\RAM[93][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2361_ (.CLK(clknet_leaf_15_clk),
    .D(_0375_),
    .Q(\RAM[93][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2362_ (.CLK(clknet_leaf_5_clk),
    .D(_0376_),
    .Q(\RAM[94][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2363_ (.CLK(clknet_leaf_7_clk),
    .D(_0377_),
    .Q(\RAM[94][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2364_ (.CLK(clknet_leaf_5_clk),
    .D(_0378_),
    .Q(\RAM[94][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2365_ (.CLK(clknet_leaf_15_clk),
    .D(_0379_),
    .Q(\RAM[94][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2366_ (.CLK(clknet_leaf_5_clk),
    .D(_0380_),
    .Q(\RAM[95][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2367_ (.CLK(clknet_leaf_8_clk),
    .D(_0381_),
    .Q(\RAM[95][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2368_ (.CLK(clknet_leaf_5_clk),
    .D(_0382_),
    .Q(\RAM[95][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2369_ (.CLK(clknet_leaf_15_clk),
    .D(_0383_),
    .Q(\RAM[95][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2370_ (.CLK(clknet_leaf_36_clk),
    .D(_0384_),
    .Q(\RAM[96][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2371_ (.CLK(clknet_leaf_34_clk),
    .D(_0385_),
    .Q(\RAM[96][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2372_ (.CLK(clknet_leaf_35_clk),
    .D(_0386_),
    .Q(\RAM[96][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2373_ (.CLK(clknet_leaf_36_clk),
    .D(_0387_),
    .Q(\RAM[96][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2374_ (.CLK(clknet_leaf_36_clk),
    .D(_0388_),
    .Q(\RAM[97][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2375_ (.CLK(clknet_leaf_35_clk),
    .D(_0389_),
    .Q(\RAM[97][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2376_ (.CLK(clknet_leaf_35_clk),
    .D(_0390_),
    .Q(\RAM[97][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2377_ (.CLK(clknet_leaf_35_clk),
    .D(_0391_),
    .Q(\RAM[97][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2378_ (.CLK(clknet_leaf_36_clk),
    .D(_0392_),
    .Q(\RAM[98][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2379_ (.CLK(clknet_leaf_35_clk),
    .D(_0393_),
    .Q(\RAM[98][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2380_ (.CLK(clknet_leaf_35_clk),
    .D(_0394_),
    .Q(\RAM[98][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2381_ (.CLK(clknet_leaf_36_clk),
    .D(_0395_),
    .Q(\RAM[98][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2382_ (.CLK(clknet_leaf_20_clk),
    .D(_0396_),
    .Q(\RAM[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2383_ (.CLK(clknet_leaf_21_clk),
    .D(_0397_),
    .Q(\RAM[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2384_ (.CLK(clknet_leaf_21_clk),
    .D(_0398_),
    .Q(\RAM[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2385_ (.CLK(clknet_leaf_20_clk),
    .D(_0399_),
    .Q(\RAM[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2386_ (.CLK(clknet_leaf_34_clk),
    .D(_0400_),
    .Q(\RAM[100][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2387_ (.CLK(clknet_leaf_34_clk),
    .D(_0401_),
    .Q(\RAM[100][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2388_ (.CLK(clknet_leaf_34_clk),
    .D(_0402_),
    .Q(\RAM[100][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2389_ (.CLK(clknet_leaf_34_clk),
    .D(_0403_),
    .Q(\RAM[100][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2390_ (.CLK(clknet_leaf_37_clk),
    .D(_0404_),
    .Q(\RAM[101][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2391_ (.CLK(clknet_leaf_34_clk),
    .D(_0405_),
    .Q(\RAM[101][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2392_ (.CLK(clknet_leaf_34_clk),
    .D(_0406_),
    .Q(\RAM[101][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2393_ (.CLK(clknet_leaf_34_clk),
    .D(_0407_),
    .Q(\RAM[101][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2394_ (.CLK(clknet_leaf_37_clk),
    .D(_0408_),
    .Q(\RAM[102][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2395_ (.CLK(clknet_leaf_35_clk),
    .D(_0409_),
    .Q(\RAM[102][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2396_ (.CLK(clknet_leaf_36_clk),
    .D(_0410_),
    .Q(\RAM[102][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2397_ (.CLK(clknet_leaf_35_clk),
    .D(_0411_),
    .Q(\RAM[102][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2398_ (.CLK(clknet_leaf_36_clk),
    .D(_0412_),
    .Q(\RAM[103][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2399_ (.CLK(clknet_leaf_35_clk),
    .D(_0413_),
    .Q(\RAM[103][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2400_ (.CLK(clknet_leaf_36_clk),
    .D(_0414_),
    .Q(\RAM[103][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2401_ (.CLK(clknet_leaf_34_clk),
    .D(_0415_),
    .Q(\RAM[103][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2402_ (.CLK(clknet_leaf_29_clk),
    .D(_0416_),
    .Q(\RAM[104][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2403_ (.CLK(clknet_leaf_32_clk),
    .D(_0417_),
    .Q(\RAM[104][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2404_ (.CLK(clknet_leaf_31_clk),
    .D(_0418_),
    .Q(\RAM[104][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2405_ (.CLK(clknet_leaf_32_clk),
    .D(_0419_),
    .Q(\RAM[104][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2406_ (.CLK(clknet_leaf_29_clk),
    .D(_0420_),
    .Q(\RAM[105][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2407_ (.CLK(clknet_leaf_32_clk),
    .D(_0421_),
    .Q(\RAM[105][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2408_ (.CLK(clknet_leaf_31_clk),
    .D(_0422_),
    .Q(\RAM[105][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2409_ (.CLK(clknet_leaf_32_clk),
    .D(_0423_),
    .Q(\RAM[105][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2410_ (.CLK(clknet_leaf_29_clk),
    .D(_0424_),
    .Q(\RAM[106][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2411_ (.CLK(clknet_leaf_32_clk),
    .D(_0425_),
    .Q(\RAM[106][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2412_ (.CLK(clknet_leaf_31_clk),
    .D(_0426_),
    .Q(\RAM[106][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2413_ (.CLK(clknet_leaf_32_clk),
    .D(_0427_),
    .Q(\RAM[106][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2414_ (.CLK(clknet_leaf_29_clk),
    .D(_0428_),
    .Q(\RAM[107][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2415_ (.CLK(clknet_leaf_31_clk),
    .D(_0429_),
    .Q(\RAM[107][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2416_ (.CLK(clknet_leaf_31_clk),
    .D(_0430_),
    .Q(\RAM[107][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2417_ (.CLK(clknet_leaf_34_clk),
    .D(_0431_),
    .Q(\RAM[107][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2418_ (.CLK(clknet_leaf_34_clk),
    .D(_0432_),
    .Q(\RAM[108][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2419_ (.CLK(clknet_leaf_33_clk),
    .D(_0433_),
    .Q(\RAM[108][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2420_ (.CLK(clknet_leaf_33_clk),
    .D(_0434_),
    .Q(\RAM[108][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2421_ (.CLK(clknet_leaf_33_clk),
    .D(_0435_),
    .Q(\RAM[108][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2422_ (.CLK(clknet_leaf_17_clk),
    .D(_0436_),
    .Q(\RAM[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2423_ (.CLK(clknet_leaf_17_clk),
    .D(_0437_),
    .Q(\RAM[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2424_ (.CLK(clknet_leaf_18_clk),
    .D(_0438_),
    .Q(\RAM[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2425_ (.CLK(clknet_leaf_18_clk),
    .D(_0439_),
    .Q(\RAM[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2426_ (.CLK(clknet_leaf_34_clk),
    .D(_0440_),
    .Q(\RAM[110][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2427_ (.CLK(clknet_leaf_34_clk),
    .D(_0441_),
    .Q(\RAM[110][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2428_ (.CLK(clknet_leaf_32_clk),
    .D(_0442_),
    .Q(\RAM[110][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2429_ (.CLK(clknet_leaf_34_clk),
    .D(_0443_),
    .Q(\RAM[110][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2430_ (.CLK(clknet_leaf_34_clk),
    .D(_0444_),
    .Q(\RAM[111][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2431_ (.CLK(clknet_leaf_34_clk),
    .D(_0445_),
    .Q(\RAM[111][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2432_ (.CLK(clknet_leaf_32_clk),
    .D(_0446_),
    .Q(\RAM[111][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2433_ (.CLK(clknet_leaf_34_clk),
    .D(_0447_),
    .Q(\RAM[111][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2434_ (.CLK(clknet_leaf_38_clk),
    .D(_0448_),
    .Q(\RAM[112][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2435_ (.CLK(clknet_leaf_36_clk),
    .D(_0449_),
    .Q(\RAM[112][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2436_ (.CLK(clknet_leaf_36_clk),
    .D(_0450_),
    .Q(\RAM[112][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2437_ (.CLK(clknet_leaf_37_clk),
    .D(_0451_),
    .Q(\RAM[112][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2438_ (.CLK(clknet_leaf_38_clk),
    .D(_0452_),
    .Q(\RAM[113][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2439_ (.CLK(clknet_leaf_40_clk),
    .D(_0453_),
    .Q(\RAM[113][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2440_ (.CLK(clknet_leaf_40_clk),
    .D(_0454_),
    .Q(\RAM[113][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2441_ (.CLK(clknet_leaf_39_clk),
    .D(_0455_),
    .Q(\RAM[113][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2442_ (.CLK(clknet_leaf_38_clk),
    .D(_0456_),
    .Q(\RAM[114][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2443_ (.CLK(clknet_leaf_40_clk),
    .D(_0457_),
    .Q(\RAM[114][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2444_ (.CLK(clknet_leaf_40_clk),
    .D(_0458_),
    .Q(\RAM[114][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2445_ (.CLK(clknet_leaf_39_clk),
    .D(_0459_),
    .Q(\RAM[114][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2446_ (.CLK(clknet_leaf_39_clk),
    .D(_0460_),
    .Q(\RAM[115][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2447_ (.CLK(clknet_leaf_40_clk),
    .D(_0461_),
    .Q(\RAM[115][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2448_ (.CLK(clknet_leaf_40_clk),
    .D(_0462_),
    .Q(\RAM[115][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2449_ (.CLK(clknet_leaf_39_clk),
    .D(_0463_),
    .Q(\RAM[115][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2450_ (.CLK(clknet_leaf_28_clk),
    .D(_0464_),
    .Q(\RAM[116][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2451_ (.CLK(clknet_leaf_28_clk),
    .D(_0465_),
    .Q(\RAM[116][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2452_ (.CLK(clknet_leaf_28_clk),
    .D(_0466_),
    .Q(\RAM[116][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2453_ (.CLK(clknet_leaf_28_clk),
    .D(_0467_),
    .Q(\RAM[116][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2454_ (.CLK(clknet_leaf_28_clk),
    .D(_0468_),
    .Q(\RAM[117][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2455_ (.CLK(clknet_leaf_28_clk),
    .D(_0469_),
    .Q(\RAM[117][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2456_ (.CLK(clknet_leaf_38_clk),
    .D(_0470_),
    .Q(\RAM[117][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2457_ (.CLK(clknet_leaf_16_clk),
    .D(_0471_),
    .Q(\RAM[117][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2458_ (.CLK(clknet_leaf_4_clk),
    .D(_0472_),
    .Q(\RAM[118][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2459_ (.CLK(clknet_leaf_4_clk),
    .D(_0473_),
    .Q(\RAM[118][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2460_ (.CLK(clknet_leaf_4_clk),
    .D(_0474_),
    .Q(\RAM[118][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2461_ (.CLK(clknet_leaf_4_clk),
    .D(_0475_),
    .Q(\RAM[118][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2462_ (.CLK(clknet_leaf_18_clk),
    .D(_0476_),
    .Q(\RAM[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2463_ (.CLK(clknet_leaf_17_clk),
    .D(_0477_),
    .Q(\RAM[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2464_ (.CLK(clknet_leaf_18_clk),
    .D(_0478_),
    .Q(\RAM[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2465_ (.CLK(clknet_leaf_18_clk),
    .D(_0479_),
    .Q(\RAM[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2466_ (.CLK(clknet_leaf_38_clk),
    .D(_0480_),
    .Q(\RAM[120][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2467_ (.CLK(clknet_leaf_37_clk),
    .D(_0481_),
    .Q(\RAM[120][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2468_ (.CLK(clknet_leaf_28_clk),
    .D(_0482_),
    .Q(\RAM[120][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2469_ (.CLK(clknet_leaf_29_clk),
    .D(_0483_),
    .Q(\RAM[120][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2470_ (.CLK(clknet_leaf_28_clk),
    .D(_0484_),
    .Q(\RAM[121][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2471_ (.CLK(clknet_leaf_37_clk),
    .D(_0485_),
    .Q(\RAM[121][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2472_ (.CLK(clknet_leaf_29_clk),
    .D(_0486_),
    .Q(\RAM[121][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2473_ (.CLK(clknet_leaf_29_clk),
    .D(_0487_),
    .Q(\RAM[121][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2474_ (.CLK(clknet_leaf_38_clk),
    .D(_0488_),
    .Q(\RAM[122][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2475_ (.CLK(clknet_leaf_38_clk),
    .D(_0489_),
    .Q(\RAM[122][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2476_ (.CLK(clknet_leaf_28_clk),
    .D(_0490_),
    .Q(\RAM[122][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2477_ (.CLK(clknet_leaf_37_clk),
    .D(_0491_),
    .Q(\RAM[122][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2478_ (.CLK(clknet_leaf_38_clk),
    .D(_0492_),
    .Q(\RAM[123][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2479_ (.CLK(clknet_leaf_38_clk),
    .D(_0493_),
    .Q(\RAM[123][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2480_ (.CLK(clknet_leaf_28_clk),
    .D(_0494_),
    .Q(\RAM[123][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2481_ (.CLK(clknet_leaf_29_clk),
    .D(_0495_),
    .Q(\RAM[123][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2482_ (.CLK(clknet_leaf_36_clk),
    .D(_0496_),
    .Q(\RAM[124][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2483_ (.CLK(clknet_leaf_35_clk),
    .D(_0497_),
    .Q(\RAM[124][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2484_ (.CLK(clknet_leaf_35_clk),
    .D(_0498_),
    .Q(\RAM[124][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2485_ (.CLK(clknet_leaf_35_clk),
    .D(_0499_),
    .Q(\RAM[124][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2486_ (.CLK(clknet_leaf_41_clk),
    .D(_0500_),
    .Q(\RAM[125][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2487_ (.CLK(clknet_leaf_41_clk),
    .D(_0501_),
    .Q(\RAM[125][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2488_ (.CLK(clknet_leaf_41_clk),
    .D(_0502_),
    .Q(\RAM[125][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2489_ (.CLK(clknet_leaf_41_clk),
    .D(_0503_),
    .Q(\RAM[125][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2490_ (.CLK(clknet_leaf_41_clk),
    .D(_0504_),
    .Q(\RAM[126][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2491_ (.CLK(clknet_leaf_41_clk),
    .D(_0505_),
    .Q(\RAM[126][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2492_ (.CLK(clknet_leaf_41_clk),
    .D(_0506_),
    .Q(\RAM[126][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2493_ (.CLK(clknet_leaf_41_clk),
    .D(_0507_),
    .Q(\RAM[126][3] ));
 sky130_fd_sc_hd__dfxtp_1 _2494_ (.CLK(clknet_leaf_17_clk),
    .D(_0508_),
    .Q(\RAM[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _2495_ (.CLK(clknet_leaf_17_clk),
    .D(_0509_),
    .Q(\RAM[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _2496_ (.CLK(clknet_leaf_21_clk),
    .D(_0510_),
    .Q(\RAM[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _2497_ (.CLK(clknet_leaf_18_clk),
    .D(_0511_),
    .Q(\RAM[9][3] ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__buf_4 fanout100 (.A(net110),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_4 fanout101 (.A(net109),
    .X(net101));
 sky130_fd_sc_hd__buf_2 fanout102 (.A(net109),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_4 fanout103 (.A(net109),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_4 fanout104 (.A(net109),
    .X(net104));
 sky130_fd_sc_hd__buf_4 fanout105 (.A(net108),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_4 fanout106 (.A(net107),
    .X(net106));
 sky130_fd_sc_hd__buf_4 fanout107 (.A(net108),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_4 fanout108 (.A(net109),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_4 fanout109 (.A(net110),
    .X(net109));
 sky130_fd_sc_hd__buf_4 fanout110 (.A(net11),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_4 fanout111 (.A(net112),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_4 fanout112 (.A(net127),
    .X(net112));
 sky130_fd_sc_hd__buf_4 fanout113 (.A(net114),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_4 fanout114 (.A(net127),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_4 fanout115 (.A(net116),
    .X(net115));
 sky130_fd_sc_hd__buf_4 fanout116 (.A(net118),
    .X(net116));
 sky130_fd_sc_hd__buf_4 fanout117 (.A(net118),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_4 fanout118 (.A(net127),
    .X(net118));
 sky130_fd_sc_hd__buf_4 fanout119 (.A(net122),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_2 fanout120 (.A(net122),
    .X(net120));
 sky130_fd_sc_hd__buf_4 fanout121 (.A(net122),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_4 fanout122 (.A(net127),
    .X(net122));
 sky130_fd_sc_hd__buf_4 fanout123 (.A(net126),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_4 fanout124 (.A(net125),
    .X(net124));
 sky130_fd_sc_hd__buf_4 fanout125 (.A(net126),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_4 fanout126 (.A(net127),
    .X(net126));
 sky130_fd_sc_hd__buf_4 fanout127 (.A(net10),
    .X(net127));
 sky130_fd_sc_hd__buf_8 fanout128 (.A(net132),
    .X(net128));
 sky130_fd_sc_hd__buf_6 fanout129 (.A(net132),
    .X(net129));
 sky130_fd_sc_hd__buf_12 fanout130 (.A(net132),
    .X(net130));
 sky130_fd_sc_hd__buf_8 fanout131 (.A(net132),
    .X(net131));
 sky130_fd_sc_hd__buf_6 fanout132 (.A(net137),
    .X(net132));
 sky130_fd_sc_hd__buf_8 fanout133 (.A(net137),
    .X(net133));
 sky130_fd_sc_hd__buf_4 fanout134 (.A(net137),
    .X(net134));
 sky130_fd_sc_hd__buf_6 fanout135 (.A(net136),
    .X(net135));
 sky130_fd_sc_hd__buf_6 fanout136 (.A(net137),
    .X(net136));
 sky130_fd_sc_hd__buf_6 fanout137 (.A(net148),
    .X(net137));
 sky130_fd_sc_hd__buf_8 fanout138 (.A(net148),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_4 fanout139 (.A(net148),
    .X(net139));
 sky130_fd_sc_hd__buf_8 fanout140 (.A(net141),
    .X(net140));
 sky130_fd_sc_hd__buf_6 fanout141 (.A(net148),
    .X(net141));
 sky130_fd_sc_hd__buf_6 fanout142 (.A(net147),
    .X(net142));
 sky130_fd_sc_hd__buf_6 fanout143 (.A(net147),
    .X(net143));
 sky130_fd_sc_hd__buf_6 fanout144 (.A(net147),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_4 fanout145 (.A(net146),
    .X(net145));
 sky130_fd_sc_hd__buf_8 fanout146 (.A(net147),
    .X(net146));
 sky130_fd_sc_hd__buf_6 fanout147 (.A(net148),
    .X(net147));
 sky130_fd_sc_hd__buf_6 fanout148 (.A(net1),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_16 fanout17 (.A(_0867_),
    .X(net17));
 sky130_fd_sc_hd__buf_12 fanout18 (.A(_0851_),
    .X(net18));
 sky130_fd_sc_hd__buf_12 fanout19 (.A(_0846_),
    .X(net19));
 sky130_fd_sc_hd__buf_12 fanout20 (.A(_0830_),
    .X(net20));
 sky130_fd_sc_hd__buf_6 fanout21 (.A(_0561_),
    .X(net21));
 sky130_fd_sc_hd__buf_8 fanout22 (.A(_0545_),
    .X(net22));
 sky130_fd_sc_hd__buf_8 fanout23 (.A(_0544_),
    .X(net23));
 sky130_fd_sc_hd__buf_6 fanout24 (.A(_0542_),
    .X(net24));
 sky130_fd_sc_hd__buf_6 fanout25 (.A(_0539_),
    .X(net25));
 sky130_fd_sc_hd__buf_6 fanout26 (.A(_0538_),
    .X(net26));
 sky130_fd_sc_hd__buf_2 fanout27 (.A(_0538_),
    .X(net27));
 sky130_fd_sc_hd__buf_6 fanout28 (.A(_0533_),
    .X(net28));
 sky130_fd_sc_hd__buf_8 fanout29 (.A(_0532_),
    .X(net29));
 sky130_fd_sc_hd__buf_2 fanout30 (.A(_0532_),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_8 fanout31 (.A(net32),
    .X(net31));
 sky130_fd_sc_hd__buf_4 fanout32 (.A(net33),
    .X(net32));
 sky130_fd_sc_hd__buf_8 fanout33 (.A(_0514_),
    .X(net33));
 sky130_fd_sc_hd__buf_4 fanout34 (.A(_0513_),
    .X(net34));
 sky130_fd_sc_hd__buf_8 fanout35 (.A(_0513_),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_4 fanout36 (.A(net37),
    .X(net36));
 sky130_fd_sc_hd__buf_4 fanout37 (.A(net39),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_4 fanout38 (.A(net39),
    .X(net38));
 sky130_fd_sc_hd__buf_4 fanout39 (.A(net44),
    .X(net39));
 sky130_fd_sc_hd__buf_4 fanout40 (.A(net44),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_4 fanout41 (.A(net44),
    .X(net41));
 sky130_fd_sc_hd__buf_4 fanout42 (.A(net44),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_2 fanout43 (.A(net44),
    .X(net43));
 sky130_fd_sc_hd__buf_4 fanout44 (.A(net9),
    .X(net44));
 sky130_fd_sc_hd__buf_4 fanout45 (.A(net48),
    .X(net45));
 sky130_fd_sc_hd__buf_4 fanout46 (.A(net48),
    .X(net46));
 sky130_fd_sc_hd__buf_2 fanout47 (.A(net48),
    .X(net47));
 sky130_fd_sc_hd__buf_4 fanout48 (.A(net9),
    .X(net48));
 sky130_fd_sc_hd__buf_4 fanout49 (.A(net52),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_4 fanout50 (.A(net52),
    .X(net50));
 sky130_fd_sc_hd__buf_4 fanout51 (.A(net52),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_4 fanout52 (.A(net9),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_4 fanout53 (.A(net54),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_4 fanout54 (.A(net8),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_4 fanout55 (.A(net56),
    .X(net55));
 sky130_fd_sc_hd__buf_4 fanout56 (.A(net8),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_4 fanout57 (.A(net59),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_4 fanout58 (.A(net59),
    .X(net58));
 sky130_fd_sc_hd__buf_4 fanout59 (.A(net8),
    .X(net59));
 sky130_fd_sc_hd__buf_4 fanout60 (.A(net68),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_2 fanout61 (.A(net68),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_4 fanout62 (.A(net68),
    .X(net62));
 sky130_fd_sc_hd__buf_2 fanout63 (.A(net68),
    .X(net63));
 sky130_fd_sc_hd__buf_4 fanout64 (.A(net67),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_2 fanout65 (.A(net67),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_4 fanout66 (.A(net67),
    .X(net66));
 sky130_fd_sc_hd__buf_4 fanout67 (.A(net68),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_4 fanout68 (.A(net8),
    .X(net68));
 sky130_fd_sc_hd__buf_8 fanout69 (.A(net5),
    .X(net69));
 sky130_fd_sc_hd__buf_8 fanout70 (.A(net4),
    .X(net70));
 sky130_fd_sc_hd__buf_4 fanout71 (.A(net72),
    .X(net71));
 sky130_fd_sc_hd__buf_6 fanout72 (.A(net4),
    .X(net72));
 sky130_fd_sc_hd__buf_8 fanout73 (.A(net76),
    .X(net73));
 sky130_fd_sc_hd__buf_4 fanout74 (.A(net75),
    .X(net74));
 sky130_fd_sc_hd__buf_6 fanout75 (.A(net76),
    .X(net75));
 sky130_fd_sc_hd__buf_6 fanout76 (.A(net3),
    .X(net76));
 sky130_fd_sc_hd__buf_6 fanout77 (.A(net85),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_4 fanout78 (.A(net85),
    .X(net78));
 sky130_fd_sc_hd__buf_8 fanout79 (.A(net85),
    .X(net79));
 sky130_fd_sc_hd__buf_4 fanout80 (.A(net85),
    .X(net80));
 sky130_fd_sc_hd__buf_6 fanout81 (.A(net85),
    .X(net81));
 sky130_fd_sc_hd__buf_4 fanout82 (.A(net85),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_8 fanout83 (.A(net85),
    .X(net83));
 sky130_fd_sc_hd__buf_4 fanout84 (.A(net85),
    .X(net84));
 sky130_fd_sc_hd__buf_8 fanout85 (.A(net2),
    .X(net85));
 sky130_fd_sc_hd__buf_6 fanout86 (.A(net89),
    .X(net86));
 sky130_fd_sc_hd__buf_6 fanout87 (.A(net89),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_4 fanout88 (.A(net89),
    .X(net88));
 sky130_fd_sc_hd__buf_4 fanout89 (.A(net94),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_8 fanout90 (.A(net94),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_4 fanout91 (.A(net94),
    .X(net91));
 sky130_fd_sc_hd__buf_6 fanout92 (.A(net94),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_4 fanout93 (.A(net94),
    .X(net93));
 sky130_fd_sc_hd__buf_4 fanout94 (.A(net2),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_4 fanout95 (.A(net97),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_4 fanout96 (.A(net97),
    .X(net96));
 sky130_fd_sc_hd__buf_4 fanout97 (.A(net110),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_4 fanout98 (.A(net100),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_4 fanout99 (.A(net100),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(ram_addr[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(w_val[2]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(w_val[3]),
    .X(net11));
 sky130_fd_sc_hd__buf_4 input12 (.A(wen),
    .X(net12));
 sky130_fd_sc_hd__buf_2 input2 (.A(ram_addr[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(ram_addr[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_8 input4 (.A(ram_addr[3]),
    .X(net4));
 sky130_fd_sc_hd__buf_2 input5 (.A(ram_addr[4]),
    .X(net5));
 sky130_fd_sc_hd__buf_8 input6 (.A(ram_addr[5]),
    .X(net6));
 sky130_fd_sc_hd__buf_6 input7 (.A(ram_addr[6]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_4 input8 (.A(w_val[0]),
    .X(net8));
 sky130_fd_sc_hd__buf_2 input9 (.A(w_val[1]),
    .X(net9));
 sky130_fd_sc_hd__buf_4 output13 (.A(net13),
    .X(r_val[0]));
 sky130_fd_sc_hd__buf_4 output14 (.A(net14),
    .X(r_val[1]));
 sky130_fd_sc_hd__buf_4 output15 (.A(net15),
    .X(r_val[2]));
 sky130_fd_sc_hd__buf_4 output16 (.A(net16),
    .X(r_val[3]));
endmodule

