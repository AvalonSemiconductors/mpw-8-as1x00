VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_tms1x00
  CLASS BLOCK ;
  FOREIGN wrapped_tms1x00 ;
  ORIGIN 0.000 0.000 ;
  SIZE 750.000 BY 700.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.670 696.000 10.950 700.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.870 696.000 204.150 700.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.190 696.000 223.470 700.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.510 696.000 242.790 700.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.830 696.000 262.110 700.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.150 696.000 281.430 700.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.470 696.000 300.750 700.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.790 696.000 320.070 700.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.110 696.000 339.390 700.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.430 696.000 358.710 700.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.750 696.000 378.030 700.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 696.000 30.270 700.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.070 696.000 397.350 700.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.390 696.000 416.670 700.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.710 696.000 435.990 700.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.030 696.000 455.310 700.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.350 696.000 474.630 700.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.670 696.000 493.950 700.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.990 696.000 513.270 700.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.310 696.000 532.590 700.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.630 696.000 551.910 700.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.950 696.000 571.230 700.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 696.000 49.590 700.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 590.270 696.000 590.550 700.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.590 696.000 609.870 700.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.910 696.000 629.190 700.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 648.230 696.000 648.510 700.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.550 696.000 667.830 700.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.870 696.000 687.150 700.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.190 696.000 706.470 700.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.510 696.000 725.790 700.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 696.000 68.910 700.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 696.000 88.230 700.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.270 696.000 107.550 700.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 696.000 126.870 700.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.910 696.000 146.190 700.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.230 696.000 165.510 700.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.550 696.000 184.830 700.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 696.000 17.390 700.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.310 696.000 210.590 700.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 696.000 229.910 700.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.950 696.000 249.230 700.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.270 696.000 268.550 700.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.590 696.000 287.870 700.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.910 696.000 307.190 700.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.230 696.000 326.510 700.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.550 696.000 345.830 700.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.870 696.000 365.150 700.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.190 696.000 384.470 700.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 696.000 36.710 700.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.510 696.000 403.790 700.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.830 696.000 423.110 700.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.150 696.000 442.430 700.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.470 696.000 461.750 700.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.790 696.000 481.070 700.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.110 696.000 500.390 700.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.430 696.000 519.710 700.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.750 696.000 539.030 700.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.070 696.000 558.350 700.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.390 696.000 577.670 700.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 696.000 56.030 700.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 596.710 696.000 596.990 700.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.030 696.000 616.310 700.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 635.350 696.000 635.630 700.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 654.670 696.000 654.950 700.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.990 696.000 674.270 700.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 693.310 696.000 693.590 700.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.630 696.000 712.910 700.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.950 696.000 732.230 700.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 696.000 75.350 700.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 696.000 94.670 700.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.710 696.000 113.990 700.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.030 696.000 133.310 700.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.350 696.000 152.630 700.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.670 696.000 171.950 700.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 696.000 191.270 700.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 696.000 23.830 700.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.750 696.000 217.030 700.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.070 696.000 236.350 700.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 696.000 255.670 700.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 696.000 274.990 700.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.030 696.000 294.310 700.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.350 696.000 313.630 700.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.670 696.000 332.950 700.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.990 696.000 352.270 700.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.310 696.000 371.590 700.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.630 696.000 390.910 700.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 696.000 43.150 700.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.950 696.000 410.230 700.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.270 696.000 429.550 700.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.590 696.000 448.870 700.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.910 696.000 468.190 700.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.230 696.000 487.510 700.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.550 696.000 506.830 700.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.870 696.000 526.150 700.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.190 696.000 545.470 700.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.510 696.000 564.790 700.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.830 696.000 584.110 700.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 696.000 62.470 700.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.150 696.000 603.430 700.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.470 696.000 622.750 700.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.790 696.000 642.070 700.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.110 696.000 661.390 700.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.430 696.000 680.710 700.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.750 696.000 700.030 700.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.070 696.000 719.350 700.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 738.390 696.000 738.670 700.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 696.000 81.790 700.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.830 696.000 101.110 700.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 696.000 120.430 700.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.470 696.000 139.750 700.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 696.000 159.070 700.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.110 696.000 178.390 700.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.430 696.000 197.710 700.000 ;
    END
  END io_out[9]
  PIN ram_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 66.680 750.000 67.280 ;
    END
  END ram_addr[0]
  PIN ram_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 197.240 750.000 197.840 ;
    END
  END ram_addr[1]
  PIN ram_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 327.800 750.000 328.400 ;
    END
  END ram_addr[2]
  PIN ram_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 458.360 750.000 458.960 ;
    END
  END ram_addr[3]
  PIN ram_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 588.920 750.000 589.520 ;
    END
  END ram_addr[4]
  PIN ram_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 632.440 750.000 633.040 ;
    END
  END ram_addr[5]
  PIN ram_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 675.960 750.000 676.560 ;
    END
  END ram_addr[6]
  PIN ram_val_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 110.200 750.000 110.800 ;
    END
  END ram_val_in[0]
  PIN ram_val_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 240.760 750.000 241.360 ;
    END
  END ram_val_in[1]
  PIN ram_val_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 371.320 750.000 371.920 ;
    END
  END ram_val_in[2]
  PIN ram_val_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 501.880 750.000 502.480 ;
    END
  END ram_val_in[3]
  PIN ram_val_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 153.720 750.000 154.320 ;
    END
  END ram_val_out[0]
  PIN ram_val_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 284.280 750.000 284.880 ;
    END
  END ram_val_out[1]
  PIN ram_val_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 414.840 750.000 415.440 ;
    END
  END ram_val_out[2]
  PIN ram_val_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 545.400 750.000 546.000 ;
    END
  END ram_val_out[3]
  PIN ram_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 23.160 750.000 23.760 ;
    END
  END ram_we
  PIN rom_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END rom_addr[0]
  PIN rom_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 4.000 64.560 ;
    END
  END rom_addr[1]
  PIN rom_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 4.000 97.200 ;
    END
  END rom_addr[2]
  PIN rom_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END rom_addr[3]
  PIN rom_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 4.000 162.480 ;
    END
  END rom_addr[4]
  PIN rom_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.520 4.000 195.120 ;
    END
  END rom_addr[5]
  PIN rom_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.160 4.000 227.760 ;
    END
  END rom_addr[6]
  PIN rom_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.800 4.000 260.400 ;
    END
  END rom_addr[7]
  PIN rom_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END rom_addr[8]
  PIN rom_csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 4.000 15.600 ;
    END
  END rom_csb
  PIN rom_value[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END rom_value[0]
  PIN rom_value[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 341.400 4.000 342.000 ;
    END
  END rom_value[10]
  PIN rom_value[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.720 4.000 358.320 ;
    END
  END rom_value[11]
  PIN rom_value[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END rom_value[12]
  PIN rom_value[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 390.360 4.000 390.960 ;
    END
  END rom_value[13]
  PIN rom_value[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 406.680 4.000 407.280 ;
    END
  END rom_value[14]
  PIN rom_value[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 423.000 4.000 423.600 ;
    END
  END rom_value[15]
  PIN rom_value[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 439.320 4.000 439.920 ;
    END
  END rom_value[16]
  PIN rom_value[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 455.640 4.000 456.240 ;
    END
  END rom_value[17]
  PIN rom_value[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 471.960 4.000 472.560 ;
    END
  END rom_value[18]
  PIN rom_value[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 488.280 4.000 488.880 ;
    END
  END rom_value[19]
  PIN rom_value[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 4.000 80.880 ;
    END
  END rom_value[1]
  PIN rom_value[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 504.600 4.000 505.200 ;
    END
  END rom_value[20]
  PIN rom_value[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.920 4.000 521.520 ;
    END
  END rom_value[21]
  PIN rom_value[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.240 4.000 537.840 ;
    END
  END rom_value[22]
  PIN rom_value[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 553.560 4.000 554.160 ;
    END
  END rom_value[23]
  PIN rom_value[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 569.880 4.000 570.480 ;
    END
  END rom_value[24]
  PIN rom_value[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 586.200 4.000 586.800 ;
    END
  END rom_value[25]
  PIN rom_value[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 602.520 4.000 603.120 ;
    END
  END rom_value[26]
  PIN rom_value[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 618.840 4.000 619.440 ;
    END
  END rom_value[27]
  PIN rom_value[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 635.160 4.000 635.760 ;
    END
  END rom_value[28]
  PIN rom_value[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 651.480 4.000 652.080 ;
    END
  END rom_value[29]
  PIN rom_value[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END rom_value[2]
  PIN rom_value[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 667.800 4.000 668.400 ;
    END
  END rom_value[30]
  PIN rom_value[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 684.120 4.000 684.720 ;
    END
  END rom_value[31]
  PIN rom_value[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END rom_value[3]
  PIN rom_value[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 4.000 178.800 ;
    END
  END rom_value[4]
  PIN rom_value[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END rom_value[5]
  PIN rom_value[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 243.480 4.000 244.080 ;
    END
  END rom_value[6]
  PIN rom_value[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.120 4.000 276.720 ;
    END
  END rom_value[7]
  PIN rom_value[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.760 4.000 309.360 ;
    END
  END rom_value[8]
  PIN rom_value[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.080 4.000 325.680 ;
    END
  END rom_value[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 688.400 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 688.400 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 0.000 10.490 4.000 ;
    END
  END wb_clk_i
  PIN wb_rom_adrb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 4.000 ;
    END
  END wb_rom_adrb[0]
  PIN wb_rom_adrb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 4.000 ;
    END
  END wb_rom_adrb[1]
  PIN wb_rom_adrb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 4.000 ;
    END
  END wb_rom_adrb[2]
  PIN wb_rom_adrb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 4.000 ;
    END
  END wb_rom_adrb[3]
  PIN wb_rom_adrb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END wb_rom_adrb[4]
  PIN wb_rom_adrb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 0.000 81.330 4.000 ;
    END
  END wb_rom_adrb[5]
  PIN wb_rom_adrb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 0.000 91.450 4.000 ;
    END
  END wb_rom_adrb[6]
  PIN wb_rom_adrb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 0.000 101.570 4.000 ;
    END
  END wb_rom_adrb[7]
  PIN wb_rom_adrb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.410 0.000 111.690 4.000 ;
    END
  END wb_rom_adrb[8]
  PIN wb_rom_csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 0.000 15.550 4.000 ;
    END
  END wb_rom_csb
  PIN wb_rom_val[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END wb_rom_val[0]
  PIN wb_rom_val[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 0.000 126.870 4.000 ;
    END
  END wb_rom_val[10]
  PIN wb_rom_val[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 0.000 131.930 4.000 ;
    END
  END wb_rom_val[11]
  PIN wb_rom_val[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 0.000 136.990 4.000 ;
    END
  END wb_rom_val[12]
  PIN wb_rom_val[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END wb_rom_val[13]
  PIN wb_rom_val[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 0.000 147.110 4.000 ;
    END
  END wb_rom_val[14]
  PIN wb_rom_val[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 0.000 152.170 4.000 ;
    END
  END wb_rom_val[15]
  PIN wb_rom_val[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.950 0.000 157.230 4.000 ;
    END
  END wb_rom_val[16]
  PIN wb_rom_val[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 0.000 162.290 4.000 ;
    END
  END wb_rom_val[17]
  PIN wb_rom_val[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.070 0.000 167.350 4.000 ;
    END
  END wb_rom_val[18]
  PIN wb_rom_val[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.130 0.000 172.410 4.000 ;
    END
  END wb_rom_val[19]
  PIN wb_rom_val[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 4.000 ;
    END
  END wb_rom_val[1]
  PIN wb_rom_val[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END wb_rom_val[20]
  PIN wb_rom_val[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 0.000 182.530 4.000 ;
    END
  END wb_rom_val[21]
  PIN wb_rom_val[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.310 0.000 187.590 4.000 ;
    END
  END wb_rom_val[22]
  PIN wb_rom_val[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 0.000 192.650 4.000 ;
    END
  END wb_rom_val[23]
  PIN wb_rom_val[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.430 0.000 197.710 4.000 ;
    END
  END wb_rom_val[24]
  PIN wb_rom_val[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.490 0.000 202.770 4.000 ;
    END
  END wb_rom_val[25]
  PIN wb_rom_val[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.550 0.000 207.830 4.000 ;
    END
  END wb_rom_val[26]
  PIN wb_rom_val[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END wb_rom_val[27]
  PIN wb_rom_val[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.670 0.000 217.950 4.000 ;
    END
  END wb_rom_val[28]
  PIN wb_rom_val[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.730 0.000 223.010 4.000 ;
    END
  END wb_rom_val[29]
  PIN wb_rom_val[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 4.000 ;
    END
  END wb_rom_val[2]
  PIN wb_rom_val[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.790 0.000 228.070 4.000 ;
    END
  END wb_rom_val[30]
  PIN wb_rom_val[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.850 0.000 233.130 4.000 ;
    END
  END wb_rom_val[31]
  PIN wb_rom_val[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 0.000 66.150 4.000 ;
    END
  END wb_rom_val[3]
  PIN wb_rom_val[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 4.000 ;
    END
  END wb_rom_val[4]
  PIN wb_rom_val[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 0.000 86.390 4.000 ;
    END
  END wb_rom_val[5]
  PIN wb_rom_val[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.230 0.000 96.510 4.000 ;
    END
  END wb_rom_val[6]
  PIN wb_rom_val[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END wb_rom_val[7]
  PIN wb_rom_val[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.470 0.000 116.750 4.000 ;
    END
  END wb_rom_val[8]
  PIN wb_rom_val[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530 0.000 121.810 4.000 ;
    END
  END wb_rom_val[9]
  PIN wb_rom_web
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 0.000 20.610 4.000 ;
    END
  END wb_rom_web
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 0.000 25.670 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.910 0.000 238.190 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.150 0.000 258.430 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.950 0.000 410.230 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 0.000 425.410 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.310 0.000 440.590 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.490 0.000 455.770 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.670 0.000 470.950 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.850 0.000 486.130 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.030 0.000 501.310 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.210 0.000 516.490 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 0.000 531.670 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.570 0.000 546.850 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.330 0.000 273.610 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.750 0.000 562.030 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.930 0.000 577.210 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.110 0.000 592.390 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 607.290 0.000 607.570 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.470 0.000 622.750 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.650 0.000 637.930 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.830 0.000 653.110 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.010 0.000 668.290 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 683.190 0.000 683.470 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.370 0.000 698.650 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 0.000 288.790 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.550 0.000 713.830 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.730 0.000 729.010 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.690 0.000 303.970 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 0.000 319.150 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.050 0.000 334.330 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.230 0.000 349.510 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.410 0.000 364.690 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.590 0.000 379.870 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.770 0.000 395.050 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 0.000 243.250 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.210 0.000 263.490 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.010 0.000 415.290 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.190 0.000 430.470 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.370 0.000 445.650 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 0.000 460.830 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.730 0.000 476.010 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.910 0.000 491.190 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.090 0.000 506.370 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.270 0.000 521.550 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.450 0.000 536.730 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.630 0.000 551.910 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.390 0.000 278.670 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.810 0.000 567.090 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.990 0.000 582.270 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.170 0.000 597.450 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.350 0.000 612.630 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.530 0.000 627.810 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 642.710 0.000 642.990 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.890 0.000 658.170 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.070 0.000 673.350 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.250 0.000 688.530 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.430 0.000 703.710 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 0.000 293.850 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.610 0.000 718.890 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.790 0.000 734.070 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.750 0.000 309.030 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.930 0.000 324.210 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.110 0.000 339.390 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 0.000 354.570 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.470 0.000 369.750 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.650 0.000 384.930 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.830 0.000 400.110 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.270 0.000 268.550 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.070 0.000 420.350 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.250 0.000 435.530 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.430 0.000 450.710 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.610 0.000 465.890 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.790 0.000 481.070 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.970 0.000 496.250 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.150 0.000 511.430 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.330 0.000 526.610 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.510 0.000 541.790 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.690 0.000 556.970 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.870 0.000 572.150 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.050 0.000 587.330 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.230 0.000 602.510 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.410 0.000 617.690 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.590 0.000 632.870 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.770 0.000 648.050 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.950 0.000 663.230 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 678.130 0.000 678.410 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 693.310 0.000 693.590 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.490 0.000 708.770 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.630 0.000 298.910 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.670 0.000 723.950 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 738.850 0.000 739.130 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.810 0.000 314.090 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.990 0.000 329.270 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.170 0.000 344.450 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.350 0.000 359.630 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.530 0.000 374.810 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 0.000 389.990 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.890 0.000 405.170 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 0.000 248.310 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.090 0.000 253.370 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 744.280 688.245 ;
      LAYER met1 ;
        RECT 2.830 0.040 744.280 688.400 ;
      LAYER met2 ;
        RECT 2.390 695.720 10.390 696.730 ;
        RECT 11.230 695.720 16.830 696.730 ;
        RECT 17.670 695.720 23.270 696.730 ;
        RECT 24.110 695.720 29.710 696.730 ;
        RECT 30.550 695.720 36.150 696.730 ;
        RECT 36.990 695.720 42.590 696.730 ;
        RECT 43.430 695.720 49.030 696.730 ;
        RECT 49.870 695.720 55.470 696.730 ;
        RECT 56.310 695.720 61.910 696.730 ;
        RECT 62.750 695.720 68.350 696.730 ;
        RECT 69.190 695.720 74.790 696.730 ;
        RECT 75.630 695.720 81.230 696.730 ;
        RECT 82.070 695.720 87.670 696.730 ;
        RECT 88.510 695.720 94.110 696.730 ;
        RECT 94.950 695.720 100.550 696.730 ;
        RECT 101.390 695.720 106.990 696.730 ;
        RECT 107.830 695.720 113.430 696.730 ;
        RECT 114.270 695.720 119.870 696.730 ;
        RECT 120.710 695.720 126.310 696.730 ;
        RECT 127.150 695.720 132.750 696.730 ;
        RECT 133.590 695.720 139.190 696.730 ;
        RECT 140.030 695.720 145.630 696.730 ;
        RECT 146.470 695.720 152.070 696.730 ;
        RECT 152.910 695.720 158.510 696.730 ;
        RECT 159.350 695.720 164.950 696.730 ;
        RECT 165.790 695.720 171.390 696.730 ;
        RECT 172.230 695.720 177.830 696.730 ;
        RECT 178.670 695.720 184.270 696.730 ;
        RECT 185.110 695.720 190.710 696.730 ;
        RECT 191.550 695.720 197.150 696.730 ;
        RECT 197.990 695.720 203.590 696.730 ;
        RECT 204.430 695.720 210.030 696.730 ;
        RECT 210.870 695.720 216.470 696.730 ;
        RECT 217.310 695.720 222.910 696.730 ;
        RECT 223.750 695.720 229.350 696.730 ;
        RECT 230.190 695.720 235.790 696.730 ;
        RECT 236.630 695.720 242.230 696.730 ;
        RECT 243.070 695.720 248.670 696.730 ;
        RECT 249.510 695.720 255.110 696.730 ;
        RECT 255.950 695.720 261.550 696.730 ;
        RECT 262.390 695.720 267.990 696.730 ;
        RECT 268.830 695.720 274.430 696.730 ;
        RECT 275.270 695.720 280.870 696.730 ;
        RECT 281.710 695.720 287.310 696.730 ;
        RECT 288.150 695.720 293.750 696.730 ;
        RECT 294.590 695.720 300.190 696.730 ;
        RECT 301.030 695.720 306.630 696.730 ;
        RECT 307.470 695.720 313.070 696.730 ;
        RECT 313.910 695.720 319.510 696.730 ;
        RECT 320.350 695.720 325.950 696.730 ;
        RECT 326.790 695.720 332.390 696.730 ;
        RECT 333.230 695.720 338.830 696.730 ;
        RECT 339.670 695.720 345.270 696.730 ;
        RECT 346.110 695.720 351.710 696.730 ;
        RECT 352.550 695.720 358.150 696.730 ;
        RECT 358.990 695.720 364.590 696.730 ;
        RECT 365.430 695.720 371.030 696.730 ;
        RECT 371.870 695.720 377.470 696.730 ;
        RECT 378.310 695.720 383.910 696.730 ;
        RECT 384.750 695.720 390.350 696.730 ;
        RECT 391.190 695.720 396.790 696.730 ;
        RECT 397.630 695.720 403.230 696.730 ;
        RECT 404.070 695.720 409.670 696.730 ;
        RECT 410.510 695.720 416.110 696.730 ;
        RECT 416.950 695.720 422.550 696.730 ;
        RECT 423.390 695.720 428.990 696.730 ;
        RECT 429.830 695.720 435.430 696.730 ;
        RECT 436.270 695.720 441.870 696.730 ;
        RECT 442.710 695.720 448.310 696.730 ;
        RECT 449.150 695.720 454.750 696.730 ;
        RECT 455.590 695.720 461.190 696.730 ;
        RECT 462.030 695.720 467.630 696.730 ;
        RECT 468.470 695.720 474.070 696.730 ;
        RECT 474.910 695.720 480.510 696.730 ;
        RECT 481.350 695.720 486.950 696.730 ;
        RECT 487.790 695.720 493.390 696.730 ;
        RECT 494.230 695.720 499.830 696.730 ;
        RECT 500.670 695.720 506.270 696.730 ;
        RECT 507.110 695.720 512.710 696.730 ;
        RECT 513.550 695.720 519.150 696.730 ;
        RECT 519.990 695.720 525.590 696.730 ;
        RECT 526.430 695.720 532.030 696.730 ;
        RECT 532.870 695.720 538.470 696.730 ;
        RECT 539.310 695.720 544.910 696.730 ;
        RECT 545.750 695.720 551.350 696.730 ;
        RECT 552.190 695.720 557.790 696.730 ;
        RECT 558.630 695.720 564.230 696.730 ;
        RECT 565.070 695.720 570.670 696.730 ;
        RECT 571.510 695.720 577.110 696.730 ;
        RECT 577.950 695.720 583.550 696.730 ;
        RECT 584.390 695.720 589.990 696.730 ;
        RECT 590.830 695.720 596.430 696.730 ;
        RECT 597.270 695.720 602.870 696.730 ;
        RECT 603.710 695.720 609.310 696.730 ;
        RECT 610.150 695.720 615.750 696.730 ;
        RECT 616.590 695.720 622.190 696.730 ;
        RECT 623.030 695.720 628.630 696.730 ;
        RECT 629.470 695.720 635.070 696.730 ;
        RECT 635.910 695.720 641.510 696.730 ;
        RECT 642.350 695.720 647.950 696.730 ;
        RECT 648.790 695.720 654.390 696.730 ;
        RECT 655.230 695.720 660.830 696.730 ;
        RECT 661.670 695.720 667.270 696.730 ;
        RECT 668.110 695.720 673.710 696.730 ;
        RECT 674.550 695.720 680.150 696.730 ;
        RECT 680.990 695.720 686.590 696.730 ;
        RECT 687.430 695.720 693.030 696.730 ;
        RECT 693.870 695.720 699.470 696.730 ;
        RECT 700.310 695.720 705.910 696.730 ;
        RECT 706.750 695.720 712.350 696.730 ;
        RECT 713.190 695.720 718.790 696.730 ;
        RECT 719.630 695.720 725.230 696.730 ;
        RECT 726.070 695.720 731.670 696.730 ;
        RECT 732.510 695.720 738.110 696.730 ;
        RECT 738.950 695.720 741.890 696.730 ;
        RECT 2.390 4.280 741.890 695.720 ;
        RECT 2.390 0.010 9.930 4.280 ;
        RECT 10.770 0.010 14.990 4.280 ;
        RECT 15.830 0.010 20.050 4.280 ;
        RECT 20.890 0.010 25.110 4.280 ;
        RECT 25.950 0.010 30.170 4.280 ;
        RECT 31.010 0.010 35.230 4.280 ;
        RECT 36.070 0.010 40.290 4.280 ;
        RECT 41.130 0.010 45.350 4.280 ;
        RECT 46.190 0.010 50.410 4.280 ;
        RECT 51.250 0.010 55.470 4.280 ;
        RECT 56.310 0.010 60.530 4.280 ;
        RECT 61.370 0.010 65.590 4.280 ;
        RECT 66.430 0.010 70.650 4.280 ;
        RECT 71.490 0.010 75.710 4.280 ;
        RECT 76.550 0.010 80.770 4.280 ;
        RECT 81.610 0.010 85.830 4.280 ;
        RECT 86.670 0.010 90.890 4.280 ;
        RECT 91.730 0.010 95.950 4.280 ;
        RECT 96.790 0.010 101.010 4.280 ;
        RECT 101.850 0.010 106.070 4.280 ;
        RECT 106.910 0.010 111.130 4.280 ;
        RECT 111.970 0.010 116.190 4.280 ;
        RECT 117.030 0.010 121.250 4.280 ;
        RECT 122.090 0.010 126.310 4.280 ;
        RECT 127.150 0.010 131.370 4.280 ;
        RECT 132.210 0.010 136.430 4.280 ;
        RECT 137.270 0.010 141.490 4.280 ;
        RECT 142.330 0.010 146.550 4.280 ;
        RECT 147.390 0.010 151.610 4.280 ;
        RECT 152.450 0.010 156.670 4.280 ;
        RECT 157.510 0.010 161.730 4.280 ;
        RECT 162.570 0.010 166.790 4.280 ;
        RECT 167.630 0.010 171.850 4.280 ;
        RECT 172.690 0.010 176.910 4.280 ;
        RECT 177.750 0.010 181.970 4.280 ;
        RECT 182.810 0.010 187.030 4.280 ;
        RECT 187.870 0.010 192.090 4.280 ;
        RECT 192.930 0.010 197.150 4.280 ;
        RECT 197.990 0.010 202.210 4.280 ;
        RECT 203.050 0.010 207.270 4.280 ;
        RECT 208.110 0.010 212.330 4.280 ;
        RECT 213.170 0.010 217.390 4.280 ;
        RECT 218.230 0.010 222.450 4.280 ;
        RECT 223.290 0.010 227.510 4.280 ;
        RECT 228.350 0.010 232.570 4.280 ;
        RECT 233.410 0.010 237.630 4.280 ;
        RECT 238.470 0.010 242.690 4.280 ;
        RECT 243.530 0.010 247.750 4.280 ;
        RECT 248.590 0.010 252.810 4.280 ;
        RECT 253.650 0.010 257.870 4.280 ;
        RECT 258.710 0.010 262.930 4.280 ;
        RECT 263.770 0.010 267.990 4.280 ;
        RECT 268.830 0.010 273.050 4.280 ;
        RECT 273.890 0.010 278.110 4.280 ;
        RECT 278.950 0.010 283.170 4.280 ;
        RECT 284.010 0.010 288.230 4.280 ;
        RECT 289.070 0.010 293.290 4.280 ;
        RECT 294.130 0.010 298.350 4.280 ;
        RECT 299.190 0.010 303.410 4.280 ;
        RECT 304.250 0.010 308.470 4.280 ;
        RECT 309.310 0.010 313.530 4.280 ;
        RECT 314.370 0.010 318.590 4.280 ;
        RECT 319.430 0.010 323.650 4.280 ;
        RECT 324.490 0.010 328.710 4.280 ;
        RECT 329.550 0.010 333.770 4.280 ;
        RECT 334.610 0.010 338.830 4.280 ;
        RECT 339.670 0.010 343.890 4.280 ;
        RECT 344.730 0.010 348.950 4.280 ;
        RECT 349.790 0.010 354.010 4.280 ;
        RECT 354.850 0.010 359.070 4.280 ;
        RECT 359.910 0.010 364.130 4.280 ;
        RECT 364.970 0.010 369.190 4.280 ;
        RECT 370.030 0.010 374.250 4.280 ;
        RECT 375.090 0.010 379.310 4.280 ;
        RECT 380.150 0.010 384.370 4.280 ;
        RECT 385.210 0.010 389.430 4.280 ;
        RECT 390.270 0.010 394.490 4.280 ;
        RECT 395.330 0.010 399.550 4.280 ;
        RECT 400.390 0.010 404.610 4.280 ;
        RECT 405.450 0.010 409.670 4.280 ;
        RECT 410.510 0.010 414.730 4.280 ;
        RECT 415.570 0.010 419.790 4.280 ;
        RECT 420.630 0.010 424.850 4.280 ;
        RECT 425.690 0.010 429.910 4.280 ;
        RECT 430.750 0.010 434.970 4.280 ;
        RECT 435.810 0.010 440.030 4.280 ;
        RECT 440.870 0.010 445.090 4.280 ;
        RECT 445.930 0.010 450.150 4.280 ;
        RECT 450.990 0.010 455.210 4.280 ;
        RECT 456.050 0.010 460.270 4.280 ;
        RECT 461.110 0.010 465.330 4.280 ;
        RECT 466.170 0.010 470.390 4.280 ;
        RECT 471.230 0.010 475.450 4.280 ;
        RECT 476.290 0.010 480.510 4.280 ;
        RECT 481.350 0.010 485.570 4.280 ;
        RECT 486.410 0.010 490.630 4.280 ;
        RECT 491.470 0.010 495.690 4.280 ;
        RECT 496.530 0.010 500.750 4.280 ;
        RECT 501.590 0.010 505.810 4.280 ;
        RECT 506.650 0.010 510.870 4.280 ;
        RECT 511.710 0.010 515.930 4.280 ;
        RECT 516.770 0.010 520.990 4.280 ;
        RECT 521.830 0.010 526.050 4.280 ;
        RECT 526.890 0.010 531.110 4.280 ;
        RECT 531.950 0.010 536.170 4.280 ;
        RECT 537.010 0.010 541.230 4.280 ;
        RECT 542.070 0.010 546.290 4.280 ;
        RECT 547.130 0.010 551.350 4.280 ;
        RECT 552.190 0.010 556.410 4.280 ;
        RECT 557.250 0.010 561.470 4.280 ;
        RECT 562.310 0.010 566.530 4.280 ;
        RECT 567.370 0.010 571.590 4.280 ;
        RECT 572.430 0.010 576.650 4.280 ;
        RECT 577.490 0.010 581.710 4.280 ;
        RECT 582.550 0.010 586.770 4.280 ;
        RECT 587.610 0.010 591.830 4.280 ;
        RECT 592.670 0.010 596.890 4.280 ;
        RECT 597.730 0.010 601.950 4.280 ;
        RECT 602.790 0.010 607.010 4.280 ;
        RECT 607.850 0.010 612.070 4.280 ;
        RECT 612.910 0.010 617.130 4.280 ;
        RECT 617.970 0.010 622.190 4.280 ;
        RECT 623.030 0.010 627.250 4.280 ;
        RECT 628.090 0.010 632.310 4.280 ;
        RECT 633.150 0.010 637.370 4.280 ;
        RECT 638.210 0.010 642.430 4.280 ;
        RECT 643.270 0.010 647.490 4.280 ;
        RECT 648.330 0.010 652.550 4.280 ;
        RECT 653.390 0.010 657.610 4.280 ;
        RECT 658.450 0.010 662.670 4.280 ;
        RECT 663.510 0.010 667.730 4.280 ;
        RECT 668.570 0.010 672.790 4.280 ;
        RECT 673.630 0.010 677.850 4.280 ;
        RECT 678.690 0.010 682.910 4.280 ;
        RECT 683.750 0.010 687.970 4.280 ;
        RECT 688.810 0.010 693.030 4.280 ;
        RECT 693.870 0.010 698.090 4.280 ;
        RECT 698.930 0.010 703.150 4.280 ;
        RECT 703.990 0.010 708.210 4.280 ;
        RECT 709.050 0.010 713.270 4.280 ;
        RECT 714.110 0.010 718.330 4.280 ;
        RECT 719.170 0.010 723.390 4.280 ;
        RECT 724.230 0.010 728.450 4.280 ;
        RECT 729.290 0.010 733.510 4.280 ;
        RECT 734.350 0.010 738.570 4.280 ;
        RECT 739.410 0.010 741.890 4.280 ;
      LAYER met3 ;
        RECT 2.365 685.120 746.000 688.325 ;
        RECT 4.400 683.720 746.000 685.120 ;
        RECT 2.365 676.960 746.000 683.720 ;
        RECT 2.365 675.560 745.600 676.960 ;
        RECT 2.365 668.800 746.000 675.560 ;
        RECT 4.400 667.400 746.000 668.800 ;
        RECT 2.365 652.480 746.000 667.400 ;
        RECT 4.400 651.080 746.000 652.480 ;
        RECT 2.365 636.160 746.000 651.080 ;
        RECT 4.400 634.760 746.000 636.160 ;
        RECT 2.365 633.440 746.000 634.760 ;
        RECT 2.365 632.040 745.600 633.440 ;
        RECT 2.365 619.840 746.000 632.040 ;
        RECT 4.400 618.440 746.000 619.840 ;
        RECT 2.365 603.520 746.000 618.440 ;
        RECT 4.400 602.120 746.000 603.520 ;
        RECT 2.365 589.920 746.000 602.120 ;
        RECT 2.365 588.520 745.600 589.920 ;
        RECT 2.365 587.200 746.000 588.520 ;
        RECT 4.400 585.800 746.000 587.200 ;
        RECT 2.365 570.880 746.000 585.800 ;
        RECT 4.400 569.480 746.000 570.880 ;
        RECT 2.365 554.560 746.000 569.480 ;
        RECT 4.400 553.160 746.000 554.560 ;
        RECT 2.365 546.400 746.000 553.160 ;
        RECT 2.365 545.000 745.600 546.400 ;
        RECT 2.365 538.240 746.000 545.000 ;
        RECT 4.400 536.840 746.000 538.240 ;
        RECT 2.365 521.920 746.000 536.840 ;
        RECT 4.400 520.520 746.000 521.920 ;
        RECT 2.365 505.600 746.000 520.520 ;
        RECT 4.400 504.200 746.000 505.600 ;
        RECT 2.365 502.880 746.000 504.200 ;
        RECT 2.365 501.480 745.600 502.880 ;
        RECT 2.365 489.280 746.000 501.480 ;
        RECT 4.400 487.880 746.000 489.280 ;
        RECT 2.365 472.960 746.000 487.880 ;
        RECT 4.400 471.560 746.000 472.960 ;
        RECT 2.365 459.360 746.000 471.560 ;
        RECT 2.365 457.960 745.600 459.360 ;
        RECT 2.365 456.640 746.000 457.960 ;
        RECT 4.400 455.240 746.000 456.640 ;
        RECT 2.365 440.320 746.000 455.240 ;
        RECT 4.400 438.920 746.000 440.320 ;
        RECT 2.365 424.000 746.000 438.920 ;
        RECT 4.400 422.600 746.000 424.000 ;
        RECT 2.365 415.840 746.000 422.600 ;
        RECT 2.365 414.440 745.600 415.840 ;
        RECT 2.365 407.680 746.000 414.440 ;
        RECT 4.400 406.280 746.000 407.680 ;
        RECT 2.365 391.360 746.000 406.280 ;
        RECT 4.400 389.960 746.000 391.360 ;
        RECT 2.365 375.040 746.000 389.960 ;
        RECT 4.400 373.640 746.000 375.040 ;
        RECT 2.365 372.320 746.000 373.640 ;
        RECT 2.365 370.920 745.600 372.320 ;
        RECT 2.365 358.720 746.000 370.920 ;
        RECT 4.400 357.320 746.000 358.720 ;
        RECT 2.365 342.400 746.000 357.320 ;
        RECT 4.400 341.000 746.000 342.400 ;
        RECT 2.365 328.800 746.000 341.000 ;
        RECT 2.365 327.400 745.600 328.800 ;
        RECT 2.365 326.080 746.000 327.400 ;
        RECT 4.400 324.680 746.000 326.080 ;
        RECT 2.365 309.760 746.000 324.680 ;
        RECT 4.400 308.360 746.000 309.760 ;
        RECT 2.365 293.440 746.000 308.360 ;
        RECT 4.400 292.040 746.000 293.440 ;
        RECT 2.365 285.280 746.000 292.040 ;
        RECT 2.365 283.880 745.600 285.280 ;
        RECT 2.365 277.120 746.000 283.880 ;
        RECT 4.400 275.720 746.000 277.120 ;
        RECT 2.365 260.800 746.000 275.720 ;
        RECT 4.400 259.400 746.000 260.800 ;
        RECT 2.365 244.480 746.000 259.400 ;
        RECT 4.400 243.080 746.000 244.480 ;
        RECT 2.365 241.760 746.000 243.080 ;
        RECT 2.365 240.360 745.600 241.760 ;
        RECT 2.365 228.160 746.000 240.360 ;
        RECT 4.400 226.760 746.000 228.160 ;
        RECT 2.365 211.840 746.000 226.760 ;
        RECT 4.400 210.440 746.000 211.840 ;
        RECT 2.365 198.240 746.000 210.440 ;
        RECT 2.365 196.840 745.600 198.240 ;
        RECT 2.365 195.520 746.000 196.840 ;
        RECT 4.400 194.120 746.000 195.520 ;
        RECT 2.365 179.200 746.000 194.120 ;
        RECT 4.400 177.800 746.000 179.200 ;
        RECT 2.365 162.880 746.000 177.800 ;
        RECT 4.400 161.480 746.000 162.880 ;
        RECT 2.365 154.720 746.000 161.480 ;
        RECT 2.365 153.320 745.600 154.720 ;
        RECT 2.365 146.560 746.000 153.320 ;
        RECT 4.400 145.160 746.000 146.560 ;
        RECT 2.365 130.240 746.000 145.160 ;
        RECT 4.400 128.840 746.000 130.240 ;
        RECT 2.365 113.920 746.000 128.840 ;
        RECT 4.400 112.520 746.000 113.920 ;
        RECT 2.365 111.200 746.000 112.520 ;
        RECT 2.365 109.800 745.600 111.200 ;
        RECT 2.365 97.600 746.000 109.800 ;
        RECT 4.400 96.200 746.000 97.600 ;
        RECT 2.365 81.280 746.000 96.200 ;
        RECT 4.400 79.880 746.000 81.280 ;
        RECT 2.365 67.680 746.000 79.880 ;
        RECT 2.365 66.280 745.600 67.680 ;
        RECT 2.365 64.960 746.000 66.280 ;
        RECT 4.400 63.560 746.000 64.960 ;
        RECT 2.365 48.640 746.000 63.560 ;
        RECT 4.400 47.240 746.000 48.640 ;
        RECT 2.365 32.320 746.000 47.240 ;
        RECT 4.400 30.920 746.000 32.320 ;
        RECT 2.365 24.160 746.000 30.920 ;
        RECT 2.365 22.760 745.600 24.160 ;
        RECT 2.365 16.000 746.000 22.760 ;
        RECT 4.400 14.600 746.000 16.000 ;
        RECT 2.365 0.175 746.000 14.600 ;
      LAYER met4 ;
        RECT 3.975 10.240 20.640 686.625 ;
        RECT 23.040 10.240 97.440 686.625 ;
        RECT 99.840 10.240 174.240 686.625 ;
        RECT 176.640 10.240 251.040 686.625 ;
        RECT 253.440 10.240 327.840 686.625 ;
        RECT 330.240 10.240 404.640 686.625 ;
        RECT 407.040 10.240 481.440 686.625 ;
        RECT 483.840 10.240 558.240 686.625 ;
        RECT 560.640 10.240 635.040 686.625 ;
        RECT 637.440 10.240 641.850 686.625 ;
        RECT 3.975 3.575 641.850 10.240 ;
  END
END wrapped_tms1x00
END LIBRARY

